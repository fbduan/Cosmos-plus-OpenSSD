// BLH dynamic attribute configuration look-up table addresses
//
// Build Summary:
//    Built By:     blh_composer 3.0001
//    Built On:     Thu Aug 15 13:33:32 2013
//    Bundle:       GTHE3_CHANNEL
//    Architecture: olympus
//    Snapshot Dir: /tmp/E0n5cwkvI1
// Environment Variables:
//    XILENV=""
//    MYXILENV=""
//

`ifdef B_GTHE3_CHANNEL_DEFINES_VH
`else
`define B_GTHE3_CHANNEL_DEFINES_VH

// Look-up table parameters
//

`define GTHE3_CHANNEL_ADDR_N  388
`define GTHE3_CHANNEL_ADDR_SZ 32
`define GTHE3_CHANNEL_DATA_SZ 88

// Attribute addresses
//

`define GTHE3_CHANNEL__ACJTAG_DEBUG_MODE   	32'h0000	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__ACJTAG_DEBUG_MODE_SZ	1

`define GTHE3_CHANNEL__ACJTAG_MODE   	32'h0001	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__ACJTAG_MODE_SZ	1

`define GTHE3_CHANNEL__ACJTAG_RESET   	32'h0002	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__ACJTAG_RESET_SZ	1

`define GTHE3_CHANNEL__ADAPT_CFG0   	32'h0003	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__ADAPT_CFG0_SZ	16

`define GTHE3_CHANNEL__ADAPT_CFG1   	32'h0004	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__ADAPT_CFG1_SZ	16

`define GTHE3_CHANNEL__ALIGN_COMMA_DOUBLE   	32'h0005	// Type=STRING; Values=FALSE,TRUE
`define GTHE3_CHANNEL__ALIGN_COMMA_DOUBLE_SZ	40

`define GTHE3_CHANNEL__ALIGN_COMMA_ENABLE   	32'h0006	// Type=BINARY; Min=10'b0000000000, Max=10'b1111111111
`define GTHE3_CHANNEL__ALIGN_COMMA_ENABLE_SZ	10

`define GTHE3_CHANNEL__ALIGN_COMMA_WORD   	32'h0007	// Type=DECIMAL; Values=1,2,4
`define GTHE3_CHANNEL__ALIGN_COMMA_WORD_SZ	32

`define GTHE3_CHANNEL__ALIGN_MCOMMA_DET   	32'h0008	// Type=STRING; Values=TRUE,FALSE
`define GTHE3_CHANNEL__ALIGN_MCOMMA_DET_SZ	40

`define GTHE3_CHANNEL__ALIGN_MCOMMA_VALUE   	32'h0009	// Type=BINARY; Min=10'b0000000000, Max=10'b1111111111
`define GTHE3_CHANNEL__ALIGN_MCOMMA_VALUE_SZ	10

`define GTHE3_CHANNEL__ALIGN_PCOMMA_DET   	32'h000a	// Type=STRING; Values=TRUE,FALSE
`define GTHE3_CHANNEL__ALIGN_PCOMMA_DET_SZ	40

`define GTHE3_CHANNEL__ALIGN_PCOMMA_VALUE   	32'h000b	// Type=BINARY; Min=10'b0000000000, Max=10'b1111111111
`define GTHE3_CHANNEL__ALIGN_PCOMMA_VALUE_SZ	10

`define GTHE3_CHANNEL__A_RXOSCALRESET   	32'h000c	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__A_RXOSCALRESET_SZ	1

`define GTHE3_CHANNEL__A_RXPROGDIVRESET   	32'h000d	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__A_RXPROGDIVRESET_SZ	1

`define GTHE3_CHANNEL__A_TXPROGDIVRESET   	32'h000e	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__A_TXPROGDIVRESET_SZ	1

`define GTHE3_CHANNEL__CBCC_DATA_SOURCE_SEL   	32'h000f	// Type=STRING; Values=DECODED,ENCODED
`define GTHE3_CHANNEL__CBCC_DATA_SOURCE_SEL_SZ	56

`define GTHE3_CHANNEL__CDR_SWAP_MODE_EN   	32'h0010	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__CDR_SWAP_MODE_EN_SZ	1

`define GTHE3_CHANNEL__CHAN_BOND_KEEP_ALIGN   	32'h0011	// Type=STRING; Values=FALSE,TRUE
`define GTHE3_CHANNEL__CHAN_BOND_KEEP_ALIGN_SZ	40

`define GTHE3_CHANNEL__CHAN_BOND_MAX_SKEW   	32'h0012	// Type=DECIMAL; Values=7,1,2,3,4,5,6,8,9,10,11,12,13,14
`define GTHE3_CHANNEL__CHAN_BOND_MAX_SKEW_SZ	32

`define GTHE3_CHANNEL__CHAN_BOND_SEQ_1_1   	32'h0013	// Type=BINARY; Min=10'b0000000000, Max=10'b1111111111
`define GTHE3_CHANNEL__CHAN_BOND_SEQ_1_1_SZ	10

`define GTHE3_CHANNEL__CHAN_BOND_SEQ_1_2   	32'h0014	// Type=BINARY; Min=10'b0000000000, Max=10'b1111111111
`define GTHE3_CHANNEL__CHAN_BOND_SEQ_1_2_SZ	10

`define GTHE3_CHANNEL__CHAN_BOND_SEQ_1_3   	32'h0015	// Type=BINARY; Min=10'b0000000000, Max=10'b1111111111
`define GTHE3_CHANNEL__CHAN_BOND_SEQ_1_3_SZ	10

`define GTHE3_CHANNEL__CHAN_BOND_SEQ_1_4   	32'h0016	// Type=BINARY; Min=10'b0000000000, Max=10'b1111111111
`define GTHE3_CHANNEL__CHAN_BOND_SEQ_1_4_SZ	10

`define GTHE3_CHANNEL__CHAN_BOND_SEQ_1_ENABLE   	32'h0017	// Type=BINARY; Min=4'b0000, Max=4'b1111
`define GTHE3_CHANNEL__CHAN_BOND_SEQ_1_ENABLE_SZ	4

`define GTHE3_CHANNEL__CHAN_BOND_SEQ_2_1   	32'h0018	// Type=BINARY; Min=10'b0000000000, Max=10'b1111111111
`define GTHE3_CHANNEL__CHAN_BOND_SEQ_2_1_SZ	10

`define GTHE3_CHANNEL__CHAN_BOND_SEQ_2_2   	32'h0019	// Type=BINARY; Min=10'b0000000000, Max=10'b1111111111
`define GTHE3_CHANNEL__CHAN_BOND_SEQ_2_2_SZ	10

`define GTHE3_CHANNEL__CHAN_BOND_SEQ_2_3   	32'h001a	// Type=BINARY; Min=10'b0000000000, Max=10'b1111111111
`define GTHE3_CHANNEL__CHAN_BOND_SEQ_2_3_SZ	10

`define GTHE3_CHANNEL__CHAN_BOND_SEQ_2_4   	32'h001b	// Type=BINARY; Min=10'b0000000000, Max=10'b1111111111
`define GTHE3_CHANNEL__CHAN_BOND_SEQ_2_4_SZ	10

`define GTHE3_CHANNEL__CHAN_BOND_SEQ_2_ENABLE   	32'h001c	// Type=BINARY; Min=4'b0000, Max=4'b1111
`define GTHE3_CHANNEL__CHAN_BOND_SEQ_2_ENABLE_SZ	4

`define GTHE3_CHANNEL__CHAN_BOND_SEQ_2_USE   	32'h001d	// Type=STRING; Values=FALSE,TRUE
`define GTHE3_CHANNEL__CHAN_BOND_SEQ_2_USE_SZ	40

`define GTHE3_CHANNEL__CHAN_BOND_SEQ_LEN   	32'h001e	// Type=DECIMAL; Values=2,1,3,4
`define GTHE3_CHANNEL__CHAN_BOND_SEQ_LEN_SZ	32

`define GTHE3_CHANNEL__CLK_CORRECT_USE   	32'h001f	// Type=STRING; Values=TRUE,FALSE
`define GTHE3_CHANNEL__CLK_CORRECT_USE_SZ	40

`define GTHE3_CHANNEL__CLK_COR_KEEP_IDLE   	32'h0020	// Type=STRING; Values=FALSE,TRUE
`define GTHE3_CHANNEL__CLK_COR_KEEP_IDLE_SZ	40

`define GTHE3_CHANNEL__CLK_COR_MAX_LAT   	32'h0021	// Type=DECIMAL; Values=20,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,21,22,23,24,25,26,27,28,29,30,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60
`define GTHE3_CHANNEL__CLK_COR_MAX_LAT_SZ	32

`define GTHE3_CHANNEL__CLK_COR_MIN_LAT   	32'h0022	// Type=DECIMAL; Values=18,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,19,20,21,22,23,24,25,26,27,28,29,30,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63
`define GTHE3_CHANNEL__CLK_COR_MIN_LAT_SZ	32

`define GTHE3_CHANNEL__CLK_COR_PRECEDENCE   	32'h0023	// Type=STRING; Values=TRUE,FALSE
`define GTHE3_CHANNEL__CLK_COR_PRECEDENCE_SZ	40

`define GTHE3_CHANNEL__CLK_COR_REPEAT_WAIT   	32'h0024	// Type=DECIMAL; Values=0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,23,24,25,26,27,28,29,30,31
`define GTHE3_CHANNEL__CLK_COR_REPEAT_WAIT_SZ	32

`define GTHE3_CHANNEL__CLK_COR_SEQ_1_1   	32'h0025	// Type=BINARY; Min=10'b0000000000, Max=10'b1111111111
`define GTHE3_CHANNEL__CLK_COR_SEQ_1_1_SZ	10

`define GTHE3_CHANNEL__CLK_COR_SEQ_1_2   	32'h0026	// Type=BINARY; Min=10'b0000000000, Max=10'b1111111111
`define GTHE3_CHANNEL__CLK_COR_SEQ_1_2_SZ	10

`define GTHE3_CHANNEL__CLK_COR_SEQ_1_3   	32'h0027	// Type=BINARY; Min=10'b0000000000, Max=10'b1111111111
`define GTHE3_CHANNEL__CLK_COR_SEQ_1_3_SZ	10

`define GTHE3_CHANNEL__CLK_COR_SEQ_1_4   	32'h0028	// Type=BINARY; Min=10'b0000000000, Max=10'b1111111111
`define GTHE3_CHANNEL__CLK_COR_SEQ_1_4_SZ	10

`define GTHE3_CHANNEL__CLK_COR_SEQ_1_ENABLE   	32'h0029	// Type=BINARY; Min=4'b0000, Max=4'b1111
`define GTHE3_CHANNEL__CLK_COR_SEQ_1_ENABLE_SZ	4

`define GTHE3_CHANNEL__CLK_COR_SEQ_2_1   	32'h002a	// Type=BINARY; Min=10'b0000000000, Max=10'b1111111111
`define GTHE3_CHANNEL__CLK_COR_SEQ_2_1_SZ	10

`define GTHE3_CHANNEL__CLK_COR_SEQ_2_2   	32'h002b	// Type=BINARY; Min=10'b0000000000, Max=10'b1111111111
`define GTHE3_CHANNEL__CLK_COR_SEQ_2_2_SZ	10

`define GTHE3_CHANNEL__CLK_COR_SEQ_2_3   	32'h002c	// Type=BINARY; Min=10'b0000000000, Max=10'b1111111111
`define GTHE3_CHANNEL__CLK_COR_SEQ_2_3_SZ	10

`define GTHE3_CHANNEL__CLK_COR_SEQ_2_4   	32'h002d	// Type=BINARY; Min=10'b0000000000, Max=10'b1111111111
`define GTHE3_CHANNEL__CLK_COR_SEQ_2_4_SZ	10

`define GTHE3_CHANNEL__CLK_COR_SEQ_2_ENABLE   	32'h002e	// Type=BINARY; Min=4'b0000, Max=4'b1111
`define GTHE3_CHANNEL__CLK_COR_SEQ_2_ENABLE_SZ	4

`define GTHE3_CHANNEL__CLK_COR_SEQ_2_USE   	32'h002f	// Type=STRING; Values=FALSE,TRUE
`define GTHE3_CHANNEL__CLK_COR_SEQ_2_USE_SZ	40

`define GTHE3_CHANNEL__CLK_COR_SEQ_LEN   	32'h0030	// Type=DECIMAL; Values=2,1,3,4
`define GTHE3_CHANNEL__CLK_COR_SEQ_LEN_SZ	32

`define GTHE3_CHANNEL__CPLL_CFG0   	32'h0031	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__CPLL_CFG0_SZ	16

`define GTHE3_CHANNEL__CPLL_CFG1   	32'h0032	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__CPLL_CFG1_SZ	16

`define GTHE3_CHANNEL__CPLL_CFG2   	32'h0033	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__CPLL_CFG2_SZ	16

`define GTHE3_CHANNEL__CPLL_CFG3   	32'h0034	// Type=HEX; Min=6'h00, Max=6'h3f
`define GTHE3_CHANNEL__CPLL_CFG3_SZ	6

`define GTHE3_CHANNEL__CPLL_FBDIV   	32'h0035	// Type=DECIMAL; Values=4,1,2,3,5,6,8,10,12,16,20
`define GTHE3_CHANNEL__CPLL_FBDIV_SZ	32

`define GTHE3_CHANNEL__CPLL_FBDIV_45   	32'h0036	// Type=DECIMAL; Values=4,5
`define GTHE3_CHANNEL__CPLL_FBDIV_45_SZ	32

`define GTHE3_CHANNEL__CPLL_INIT_CFG0   	32'h0037	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__CPLL_INIT_CFG0_SZ	16

`define GTHE3_CHANNEL__CPLL_INIT_CFG1   	32'h0038	// Type=HEX; Min=8'h00, Max=8'hff
`define GTHE3_CHANNEL__CPLL_INIT_CFG1_SZ	8

`define GTHE3_CHANNEL__CPLL_LOCK_CFG   	32'h0039	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__CPLL_LOCK_CFG_SZ	16

`define GTHE3_CHANNEL__CPLL_REFCLK_DIV   	32'h003a	// Type=DECIMAL; Values=1,2,3,4,5,6,8,10,12,16,20
`define GTHE3_CHANNEL__CPLL_REFCLK_DIV_SZ	32

`define GTHE3_CHANNEL__DDI_CTRL   	32'h003b	// Type=BINARY; Min=2'b00, Max=2'b11
`define GTHE3_CHANNEL__DDI_CTRL_SZ	2

`define GTHE3_CHANNEL__DDI_REALIGN_WAIT   	32'h003c	// Type=DECIMAL; Values=15,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,16,17,18,19,20,21,22,23,24,25,26,27,28,29,30,31
`define GTHE3_CHANNEL__DDI_REALIGN_WAIT_SZ	32

`define GTHE3_CHANNEL__DEC_MCOMMA_DETECT   	32'h003d	// Type=STRING; Values=TRUE,FALSE
`define GTHE3_CHANNEL__DEC_MCOMMA_DETECT_SZ	40

`define GTHE3_CHANNEL__DEC_PCOMMA_DETECT   	32'h003e	// Type=STRING; Values=TRUE,FALSE
`define GTHE3_CHANNEL__DEC_PCOMMA_DETECT_SZ	40

`define GTHE3_CHANNEL__DEC_VALID_COMMA_ONLY   	32'h003f	// Type=STRING; Values=TRUE,FALSE
`define GTHE3_CHANNEL__DEC_VALID_COMMA_ONLY_SZ	40

`define GTHE3_CHANNEL__DFE_D_X_REL_POS   	32'h0040	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__DFE_D_X_REL_POS_SZ	1

`define GTHE3_CHANNEL__DFE_VCM_COMP_EN   	32'h0041	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__DFE_VCM_COMP_EN_SZ	1

`define GTHE3_CHANNEL__DMONITOR_CFG0   	32'h0042	// Type=HEX; Min=10'h000, Max=10'h3ff
`define GTHE3_CHANNEL__DMONITOR_CFG0_SZ	10

`define GTHE3_CHANNEL__DMONITOR_CFG1   	32'h0043	// Type=HEX; Min=8'h00, Max=8'hff
`define GTHE3_CHANNEL__DMONITOR_CFG1_SZ	8

`define GTHE3_CHANNEL__ES_CLK_PHASE_SEL   	32'h0044	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__ES_CLK_PHASE_SEL_SZ	1

`define GTHE3_CHANNEL__ES_CONTROL   	32'h0045	// Type=BINARY; Min=6'b000000, Max=6'b111111
`define GTHE3_CHANNEL__ES_CONTROL_SZ	6

`define GTHE3_CHANNEL__ES_ERRDET_EN   	32'h0046	// Type=STRING; Values=FALSE,TRUE
`define GTHE3_CHANNEL__ES_ERRDET_EN_SZ	40

`define GTHE3_CHANNEL__ES_EYE_SCAN_EN   	32'h0047	// Type=STRING; Values=FALSE,TRUE
`define GTHE3_CHANNEL__ES_EYE_SCAN_EN_SZ	40

`define GTHE3_CHANNEL__ES_HORZ_OFFSET   	32'h0048	// Type=HEX; Min=12'h000, Max=12'hfff
`define GTHE3_CHANNEL__ES_HORZ_OFFSET_SZ	12

`define GTHE3_CHANNEL__ES_PMA_CFG   	32'h0049	// Type=BINARY; Min=10'b0000000000, Max=10'b1111111111
`define GTHE3_CHANNEL__ES_PMA_CFG_SZ	10

`define GTHE3_CHANNEL__ES_PRESCALE   	32'h004a	// Type=BINARY; Min=5'b00000, Max=5'b11111
`define GTHE3_CHANNEL__ES_PRESCALE_SZ	5

`define GTHE3_CHANNEL__ES_QUALIFIER0   	32'h004b	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__ES_QUALIFIER0_SZ	16

`define GTHE3_CHANNEL__ES_QUALIFIER1   	32'h004c	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__ES_QUALIFIER1_SZ	16

`define GTHE3_CHANNEL__ES_QUALIFIER2   	32'h004d	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__ES_QUALIFIER2_SZ	16

`define GTHE3_CHANNEL__ES_QUALIFIER3   	32'h004e	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__ES_QUALIFIER3_SZ	16

`define GTHE3_CHANNEL__ES_QUALIFIER4   	32'h004f	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__ES_QUALIFIER4_SZ	16

`define GTHE3_CHANNEL__ES_QUAL_MASK0   	32'h0050	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__ES_QUAL_MASK0_SZ	16

`define GTHE3_CHANNEL__ES_QUAL_MASK1   	32'h0051	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__ES_QUAL_MASK1_SZ	16

`define GTHE3_CHANNEL__ES_QUAL_MASK2   	32'h0052	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__ES_QUAL_MASK2_SZ	16

`define GTHE3_CHANNEL__ES_QUAL_MASK3   	32'h0053	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__ES_QUAL_MASK3_SZ	16

`define GTHE3_CHANNEL__ES_QUAL_MASK4   	32'h0054	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__ES_QUAL_MASK4_SZ	16

`define GTHE3_CHANNEL__ES_SDATA_MASK0   	32'h0055	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__ES_SDATA_MASK0_SZ	16

`define GTHE3_CHANNEL__ES_SDATA_MASK1   	32'h0056	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__ES_SDATA_MASK1_SZ	16

`define GTHE3_CHANNEL__ES_SDATA_MASK2   	32'h0057	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__ES_SDATA_MASK2_SZ	16

`define GTHE3_CHANNEL__ES_SDATA_MASK3   	32'h0058	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__ES_SDATA_MASK3_SZ	16

`define GTHE3_CHANNEL__ES_SDATA_MASK4   	32'h0059	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__ES_SDATA_MASK4_SZ	16

`define GTHE3_CHANNEL__EVODD_PHI_CFG   	32'h005a	// Type=BINARY; Min=11'b00000000000, Max=11'b11111111111
`define GTHE3_CHANNEL__EVODD_PHI_CFG_SZ	11

`define GTHE3_CHANNEL__EYE_SCAN_SWAP_EN   	32'h005b	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__EYE_SCAN_SWAP_EN_SZ	1

`define GTHE3_CHANNEL__FTS_DESKEW_SEQ_ENABLE   	32'h005c	// Type=BINARY; Min=4'b0000, Max=4'b1111
`define GTHE3_CHANNEL__FTS_DESKEW_SEQ_ENABLE_SZ	4

`define GTHE3_CHANNEL__FTS_LANE_DESKEW_CFG   	32'h005d	// Type=BINARY; Min=4'b0000, Max=4'b1111
`define GTHE3_CHANNEL__FTS_LANE_DESKEW_CFG_SZ	4

`define GTHE3_CHANNEL__FTS_LANE_DESKEW_EN   	32'h005e	// Type=STRING; Values=FALSE,TRUE
`define GTHE3_CHANNEL__FTS_LANE_DESKEW_EN_SZ	40

`define GTHE3_CHANNEL__GEARBOX_MODE   	32'h005f	// Type=BINARY; Min=5'b00000, Max=5'b11111
`define GTHE3_CHANNEL__GEARBOX_MODE_SZ	5

`define GTHE3_CHANNEL__GM_BIAS_SELECT   	32'h0060	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__GM_BIAS_SELECT_SZ	1

`define GTHE3_CHANNEL__LOCAL_MASTER   	32'h0061	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__LOCAL_MASTER_SZ	1

`define GTHE3_CHANNEL__OOBDIVCTL   	32'h0062	// Type=BINARY; Min=2'b00, Max=2'b11
`define GTHE3_CHANNEL__OOBDIVCTL_SZ	2

`define GTHE3_CHANNEL__OOB_PWRUP   	32'h0063	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__OOB_PWRUP_SZ	1

`define GTHE3_CHANNEL__PCI3_AUTO_REALIGN   	32'h0064	// Type=STRING; Values=FRST_SMPL,OVR_1K_BLK,OVR_8_BLK,OVR_64_BLK
`define GTHE3_CHANNEL__PCI3_AUTO_REALIGN_SZ	80

`define GTHE3_CHANNEL__PCI3_PIPE_RX_ELECIDLE   	32'h0065	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__PCI3_PIPE_RX_ELECIDLE_SZ	1

`define GTHE3_CHANNEL__PCI3_RX_ASYNC_EBUF_BYPASS   	32'h0066	// Type=BINARY; Min=2'b00, Max=2'b11
`define GTHE3_CHANNEL__PCI3_RX_ASYNC_EBUF_BYPASS_SZ	2

`define GTHE3_CHANNEL__PCI3_RX_ELECIDLE_EI2_ENABLE   	32'h0067	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__PCI3_RX_ELECIDLE_EI2_ENABLE_SZ	1

`define GTHE3_CHANNEL__PCI3_RX_ELECIDLE_H2L_COUNT   	32'h0068	// Type=BINARY; Min=6'b000000, Max=6'b111111
`define GTHE3_CHANNEL__PCI3_RX_ELECIDLE_H2L_COUNT_SZ	6

`define GTHE3_CHANNEL__PCI3_RX_ELECIDLE_H2L_DISABLE   	32'h0069	// Type=BINARY; Min=3'b000, Max=3'b111
`define GTHE3_CHANNEL__PCI3_RX_ELECIDLE_H2L_DISABLE_SZ	3

`define GTHE3_CHANNEL__PCI3_RX_ELECIDLE_HI_COUNT   	32'h006a	// Type=BINARY; Min=6'b000000, Max=6'b111111
`define GTHE3_CHANNEL__PCI3_RX_ELECIDLE_HI_COUNT_SZ	6

`define GTHE3_CHANNEL__PCI3_RX_ELECIDLE_LP4_DISABLE   	32'h006b	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__PCI3_RX_ELECIDLE_LP4_DISABLE_SZ	1

`define GTHE3_CHANNEL__PCI3_RX_FIFO_DISABLE   	32'h006c	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__PCI3_RX_FIFO_DISABLE_SZ	1

`define GTHE3_CHANNEL__PCIE_BUFG_DIV_CTRL   	32'h006d	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__PCIE_BUFG_DIV_CTRL_SZ	16

`define GTHE3_CHANNEL__PCIE_RXPCS_CFG_GEN3   	32'h006e	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__PCIE_RXPCS_CFG_GEN3_SZ	16

`define GTHE3_CHANNEL__PCIE_RXPMA_CFG   	32'h006f	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__PCIE_RXPMA_CFG_SZ	16

`define GTHE3_CHANNEL__PCIE_TXPCS_CFG_GEN3   	32'h0070	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__PCIE_TXPCS_CFG_GEN3_SZ	16

`define GTHE3_CHANNEL__PCIE_TXPMA_CFG   	32'h0071	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__PCIE_TXPMA_CFG_SZ	16

`define GTHE3_CHANNEL__PCS_PCIE_EN   	32'h0072	// Type=STRING; Values=FALSE,TRUE
`define GTHE3_CHANNEL__PCS_PCIE_EN_SZ	40

`define GTHE3_CHANNEL__PCS_RSVD0   	32'h0073	// Type=BINARY; Min=16'b0000000000000000, Max=16'b1111111111111111
`define GTHE3_CHANNEL__PCS_RSVD0_SZ	16

`define GTHE3_CHANNEL__PCS_RSVD1   	32'h0074	// Type=BINARY; Min=3'b000, Max=3'b111
`define GTHE3_CHANNEL__PCS_RSVD1_SZ	3

`define GTHE3_CHANNEL__PD_TRANS_TIME_FROM_P2   	32'h0075	// Type=HEX; Min=12'h000, Max=12'hfff
`define GTHE3_CHANNEL__PD_TRANS_TIME_FROM_P2_SZ	12

`define GTHE3_CHANNEL__PD_TRANS_TIME_NONE_P2   	32'h0076	// Type=HEX; Min=8'h00, Max=8'hff
`define GTHE3_CHANNEL__PD_TRANS_TIME_NONE_P2_SZ	8

`define GTHE3_CHANNEL__PD_TRANS_TIME_TO_P2   	32'h0077	// Type=HEX; Min=8'h00, Max=8'hff
`define GTHE3_CHANNEL__PD_TRANS_TIME_TO_P2_SZ	8

`define GTHE3_CHANNEL__PLL_SEL_MODE_GEN12   	32'h0078	// Type=HEX; Min=2'h0, Max=2'h3
`define GTHE3_CHANNEL__PLL_SEL_MODE_GEN12_SZ	2

`define GTHE3_CHANNEL__PLL_SEL_MODE_GEN3   	32'h0079	// Type=HEX; Min=2'h0, Max=2'h3
`define GTHE3_CHANNEL__PLL_SEL_MODE_GEN3_SZ	2

`define GTHE3_CHANNEL__PMA_RSV1   	32'h007a	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__PMA_RSV1_SZ	16

`define GTHE3_CHANNEL__PROCESS_PAR   	32'h007b	// Type=BINARY; Min=3'b000, Max=3'b111
`define GTHE3_CHANNEL__PROCESS_PAR_SZ	3

`define GTHE3_CHANNEL__RATE_SW_USE_DRP   	32'h007c	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RATE_SW_USE_DRP_SZ	1

`define GTHE3_CHANNEL__RESET_POWERSAVE_DISABLE   	32'h007d	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RESET_POWERSAVE_DISABLE_SZ	1

`define GTHE3_CHANNEL__RXBUFRESET_TIME   	32'h007e	// Type=BINARY; Min=5'b00000, Max=5'b11111
`define GTHE3_CHANNEL__RXBUFRESET_TIME_SZ	5

`define GTHE3_CHANNEL__RXBUF_ADDR_MODE   	32'h007f	// Type=STRING; Values=FULL,FAST
`define GTHE3_CHANNEL__RXBUF_ADDR_MODE_SZ	32

`define GTHE3_CHANNEL__RXBUF_EIDLE_HI_CNT   	32'h0080	// Type=BINARY; Min=4'b0000, Max=4'b1111
`define GTHE3_CHANNEL__RXBUF_EIDLE_HI_CNT_SZ	4

`define GTHE3_CHANNEL__RXBUF_EIDLE_LO_CNT   	32'h0081	// Type=BINARY; Min=4'b0000, Max=4'b1111
`define GTHE3_CHANNEL__RXBUF_EIDLE_LO_CNT_SZ	4

`define GTHE3_CHANNEL__RXBUF_EN   	32'h0082	// Type=STRING; Values=TRUE,FALSE
`define GTHE3_CHANNEL__RXBUF_EN_SZ	40

`define GTHE3_CHANNEL__RXBUF_RESET_ON_CB_CHANGE   	32'h0083	// Type=STRING; Values=TRUE,FALSE
`define GTHE3_CHANNEL__RXBUF_RESET_ON_CB_CHANGE_SZ	40

`define GTHE3_CHANNEL__RXBUF_RESET_ON_COMMAALIGN   	32'h0084	// Type=STRING; Values=FALSE,TRUE
`define GTHE3_CHANNEL__RXBUF_RESET_ON_COMMAALIGN_SZ	40

`define GTHE3_CHANNEL__RXBUF_RESET_ON_EIDLE   	32'h0085	// Type=STRING; Values=FALSE,TRUE
`define GTHE3_CHANNEL__RXBUF_RESET_ON_EIDLE_SZ	40

`define GTHE3_CHANNEL__RXBUF_RESET_ON_RATE_CHANGE   	32'h0086	// Type=STRING; Values=TRUE,FALSE
`define GTHE3_CHANNEL__RXBUF_RESET_ON_RATE_CHANGE_SZ	40

`define GTHE3_CHANNEL__RXBUF_THRESH_OVFLW   	32'h0087	// Type=DECIMAL; Values=0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,23,24,25,26,27,28,29,30,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63
`define GTHE3_CHANNEL__RXBUF_THRESH_OVFLW_SZ	32

`define GTHE3_CHANNEL__RXBUF_THRESH_OVRD   	32'h0088	// Type=STRING; Values=FALSE,TRUE
`define GTHE3_CHANNEL__RXBUF_THRESH_OVRD_SZ	40

`define GTHE3_CHANNEL__RXBUF_THRESH_UNDFLW   	32'h0089	// Type=DECIMAL; Values=4,0,1,2,3,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,23,24,25,26,27,28,29,30,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63
`define GTHE3_CHANNEL__RXBUF_THRESH_UNDFLW_SZ	32

`define GTHE3_CHANNEL__RXCDRFREQRESET_TIME   	32'h008a	// Type=BINARY; Min=5'b00000, Max=5'b11111
`define GTHE3_CHANNEL__RXCDRFREQRESET_TIME_SZ	5

`define GTHE3_CHANNEL__RXCDRPHRESET_TIME   	32'h008b	// Type=BINARY; Min=5'b00000, Max=5'b11111
`define GTHE3_CHANNEL__RXCDRPHRESET_TIME_SZ	5

`define GTHE3_CHANNEL__RXCDR_CFG0   	32'h008c	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXCDR_CFG0_SZ	16

`define GTHE3_CHANNEL__RXCDR_CFG0_GEN3   	32'h008d	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXCDR_CFG0_GEN3_SZ	16

`define GTHE3_CHANNEL__RXCDR_CFG1   	32'h008e	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXCDR_CFG1_SZ	16

`define GTHE3_CHANNEL__RXCDR_CFG1_GEN3   	32'h008f	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXCDR_CFG1_GEN3_SZ	16

`define GTHE3_CHANNEL__RXCDR_CFG2   	32'h0090	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXCDR_CFG2_SZ	16

`define GTHE3_CHANNEL__RXCDR_CFG2_GEN3   	32'h0091	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXCDR_CFG2_GEN3_SZ	16

`define GTHE3_CHANNEL__RXCDR_CFG3   	32'h0092	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXCDR_CFG3_SZ	16

`define GTHE3_CHANNEL__RXCDR_CFG3_GEN3   	32'h0093	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXCDR_CFG3_GEN3_SZ	16

`define GTHE3_CHANNEL__RXCDR_CFG4   	32'h0094	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXCDR_CFG4_SZ	16

`define GTHE3_CHANNEL__RXCDR_CFG4_GEN3   	32'h0095	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXCDR_CFG4_GEN3_SZ	16

`define GTHE3_CHANNEL__RXCDR_CFG5   	32'h0096	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXCDR_CFG5_SZ	16

`define GTHE3_CHANNEL__RXCDR_CFG5_GEN3   	32'h0097	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXCDR_CFG5_GEN3_SZ	16

`define GTHE3_CHANNEL__RXCDR_FR_RESET_ON_EIDLE   	32'h0098	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RXCDR_FR_RESET_ON_EIDLE_SZ	1

`define GTHE3_CHANNEL__RXCDR_HOLD_DURING_EIDLE   	32'h0099	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RXCDR_HOLD_DURING_EIDLE_SZ	1

`define GTHE3_CHANNEL__RXCDR_LOCK_CFG0   	32'h009a	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXCDR_LOCK_CFG0_SZ	16

`define GTHE3_CHANNEL__RXCDR_LOCK_CFG1   	32'h009b	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXCDR_LOCK_CFG1_SZ	16

`define GTHE3_CHANNEL__RXCDR_LOCK_CFG2   	32'h009c	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXCDR_LOCK_CFG2_SZ	16

`define GTHE3_CHANNEL__RXCDR_PH_RESET_ON_EIDLE   	32'h009d	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RXCDR_PH_RESET_ON_EIDLE_SZ	1

`define GTHE3_CHANNEL__RXCFOK_CFG0   	32'h009e	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXCFOK_CFG0_SZ	16

`define GTHE3_CHANNEL__RXCFOK_CFG1   	32'h009f	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXCFOK_CFG1_SZ	16

`define GTHE3_CHANNEL__RXCFOK_CFG2   	32'h00a0	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXCFOK_CFG2_SZ	16

`define GTHE3_CHANNEL__RXDFELPMRESET_TIME   	32'h00a1	// Type=BINARY; Min=7'b0000000, Max=7'b1111111
`define GTHE3_CHANNEL__RXDFELPMRESET_TIME_SZ	7

`define GTHE3_CHANNEL__RXDFELPM_KL_CFG0   	32'h00a2	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFELPM_KL_CFG0_SZ	16

`define GTHE3_CHANNEL__RXDFELPM_KL_CFG1   	32'h00a3	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFELPM_KL_CFG1_SZ	16

`define GTHE3_CHANNEL__RXDFELPM_KL_CFG2   	32'h00a4	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFELPM_KL_CFG2_SZ	16

`define GTHE3_CHANNEL__RXDFE_CFG0   	32'h00a5	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_CFG0_SZ	16

`define GTHE3_CHANNEL__RXDFE_CFG1   	32'h00a6	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_CFG1_SZ	16

`define GTHE3_CHANNEL__RXDFE_GC_CFG0   	32'h00a7	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_GC_CFG0_SZ	16

`define GTHE3_CHANNEL__RXDFE_GC_CFG1   	32'h00a8	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_GC_CFG1_SZ	16

`define GTHE3_CHANNEL__RXDFE_GC_CFG2   	32'h00a9	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_GC_CFG2_SZ	16

`define GTHE3_CHANNEL__RXDFE_H2_CFG0   	32'h00aa	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_H2_CFG0_SZ	16

`define GTHE3_CHANNEL__RXDFE_H2_CFG1   	32'h00ab	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_H2_CFG1_SZ	16

`define GTHE3_CHANNEL__RXDFE_H3_CFG0   	32'h00ac	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_H3_CFG0_SZ	16

`define GTHE3_CHANNEL__RXDFE_H3_CFG1   	32'h00ad	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_H3_CFG1_SZ	16

`define GTHE3_CHANNEL__RXDFE_H4_CFG0   	32'h00ae	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_H4_CFG0_SZ	16

`define GTHE3_CHANNEL__RXDFE_H4_CFG1   	32'h00af	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_H4_CFG1_SZ	16

`define GTHE3_CHANNEL__RXDFE_H5_CFG0   	32'h00b0	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_H5_CFG0_SZ	16

`define GTHE3_CHANNEL__RXDFE_H5_CFG1   	32'h00b1	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_H5_CFG1_SZ	16

`define GTHE3_CHANNEL__RXDFE_H6_CFG0   	32'h00b2	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_H6_CFG0_SZ	16

`define GTHE3_CHANNEL__RXDFE_H6_CFG1   	32'h00b3	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_H6_CFG1_SZ	16

`define GTHE3_CHANNEL__RXDFE_H7_CFG0   	32'h00b4	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_H7_CFG0_SZ	16

`define GTHE3_CHANNEL__RXDFE_H7_CFG1   	32'h00b5	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_H7_CFG1_SZ	16

`define GTHE3_CHANNEL__RXDFE_H8_CFG0   	32'h00b6	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_H8_CFG0_SZ	16

`define GTHE3_CHANNEL__RXDFE_H8_CFG1   	32'h00b7	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_H8_CFG1_SZ	16

`define GTHE3_CHANNEL__RXDFE_H9_CFG0   	32'h00b8	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_H9_CFG0_SZ	16

`define GTHE3_CHANNEL__RXDFE_H9_CFG1   	32'h00b9	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_H9_CFG1_SZ	16

`define GTHE3_CHANNEL__RXDFE_HA_CFG0   	32'h00ba	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_HA_CFG0_SZ	16

`define GTHE3_CHANNEL__RXDFE_HA_CFG1   	32'h00bb	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_HA_CFG1_SZ	16

`define GTHE3_CHANNEL__RXDFE_HB_CFG0   	32'h00bc	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_HB_CFG0_SZ	16

`define GTHE3_CHANNEL__RXDFE_HB_CFG1   	32'h00bd	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_HB_CFG1_SZ	16

`define GTHE3_CHANNEL__RXDFE_HC_CFG0   	32'h00be	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_HC_CFG0_SZ	16

`define GTHE3_CHANNEL__RXDFE_HC_CFG1   	32'h00bf	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_HC_CFG1_SZ	16

`define GTHE3_CHANNEL__RXDFE_HD_CFG0   	32'h00c0	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_HD_CFG0_SZ	16

`define GTHE3_CHANNEL__RXDFE_HD_CFG1   	32'h00c1	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_HD_CFG1_SZ	16

`define GTHE3_CHANNEL__RXDFE_HE_CFG0   	32'h00c2	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_HE_CFG0_SZ	16

`define GTHE3_CHANNEL__RXDFE_HE_CFG1   	32'h00c3	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_HE_CFG1_SZ	16

`define GTHE3_CHANNEL__RXDFE_HF_CFG0   	32'h00c4	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_HF_CFG0_SZ	16

`define GTHE3_CHANNEL__RXDFE_HF_CFG1   	32'h00c5	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_HF_CFG1_SZ	16

`define GTHE3_CHANNEL__RXDFE_OS_CFG0   	32'h00c6	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_OS_CFG0_SZ	16

`define GTHE3_CHANNEL__RXDFE_OS_CFG1   	32'h00c7	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_OS_CFG1_SZ	16

`define GTHE3_CHANNEL__RXDFE_UT_CFG0   	32'h00c8	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_UT_CFG0_SZ	16

`define GTHE3_CHANNEL__RXDFE_UT_CFG1   	32'h00c9	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_UT_CFG1_SZ	16

`define GTHE3_CHANNEL__RXDFE_VP_CFG0   	32'h00ca	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_VP_CFG0_SZ	16

`define GTHE3_CHANNEL__RXDFE_VP_CFG1   	32'h00cb	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDFE_VP_CFG1_SZ	16

`define GTHE3_CHANNEL__RXDLY_CFG   	32'h00cc	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDLY_CFG_SZ	16

`define GTHE3_CHANNEL__RXDLY_LCFG   	32'h00cd	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXDLY_LCFG_SZ	16

`define GTHE3_CHANNEL__RXELECIDLE_CFG   	32'h00ce	// Type=STRING; Values=Sigcfg_4,Sigcfg_1,Sigcfg_2,Sigcfg_3,Sigcfg_6,Sigcfg_8,Sigcfg_12,Sigcfg_16
`define GTHE3_CHANNEL__RXELECIDLE_CFG_SZ	72

`define GTHE3_CHANNEL__RXGBOX_FIFO_INIT_RD_ADDR   	32'h00cf	// Type=DECIMAL; Values=4,2,3,5
`define GTHE3_CHANNEL__RXGBOX_FIFO_INIT_RD_ADDR_SZ	32

`define GTHE3_CHANNEL__RXGEARBOX_EN   	32'h00d0	// Type=STRING; Values=FALSE,TRUE
`define GTHE3_CHANNEL__RXGEARBOX_EN_SZ	40

`define GTHE3_CHANNEL__RXISCANRESET_TIME   	32'h00d1	// Type=BINARY; Min=5'b00000, Max=5'b11111
`define GTHE3_CHANNEL__RXISCANRESET_TIME_SZ	5

`define GTHE3_CHANNEL__RXLPM_CFG   	32'h00d2	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXLPM_CFG_SZ	16

`define GTHE3_CHANNEL__RXLPM_GC_CFG   	32'h00d3	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXLPM_GC_CFG_SZ	16

`define GTHE3_CHANNEL__RXLPM_KH_CFG0   	32'h00d4	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXLPM_KH_CFG0_SZ	16

`define GTHE3_CHANNEL__RXLPM_KH_CFG1   	32'h00d5	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXLPM_KH_CFG1_SZ	16

`define GTHE3_CHANNEL__RXLPM_OS_CFG0   	32'h00d6	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXLPM_OS_CFG0_SZ	16

`define GTHE3_CHANNEL__RXLPM_OS_CFG1   	32'h00d7	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXLPM_OS_CFG1_SZ	16

`define GTHE3_CHANNEL__RXOOB_CFG   	32'h00d8	// Type=BINARY; Min=9'b000000000, Max=9'b111111111
`define GTHE3_CHANNEL__RXOOB_CFG_SZ	9

`define GTHE3_CHANNEL__RXOOB_CLK_CFG   	32'h00d9	// Type=STRING; Values=PMA,FABRIC
`define GTHE3_CHANNEL__RXOOB_CLK_CFG_SZ	48

`define GTHE3_CHANNEL__RXOSCALRESET_TIME   	32'h00da	// Type=BINARY; Min=5'b00000, Max=5'b11111
`define GTHE3_CHANNEL__RXOSCALRESET_TIME_SZ	5

`define GTHE3_CHANNEL__RXOUT_DIV   	32'h00db	// Type=DECIMAL; Values=4,1,2,8,16
`define GTHE3_CHANNEL__RXOUT_DIV_SZ	32

`define GTHE3_CHANNEL__RXPCSRESET_TIME   	32'h00dc	// Type=BINARY; Min=5'b00000, Max=5'b11111
`define GTHE3_CHANNEL__RXPCSRESET_TIME_SZ	5

`define GTHE3_CHANNEL__RXPHBEACON_CFG   	32'h00dd	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXPHBEACON_CFG_SZ	16

`define GTHE3_CHANNEL__RXPHDLY_CFG   	32'h00de	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXPHDLY_CFG_SZ	16

`define GTHE3_CHANNEL__RXPHSAMP_CFG   	32'h00df	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXPHSAMP_CFG_SZ	16

`define GTHE3_CHANNEL__RXPHSLIP_CFG   	32'h00e0	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RXPHSLIP_CFG_SZ	16

`define GTHE3_CHANNEL__RXPH_MONITOR_SEL   	32'h00e1	// Type=BINARY; Min=5'b00000, Max=5'b11111
`define GTHE3_CHANNEL__RXPH_MONITOR_SEL_SZ	5

`define GTHE3_CHANNEL__RXPI_CFG0   	32'h00e2	// Type=BINARY; Min=2'b00, Max=2'b11
`define GTHE3_CHANNEL__RXPI_CFG0_SZ	2

`define GTHE3_CHANNEL__RXPI_CFG1   	32'h00e3	// Type=BINARY; Min=2'b00, Max=2'b11
`define GTHE3_CHANNEL__RXPI_CFG1_SZ	2

`define GTHE3_CHANNEL__RXPI_CFG2   	32'h00e4	// Type=BINARY; Min=2'b00, Max=2'b11
`define GTHE3_CHANNEL__RXPI_CFG2_SZ	2

`define GTHE3_CHANNEL__RXPI_CFG3   	32'h00e5	// Type=BINARY; Min=2'b00, Max=2'b11
`define GTHE3_CHANNEL__RXPI_CFG3_SZ	2

`define GTHE3_CHANNEL__RXPI_CFG4   	32'h00e6	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RXPI_CFG4_SZ	1

`define GTHE3_CHANNEL__RXPI_CFG5   	32'h00e7	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RXPI_CFG5_SZ	1

`define GTHE3_CHANNEL__RXPI_CFG6   	32'h00e8	// Type=BINARY; Min=3'b000, Max=3'b111
`define GTHE3_CHANNEL__RXPI_CFG6_SZ	3

`define GTHE3_CHANNEL__RXPI_LPM   	32'h00e9	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RXPI_LPM_SZ	1

`define GTHE3_CHANNEL__RXPI_VREFSEL   	32'h00ea	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RXPI_VREFSEL_SZ	1

`define GTHE3_CHANNEL__RXPMACLK_SEL   	32'h00eb	// Type=STRING; Values=DATA,CROSSING,EYESCAN
`define GTHE3_CHANNEL__RXPMACLK_SEL_SZ	64

`define GTHE3_CHANNEL__RXPMARESET_TIME   	32'h00ec	// Type=BINARY; Min=5'b00000, Max=5'b11111
`define GTHE3_CHANNEL__RXPMARESET_TIME_SZ	5

`define GTHE3_CHANNEL__RXPRBS_ERR_LOOPBACK   	32'h00ed	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RXPRBS_ERR_LOOPBACK_SZ	1

`define GTHE3_CHANNEL__RXPRBS_LINKACQ_CNT   	32'h00ee	// Type=DECIMAL; Values=15,16,17,18,19,20,21,22,23,24,25,26,27,28,29,30,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,148,149,150,151,152,153,154,155,156,157,158,159,160,161,162,163,164,165,166,167,168,169,170,171,172,173,174,175,176,177,178,179,180,181,182,183,184,185,186,187,188,189,190,191,192,193,194,195,196,197,198,199,200,201,202,203,204,205,206,207,208,209,210,211,212,213,214,215,216,217,218,219,220,221,222,223,224,225,226,227,228,229,230,231,232,233,234,235,236,237,238,239,240,241,242,243,244,245,246,247,248,249,250,251,252,253,254,255
`define GTHE3_CHANNEL__RXPRBS_LINKACQ_CNT_SZ	32

`define GTHE3_CHANNEL__RXSLIDE_AUTO_WAIT   	32'h00ef	// Type=DECIMAL; Values=7,1,2,3,4,5,6,8,9,10,11,12,13,14,15
`define GTHE3_CHANNEL__RXSLIDE_AUTO_WAIT_SZ	32

`define GTHE3_CHANNEL__RXSLIDE_MODE   	32'h00f0	// Type=STRING; Values=OFF,AUTO,PCS,PMA
`define GTHE3_CHANNEL__RXSLIDE_MODE_SZ	32

`define GTHE3_CHANNEL__RXSYNC_MULTILANE   	32'h00f1	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RXSYNC_MULTILANE_SZ	1

`define GTHE3_CHANNEL__RXSYNC_OVRD   	32'h00f2	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RXSYNC_OVRD_SZ	1

`define GTHE3_CHANNEL__RXSYNC_SKIP_DA   	32'h00f3	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RXSYNC_SKIP_DA_SZ	1

`define GTHE3_CHANNEL__RX_AFE_CM_EN   	32'h00f4	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RX_AFE_CM_EN_SZ	1

`define GTHE3_CHANNEL__RX_BIAS_CFG0   	32'h00f5	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__RX_BIAS_CFG0_SZ	16

`define GTHE3_CHANNEL__RX_BUFFER_CFG   	32'h00f6	// Type=BINARY; Min=6'b000000, Max=6'b111111
`define GTHE3_CHANNEL__RX_BUFFER_CFG_SZ	6

`define GTHE3_CHANNEL__RX_CAPFF_SARC_ENB   	32'h00f7	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RX_CAPFF_SARC_ENB_SZ	1

`define GTHE3_CHANNEL__RX_CLK25_DIV   	32'h00f8	// Type=DECIMAL; Values=8,1,2,3,4,5,6,7,9,10,11,12,13,14,15,16,17,18,19,20,21,22,23,24,25,26,27,28,29,30,31,32
`define GTHE3_CHANNEL__RX_CLK25_DIV_SZ	32

`define GTHE3_CHANNEL__RX_CLKMUX_EN   	32'h00f9	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RX_CLKMUX_EN_SZ	1

`define GTHE3_CHANNEL__RX_CLK_SLIP_OVRD   	32'h00fa	// Type=BINARY; Min=5'b00000, Max=5'b11111
`define GTHE3_CHANNEL__RX_CLK_SLIP_OVRD_SZ	5

`define GTHE3_CHANNEL__RX_CM_BUF_CFG   	32'h00fb	// Type=BINARY; Min=4'b0000, Max=4'b1111
`define GTHE3_CHANNEL__RX_CM_BUF_CFG_SZ	4

`define GTHE3_CHANNEL__RX_CM_BUF_PD   	32'h00fc	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RX_CM_BUF_PD_SZ	1

`define GTHE3_CHANNEL__RX_CM_SEL   	32'h00fd	// Type=BINARY; Min=2'b00, Max=2'b11
`define GTHE3_CHANNEL__RX_CM_SEL_SZ	2

`define GTHE3_CHANNEL__RX_CM_TRIM   	32'h00fe	// Type=BINARY; Min=4'b0000, Max=4'b1111
`define GTHE3_CHANNEL__RX_CM_TRIM_SZ	4

`define GTHE3_CHANNEL__RX_CTLE3_LPF   	32'h00ff	// Type=BINARY; Min=8'b00000000, Max=8'b11111111
`define GTHE3_CHANNEL__RX_CTLE3_LPF_SZ	8

`define GTHE3_CHANNEL__RX_DATA_WIDTH   	32'h0100	// Type=DECIMAL; Values=20,16,32,40,64,80,128,160
`define GTHE3_CHANNEL__RX_DATA_WIDTH_SZ	32

`define GTHE3_CHANNEL__RX_DDI_SEL   	32'h0101	// Type=BINARY; Min=6'b000000, Max=6'b111111
`define GTHE3_CHANNEL__RX_DDI_SEL_SZ	6

`define GTHE3_CHANNEL__RX_DEFER_RESET_BUF_EN   	32'h0102	// Type=STRING; Values=TRUE,FALSE
`define GTHE3_CHANNEL__RX_DEFER_RESET_BUF_EN_SZ	40

`define GTHE3_CHANNEL__RX_DFELPM_CFG0   	32'h0103	// Type=BINARY; Min=4'b0000, Max=4'b1111
`define GTHE3_CHANNEL__RX_DFELPM_CFG0_SZ	4

`define GTHE3_CHANNEL__RX_DFELPM_CFG1   	32'h0104	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RX_DFELPM_CFG1_SZ	1

`define GTHE3_CHANNEL__RX_DFELPM_KLKH_AGC_STUP_EN   	32'h0105	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RX_DFELPM_KLKH_AGC_STUP_EN_SZ	1

`define GTHE3_CHANNEL__RX_DFE_AGC_CFG0   	32'h0106	// Type=BINARY; Min=2'b00, Max=2'b11
`define GTHE3_CHANNEL__RX_DFE_AGC_CFG0_SZ	2

`define GTHE3_CHANNEL__RX_DFE_AGC_CFG1   	32'h0107	// Type=BINARY; Min=3'b000, Max=3'b111
`define GTHE3_CHANNEL__RX_DFE_AGC_CFG1_SZ	3

`define GTHE3_CHANNEL__RX_DFE_KL_LPM_KH_CFG0   	32'h0108	// Type=BINARY; Min=2'b00, Max=2'b11
`define GTHE3_CHANNEL__RX_DFE_KL_LPM_KH_CFG0_SZ	2

`define GTHE3_CHANNEL__RX_DFE_KL_LPM_KH_CFG1   	32'h0109	// Type=BINARY; Min=3'b000, Max=3'b111
`define GTHE3_CHANNEL__RX_DFE_KL_LPM_KH_CFG1_SZ	3

`define GTHE3_CHANNEL__RX_DFE_KL_LPM_KL_CFG0   	32'h010a	// Type=BINARY; Min=2'b00, Max=2'b11
`define GTHE3_CHANNEL__RX_DFE_KL_LPM_KL_CFG0_SZ	2

`define GTHE3_CHANNEL__RX_DFE_KL_LPM_KL_CFG1   	32'h010b	// Type=BINARY; Min=3'b000, Max=3'b111
`define GTHE3_CHANNEL__RX_DFE_KL_LPM_KL_CFG1_SZ	3

`define GTHE3_CHANNEL__RX_DFE_LPM_HOLD_DURING_EIDLE   	32'h010c	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RX_DFE_LPM_HOLD_DURING_EIDLE_SZ	1

`define GTHE3_CHANNEL__RX_DISPERR_SEQ_MATCH   	32'h010d	// Type=STRING; Values=TRUE,FALSE
`define GTHE3_CHANNEL__RX_DISPERR_SEQ_MATCH_SZ	40

`define GTHE3_CHANNEL__RX_DIVRESET_TIME   	32'h010e	// Type=BINARY; Min=5'b00000, Max=5'b11111
`define GTHE3_CHANNEL__RX_DIVRESET_TIME_SZ	5

`define GTHE3_CHANNEL__RX_EN_HI_LR   	32'h010f	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RX_EN_HI_LR_SZ	1

`define GTHE3_CHANNEL__RX_EYESCAN_VS_CODE   	32'h0110	// Type=BINARY; Min=7'b0000000, Max=7'b1111111
`define GTHE3_CHANNEL__RX_EYESCAN_VS_CODE_SZ	7

`define GTHE3_CHANNEL__RX_EYESCAN_VS_NEG_DIR   	32'h0111	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RX_EYESCAN_VS_NEG_DIR_SZ	1

`define GTHE3_CHANNEL__RX_EYESCAN_VS_RANGE   	32'h0112	// Type=BINARY; Min=2'b00, Max=2'b11
`define GTHE3_CHANNEL__RX_EYESCAN_VS_RANGE_SZ	2

`define GTHE3_CHANNEL__RX_EYESCAN_VS_UT_SIGN   	32'h0113	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RX_EYESCAN_VS_UT_SIGN_SZ	1

`define GTHE3_CHANNEL__RX_FABINT_USRCLK_FLOP   	32'h0114	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RX_FABINT_USRCLK_FLOP_SZ	1

`define GTHE3_CHANNEL__RX_INT_DATAWIDTH   	32'h0115	// Type=DECIMAL; Values=1,0,2
`define GTHE3_CHANNEL__RX_INT_DATAWIDTH_SZ	32

`define GTHE3_CHANNEL__RX_PMA_POWER_SAVE   	32'h0116	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RX_PMA_POWER_SAVE_SZ	1

`define GTHE3_CHANNEL__RX_PROGDIV_CFG   	32'h0117	// Type=FLOAT; Values=4.0,5.0,8.0,10.0,16.0,16.5,20.0,32.0,33.0,40.0,64.0,66.0
`define GTHE3_CHANNEL__RX_PROGDIV_CFG_SZ	64

`define GTHE3_CHANNEL__RX_SAMPLE_PERIOD   	32'h0118	// Type=BINARY; Min=3'b000, Max=3'b111
`define GTHE3_CHANNEL__RX_SAMPLE_PERIOD_SZ	3

`define GTHE3_CHANNEL__RX_SIG_VALID_DLY   	32'h0119	// Type=DECIMAL; Values=11,1,2,3,4,5,6,7,8,9,10,12,13,14,15,16,17,18,19,20,21,22,23,24,25,26,27,28,29,30,31,32
`define GTHE3_CHANNEL__RX_SIG_VALID_DLY_SZ	32

`define GTHE3_CHANNEL__RX_SUM_DFETAPREP_EN   	32'h011a	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RX_SUM_DFETAPREP_EN_SZ	1

`define GTHE3_CHANNEL__RX_SUM_IREF_TUNE   	32'h011b	// Type=BINARY; Min=4'b0000, Max=4'b1111
`define GTHE3_CHANNEL__RX_SUM_IREF_TUNE_SZ	4

`define GTHE3_CHANNEL__RX_SUM_RES_CTRL   	32'h011c	// Type=BINARY; Min=2'b00, Max=2'b11
`define GTHE3_CHANNEL__RX_SUM_RES_CTRL_SZ	2

`define GTHE3_CHANNEL__RX_SUM_VCMTUNE   	32'h011d	// Type=BINARY; Min=4'b0000, Max=4'b1111
`define GTHE3_CHANNEL__RX_SUM_VCMTUNE_SZ	4

`define GTHE3_CHANNEL__RX_SUM_VCM_OVWR   	32'h011e	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RX_SUM_VCM_OVWR_SZ	1

`define GTHE3_CHANNEL__RX_SUM_VREF_TUNE   	32'h011f	// Type=BINARY; Min=3'b000, Max=3'b111
`define GTHE3_CHANNEL__RX_SUM_VREF_TUNE_SZ	3

`define GTHE3_CHANNEL__RX_TUNE_AFE_OS   	32'h0120	// Type=BINARY; Min=2'b00, Max=2'b11
`define GTHE3_CHANNEL__RX_TUNE_AFE_OS_SZ	2

`define GTHE3_CHANNEL__RX_WIDEMODE_CDR   	32'h0121	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__RX_WIDEMODE_CDR_SZ	1

`define GTHE3_CHANNEL__RX_XCLK_SEL   	32'h0122	// Type=STRING; Values=RXDES,RXPMA,RXUSR
`define GTHE3_CHANNEL__RX_XCLK_SEL_SZ	40

`define GTHE3_CHANNEL__SAS_MAX_COM   	32'h0123	// Type=DECIMAL; Values=64,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,23,24,25,26,27,28,29,30,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127
`define GTHE3_CHANNEL__SAS_MAX_COM_SZ	32

`define GTHE3_CHANNEL__SAS_MIN_COM   	32'h0124	// Type=DECIMAL; Values=36,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,23,24,25,26,27,28,29,30,31,32,33,34,35,37,38,39,40,41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63
`define GTHE3_CHANNEL__SAS_MIN_COM_SZ	32

`define GTHE3_CHANNEL__SATA_BURST_SEQ_LEN   	32'h0125	// Type=BINARY; Min=4'b0000, Max=4'b1111
`define GTHE3_CHANNEL__SATA_BURST_SEQ_LEN_SZ	4

`define GTHE3_CHANNEL__SATA_BURST_VAL   	32'h0126	// Type=BINARY; Min=3'b000, Max=3'b111
`define GTHE3_CHANNEL__SATA_BURST_VAL_SZ	3

`define GTHE3_CHANNEL__SATA_CPLL_CFG   	32'h0127	// Type=STRING; Values=VCO_3000MHZ,VCO_750MHZ,VCO_1500MHZ
`define GTHE3_CHANNEL__SATA_CPLL_CFG_SZ	88

`define GTHE3_CHANNEL__SATA_EIDLE_VAL   	32'h0128	// Type=BINARY; Min=3'b000, Max=3'b111
`define GTHE3_CHANNEL__SATA_EIDLE_VAL_SZ	3

`define GTHE3_CHANNEL__SATA_MAX_BURST   	32'h0129	// Type=DECIMAL; Values=8,1,2,3,4,5,6,7,9,10,11,12,13,14,15,16,17,18,19,20,21,22,23,24,25,26,27,28,29,30,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63
`define GTHE3_CHANNEL__SATA_MAX_BURST_SZ	32

`define GTHE3_CHANNEL__SATA_MAX_INIT   	32'h012a	// Type=DECIMAL; Values=21,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,22,23,24,25,26,27,28,29,30,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63
`define GTHE3_CHANNEL__SATA_MAX_INIT_SZ	32

`define GTHE3_CHANNEL__SATA_MAX_WAKE   	32'h012b	// Type=DECIMAL; Values=7,1,2,3,4,5,6,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,23,24,25,26,27,28,29,30,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63
`define GTHE3_CHANNEL__SATA_MAX_WAKE_SZ	32

`define GTHE3_CHANNEL__SATA_MIN_BURST   	32'h012c	// Type=DECIMAL; Values=4,1,2,3,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,23,24,25,26,27,28,29,30,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61
`define GTHE3_CHANNEL__SATA_MIN_BURST_SZ	32

`define GTHE3_CHANNEL__SATA_MIN_INIT   	32'h012d	// Type=DECIMAL; Values=12,1,2,3,4,5,6,7,8,9,10,11,13,14,15,16,17,18,19,20,21,22,23,24,25,26,27,28,29,30,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63
`define GTHE3_CHANNEL__SATA_MIN_INIT_SZ	32

`define GTHE3_CHANNEL__SATA_MIN_WAKE   	32'h012e	// Type=DECIMAL; Values=4,1,2,3,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,23,24,25,26,27,28,29,30,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63
`define GTHE3_CHANNEL__SATA_MIN_WAKE_SZ	32

`define GTHE3_CHANNEL__SHOW_REALIGN_COMMA   	32'h012f	// Type=STRING; Values=TRUE,FALSE
`define GTHE3_CHANNEL__SHOW_REALIGN_COMMA_SZ	40

`define GTHE3_CHANNEL__SIM_CPLLREFCLK_SEL   	32'h0130	// Type=BINARY; Min=3'b000, Max=3'b111
`define GTHE3_CHANNEL__SIM_CPLLREFCLK_SEL_SZ	3

`define GTHE3_CHANNEL__SIM_RECEIVER_DETECT_PASS   	32'h0131	// Type=STRING; Values=TRUE,FALSE
`define GTHE3_CHANNEL__SIM_RECEIVER_DETECT_PASS_SZ	40

`define GTHE3_CHANNEL__SIM_RESET_SPEEDUP   	32'h0132	// Type=STRING; Values=TRUE,FALSE
`define GTHE3_CHANNEL__SIM_RESET_SPEEDUP_SZ	40

`define GTHE3_CHANNEL__SIM_TX_EIDLE_DRIVE_LEVEL   	32'h0133	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__SIM_TX_EIDLE_DRIVE_LEVEL_SZ	1

`define GTHE3_CHANNEL__SIM_VERSION   	32'h0134	// Type=STRING; Values=Ver_1,Ver_1_1,Ver_2
`define GTHE3_CHANNEL__SIM_VERSION_SZ	56

`define GTHE3_CHANNEL__TAPDLY_SET_TX   	32'h0135	// Type=HEX; Min=2'h0, Max=2'h3
`define GTHE3_CHANNEL__TAPDLY_SET_TX_SZ	2

`define GTHE3_CHANNEL__TEMPERATUR_PAR   	32'h0136	// Type=BINARY; Min=4'b0000, Max=4'b1111
`define GTHE3_CHANNEL__TEMPERATUR_PAR_SZ	4

`define GTHE3_CHANNEL__TERM_RCAL_CFG   	32'h0137	// Type=BINARY; Min=15'b000000000000000, Max=15'b111111111111111
`define GTHE3_CHANNEL__TERM_RCAL_CFG_SZ	15

`define GTHE3_CHANNEL__TERM_RCAL_OVRD   	32'h0138	// Type=BINARY; Min=3'b000, Max=3'b111
`define GTHE3_CHANNEL__TERM_RCAL_OVRD_SZ	3

`define GTHE3_CHANNEL__TRANS_TIME_RATE   	32'h0139	// Type=HEX; Min=8'h00, Max=8'hff
`define GTHE3_CHANNEL__TRANS_TIME_RATE_SZ	8

`define GTHE3_CHANNEL__TST_RSV0   	32'h013a	// Type=HEX; Min=8'h00, Max=8'hff
`define GTHE3_CHANNEL__TST_RSV0_SZ	8

`define GTHE3_CHANNEL__TST_RSV1   	32'h013b	// Type=HEX; Min=8'h00, Max=8'hff
`define GTHE3_CHANNEL__TST_RSV1_SZ	8

`define GTHE3_CHANNEL__TXBUF_EN   	32'h013c	// Type=STRING; Values=TRUE,FALSE
`define GTHE3_CHANNEL__TXBUF_EN_SZ	40

`define GTHE3_CHANNEL__TXBUF_RESET_ON_RATE_CHANGE   	32'h013d	// Type=STRING; Values=FALSE,TRUE
`define GTHE3_CHANNEL__TXBUF_RESET_ON_RATE_CHANGE_SZ	40

`define GTHE3_CHANNEL__TXDLY_CFG   	32'h013e	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__TXDLY_CFG_SZ	16

`define GTHE3_CHANNEL__TXDLY_LCFG   	32'h013f	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__TXDLY_LCFG_SZ	16

`define GTHE3_CHANNEL__TXDRVBIAS_N   	32'h0140	// Type=BINARY; Min=4'b0000, Max=4'b1111
`define GTHE3_CHANNEL__TXDRVBIAS_N_SZ	4

`define GTHE3_CHANNEL__TXDRVBIAS_P   	32'h0141	// Type=BINARY; Min=4'b0000, Max=4'b1111
`define GTHE3_CHANNEL__TXDRVBIAS_P_SZ	4

`define GTHE3_CHANNEL__TXFIFO_ADDR_CFG   	32'h0142	// Type=STRING; Values=LOW,HIGH
`define GTHE3_CHANNEL__TXFIFO_ADDR_CFG_SZ	32

`define GTHE3_CHANNEL__TXGBOX_FIFO_INIT_RD_ADDR   	32'h0143	// Type=DECIMAL; Values=4,2,3,5,6
`define GTHE3_CHANNEL__TXGBOX_FIFO_INIT_RD_ADDR_SZ	32

`define GTHE3_CHANNEL__TXGEARBOX_EN   	32'h0144	// Type=STRING; Values=FALSE,TRUE
`define GTHE3_CHANNEL__TXGEARBOX_EN_SZ	40

`define GTHE3_CHANNEL__TXOUT_DIV   	32'h0145	// Type=DECIMAL; Values=4,1,2,8,16
`define GTHE3_CHANNEL__TXOUT_DIV_SZ	32

`define GTHE3_CHANNEL__TXPCSRESET_TIME   	32'h0146	// Type=BINARY; Min=5'b00000, Max=5'b11111
`define GTHE3_CHANNEL__TXPCSRESET_TIME_SZ	5

`define GTHE3_CHANNEL__TXPHDLY_CFG0   	32'h0147	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__TXPHDLY_CFG0_SZ	16

`define GTHE3_CHANNEL__TXPHDLY_CFG1   	32'h0148	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__TXPHDLY_CFG1_SZ	16

`define GTHE3_CHANNEL__TXPH_CFG   	32'h0149	// Type=HEX; Min=16'h0000, Max=16'hffff
`define GTHE3_CHANNEL__TXPH_CFG_SZ	16

`define GTHE3_CHANNEL__TXPH_MONITOR_SEL   	32'h014a	// Type=BINARY; Min=5'b00000, Max=5'b11111
`define GTHE3_CHANNEL__TXPH_MONITOR_SEL_SZ	5

`define GTHE3_CHANNEL__TXPI_CFG0   	32'h014b	// Type=BINARY; Min=2'b00, Max=2'b11
`define GTHE3_CHANNEL__TXPI_CFG0_SZ	2

`define GTHE3_CHANNEL__TXPI_CFG1   	32'h014c	// Type=BINARY; Min=2'b00, Max=2'b11
`define GTHE3_CHANNEL__TXPI_CFG1_SZ	2

`define GTHE3_CHANNEL__TXPI_CFG2   	32'h014d	// Type=BINARY; Min=2'b00, Max=2'b11
`define GTHE3_CHANNEL__TXPI_CFG2_SZ	2

`define GTHE3_CHANNEL__TXPI_CFG3   	32'h014e	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__TXPI_CFG3_SZ	1

`define GTHE3_CHANNEL__TXPI_CFG4   	32'h014f	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__TXPI_CFG4_SZ	1

`define GTHE3_CHANNEL__TXPI_CFG5   	32'h0150	// Type=BINARY; Min=3'b000, Max=3'b111
`define GTHE3_CHANNEL__TXPI_CFG5_SZ	3

`define GTHE3_CHANNEL__TXPI_GRAY_SEL   	32'h0151	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__TXPI_GRAY_SEL_SZ	1

`define GTHE3_CHANNEL__TXPI_INVSTROBE_SEL   	32'h0152	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__TXPI_INVSTROBE_SEL_SZ	1

`define GTHE3_CHANNEL__TXPI_LPM   	32'h0153	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__TXPI_LPM_SZ	1

`define GTHE3_CHANNEL__TXPI_PPMCLK_SEL   	32'h0154	// Type=STRING; Values=TXUSRCLK2,TXUSRCLK
`define GTHE3_CHANNEL__TXPI_PPMCLK_SEL_SZ	72

`define GTHE3_CHANNEL__TXPI_PPM_CFG   	32'h0155	// Type=BINARY; Min=8'b00000000, Max=8'b11111111
`define GTHE3_CHANNEL__TXPI_PPM_CFG_SZ	8

`define GTHE3_CHANNEL__TXPI_SYNFREQ_PPM   	32'h0156	// Type=BINARY; Min=3'b000, Max=3'b111
`define GTHE3_CHANNEL__TXPI_SYNFREQ_PPM_SZ	3

`define GTHE3_CHANNEL__TXPI_VREFSEL   	32'h0157	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__TXPI_VREFSEL_SZ	1

`define GTHE3_CHANNEL__TXPMARESET_TIME   	32'h0158	// Type=BINARY; Min=5'b00000, Max=5'b11111
`define GTHE3_CHANNEL__TXPMARESET_TIME_SZ	5

`define GTHE3_CHANNEL__TXSYNC_MULTILANE   	32'h0159	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__TXSYNC_MULTILANE_SZ	1

`define GTHE3_CHANNEL__TXSYNC_OVRD   	32'h015a	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__TXSYNC_OVRD_SZ	1

`define GTHE3_CHANNEL__TXSYNC_SKIP_DA   	32'h015b	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__TXSYNC_SKIP_DA_SZ	1

`define GTHE3_CHANNEL__TX_CLK25_DIV   	32'h015c	// Type=DECIMAL; Values=8,1,2,3,4,5,6,7,9,10,11,12,13,14,15,16,17,18,19,20,21,22,23,24,25,26,27,28,29,30,31,32
`define GTHE3_CHANNEL__TX_CLK25_DIV_SZ	32

`define GTHE3_CHANNEL__TX_CLKMUX_EN   	32'h015d	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__TX_CLKMUX_EN_SZ	1

`define GTHE3_CHANNEL__TX_DATA_WIDTH   	32'h015e	// Type=DECIMAL; Values=20,16,32,40,64,80,128,160
`define GTHE3_CHANNEL__TX_DATA_WIDTH_SZ	32

`define GTHE3_CHANNEL__TX_DCD_CFG   	32'h015f	// Type=BINARY; Min=6'b000000, Max=6'b111111
`define GTHE3_CHANNEL__TX_DCD_CFG_SZ	6

`define GTHE3_CHANNEL__TX_DCD_EN   	32'h0160	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__TX_DCD_EN_SZ	1

`define GTHE3_CHANNEL__TX_DEEMPH0   	32'h0161	// Type=BINARY; Min=6'b000000, Max=6'b111111
`define GTHE3_CHANNEL__TX_DEEMPH0_SZ	6

`define GTHE3_CHANNEL__TX_DEEMPH1   	32'h0162	// Type=BINARY; Min=6'b000000, Max=6'b111111
`define GTHE3_CHANNEL__TX_DEEMPH1_SZ	6

`define GTHE3_CHANNEL__TX_DIVRESET_TIME   	32'h0163	// Type=BINARY; Min=5'b00000, Max=5'b11111
`define GTHE3_CHANNEL__TX_DIVRESET_TIME_SZ	5

`define GTHE3_CHANNEL__TX_DRIVE_MODE   	32'h0164	// Type=STRING; Values=DIRECT,PIPE,PIPEGEN3
`define GTHE3_CHANNEL__TX_DRIVE_MODE_SZ	64

`define GTHE3_CHANNEL__TX_EIDLE_ASSERT_DELAY   	32'h0165	// Type=BINARY; Min=3'b000, Max=3'b111
`define GTHE3_CHANNEL__TX_EIDLE_ASSERT_DELAY_SZ	3

`define GTHE3_CHANNEL__TX_EIDLE_DEASSERT_DELAY   	32'h0166	// Type=BINARY; Min=3'b000, Max=3'b111
`define GTHE3_CHANNEL__TX_EIDLE_DEASSERT_DELAY_SZ	3

`define GTHE3_CHANNEL__TX_EML_PHI_TUNE   	32'h0167	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__TX_EML_PHI_TUNE_SZ	1

`define GTHE3_CHANNEL__TX_FABINT_USRCLK_FLOP   	32'h0168	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__TX_FABINT_USRCLK_FLOP_SZ	1

`define GTHE3_CHANNEL__TX_IDLE_DATA_ZERO   	32'h0169	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__TX_IDLE_DATA_ZERO_SZ	1

`define GTHE3_CHANNEL__TX_INT_DATAWIDTH   	32'h016a	// Type=DECIMAL; Values=1,0,2
`define GTHE3_CHANNEL__TX_INT_DATAWIDTH_SZ	32

`define GTHE3_CHANNEL__TX_LOOPBACK_DRIVE_HIZ   	32'h016b	// Type=STRING; Values=FALSE,TRUE
`define GTHE3_CHANNEL__TX_LOOPBACK_DRIVE_HIZ_SZ	40

`define GTHE3_CHANNEL__TX_MAINCURSOR_SEL   	32'h016c	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__TX_MAINCURSOR_SEL_SZ	1

`define GTHE3_CHANNEL__TX_MARGIN_FULL_0   	32'h016d	// Type=BINARY; Min=7'b0000000, Max=7'b1111111
`define GTHE3_CHANNEL__TX_MARGIN_FULL_0_SZ	7

`define GTHE3_CHANNEL__TX_MARGIN_FULL_1   	32'h016e	// Type=BINARY; Min=7'b0000000, Max=7'b1111111
`define GTHE3_CHANNEL__TX_MARGIN_FULL_1_SZ	7

`define GTHE3_CHANNEL__TX_MARGIN_FULL_2   	32'h016f	// Type=BINARY; Min=7'b0000000, Max=7'b1111111
`define GTHE3_CHANNEL__TX_MARGIN_FULL_2_SZ	7

`define GTHE3_CHANNEL__TX_MARGIN_FULL_3   	32'h0170	// Type=BINARY; Min=7'b0000000, Max=7'b1111111
`define GTHE3_CHANNEL__TX_MARGIN_FULL_3_SZ	7

`define GTHE3_CHANNEL__TX_MARGIN_FULL_4   	32'h0171	// Type=BINARY; Min=7'b0000000, Max=7'b1111111
`define GTHE3_CHANNEL__TX_MARGIN_FULL_4_SZ	7

`define GTHE3_CHANNEL__TX_MARGIN_LOW_0   	32'h0172	// Type=BINARY; Min=7'b0000000, Max=7'b1111111
`define GTHE3_CHANNEL__TX_MARGIN_LOW_0_SZ	7

`define GTHE3_CHANNEL__TX_MARGIN_LOW_1   	32'h0173	// Type=BINARY; Min=7'b0000000, Max=7'b1111111
`define GTHE3_CHANNEL__TX_MARGIN_LOW_1_SZ	7

`define GTHE3_CHANNEL__TX_MARGIN_LOW_2   	32'h0174	// Type=BINARY; Min=7'b0000000, Max=7'b1111111
`define GTHE3_CHANNEL__TX_MARGIN_LOW_2_SZ	7

`define GTHE3_CHANNEL__TX_MARGIN_LOW_3   	32'h0175	// Type=BINARY; Min=7'b0000000, Max=7'b1111111
`define GTHE3_CHANNEL__TX_MARGIN_LOW_3_SZ	7

`define GTHE3_CHANNEL__TX_MARGIN_LOW_4   	32'h0176	// Type=BINARY; Min=7'b0000000, Max=7'b1111111
`define GTHE3_CHANNEL__TX_MARGIN_LOW_4_SZ	7

`define GTHE3_CHANNEL__TX_MODE_SEL   	32'h0177	// Type=BINARY; Min=3'b000, Max=3'b111
`define GTHE3_CHANNEL__TX_MODE_SEL_SZ	3

`define GTHE3_CHANNEL__TX_PMADATA_OPT   	32'h0178	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__TX_PMADATA_OPT_SZ	1

`define GTHE3_CHANNEL__TX_PMA_POWER_SAVE   	32'h0179	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__TX_PMA_POWER_SAVE_SZ	1

`define GTHE3_CHANNEL__TX_PROGCLK_SEL   	32'h017a	// Type=STRING; Values=POSTPI,CPLL,PREPI
`define GTHE3_CHANNEL__TX_PROGCLK_SEL_SZ	48

`define GTHE3_CHANNEL__TX_PROGDIV_CFG   	32'h017b	// Type=FLOAT; Values=4.0,5.0,8.0,10.0,16.0,16.5,20.0,32.0,33.0,40.0,64.0,66.0
`define GTHE3_CHANNEL__TX_PROGDIV_CFG_SZ	64

`define GTHE3_CHANNEL__TX_QPI_STATUS_EN   	32'h017c	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__TX_QPI_STATUS_EN_SZ	1

`define GTHE3_CHANNEL__TX_RXDETECT_CFG   	32'h017d	// Type=HEX; Min=14'h0000, Max=14'h3fff
`define GTHE3_CHANNEL__TX_RXDETECT_CFG_SZ	14

`define GTHE3_CHANNEL__TX_RXDETECT_REF   	32'h017e	// Type=BINARY; Min=3'b000, Max=3'b111
`define GTHE3_CHANNEL__TX_RXDETECT_REF_SZ	3

`define GTHE3_CHANNEL__TX_SAMPLE_PERIOD   	32'h017f	// Type=BINARY; Min=3'b000, Max=3'b111
`define GTHE3_CHANNEL__TX_SAMPLE_PERIOD_SZ	3

`define GTHE3_CHANNEL__TX_SARC_LPBK_ENB   	32'h0180	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__TX_SARC_LPBK_ENB_SZ	1

`define GTHE3_CHANNEL__TX_XCLK_SEL   	32'h0181	// Type=STRING; Values=TXOUT,TXUSR
`define GTHE3_CHANNEL__TX_XCLK_SEL_SZ	40

`define GTHE3_CHANNEL__USE_PCS_CLK_PHASE_SEL   	32'h0182	// Type=BINARY; Min=1'b0, Max=1'b1
`define GTHE3_CHANNEL__USE_PCS_CLK_PHASE_SEL_SZ	1

`define GTHE3_CHANNEL__WB_MODE   	32'h0183	// Type=BINARY; Min=2'b00, Max=2'b11
`define GTHE3_CHANNEL__WB_MODE_SZ	2

`endif  // B_GTHE3_CHANNEL_DEFINES_VH
