`include "B_ODELAYE3_defines.vh"

reg [`ODELAYE3_DATA_SZ-1:0] ATTR [0:`ODELAYE3_ADDR_N-1];
reg [96:1] CASCADE_REG = CASCADE;
reg [40:1] DELAY_FORMAT_REG = DELAY_FORMAT;
reg [64:1] DELAY_TYPE_REG = DELAY_TYPE;
reg [10:0] DELAY_VALUE_REG = DELAY_VALUE;
reg IS_CLK_INVERTED_REG = IS_CLK_INVERTED;
reg IS_RST_INVERTED_REG = IS_RST_INVERTED;
real REFCLK_FREQUENCY_REG = REFCLK_FREQUENCY;
real SIM_VERSION_REG = SIM_VERSION;
reg [48:1] UPDATE_MODE_REG = UPDATE_MODE;

initial begin
ATTR[`ODELAYE3__CASCADE] = CASCADE;
ATTR[`ODELAYE3__DELAY_FORMAT] = DELAY_FORMAT;
ATTR[`ODELAYE3__DELAY_TYPE] = DELAY_TYPE;
ATTR[`ODELAYE3__DELAY_VALUE] = DELAY_VALUE;
ATTR[`ODELAYE3__IS_CLK_INVERTED] = IS_CLK_INVERTED;
ATTR[`ODELAYE3__IS_RST_INVERTED] = IS_RST_INVERTED;
ATTR[`ODELAYE3__REFCLK_FREQUENCY] = $realtobits(REFCLK_FREQUENCY);
ATTR[`ODELAYE3__SIM_VERSION] = $realtobits(SIM_VERSION);
ATTR[`ODELAYE3__UPDATE_MODE] = UPDATE_MODE;
end

always @(trig_attr) begin
CASCADE_REG = ATTR[`ODELAYE3__CASCADE];
DELAY_FORMAT_REG = ATTR[`ODELAYE3__DELAY_FORMAT];
DELAY_TYPE_REG = ATTR[`ODELAYE3__DELAY_TYPE];
DELAY_VALUE_REG = ATTR[`ODELAYE3__DELAY_VALUE];
IS_CLK_INVERTED_REG = ATTR[`ODELAYE3__IS_CLK_INVERTED];
IS_RST_INVERTED_REG = ATTR[`ODELAYE3__IS_RST_INVERTED];
REFCLK_FREQUENCY_REG = $bitstoreal(ATTR[`ODELAYE3__REFCLK_FREQUENCY]);
SIM_VERSION_REG = $bitstoreal(ATTR[`ODELAYE3__SIM_VERSION]);
UPDATE_MODE_REG = ATTR[`ODELAYE3__UPDATE_MODE];
end

// procedures to override, read attribute values

task write_attr;
  input  [`ODELAYE3_ADDR_SZ-1:0] addr;
  input  [`ODELAYE3_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`ODELAYE3_DATA_SZ-1:0] read_attr;
  input  [`ODELAYE3_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
    trig_attr = ~trig_attr;
  end
endtask
