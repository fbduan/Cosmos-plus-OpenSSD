// BLH dynamic attribute configuration look-up table addresses
//
// Build Summary:
//    Built By:     mk_defines_vh 3.0001
//    Built On:     Wed May 21 17:07:22 2014
//    Bundle:       XIPHY
//    Architecture: olympus
//    Snapshot Dir: /tmp/MgzBFkdK57
// Environment Variables:
//    XILENV="/build/xfndry/HEAD/env"
//    MYXILENV=""
//

`ifdef B_RXTX_BITSLICE_DEFINES_VH
`else
`define B_RXTX_BITSLICE_DEFINES_VH

// Look-up table parameters
//

`define RXTX_BITSLICE_ADDR_N  27
`define RXTX_BITSLICE_ADDR_SZ 32
`define RXTX_BITSLICE_DATA_SZ 112

// Attribute addresses
//

`define RXTX_BITSLICE__ENABLE_PRE_EMPHASIS   	32'h0000	// Type=BOOLSTRING; Values=FALSE,TRUE
`define RXTX_BITSLICE__ENABLE_PRE_EMPHASIS_SZ	40

`define RXTX_BITSLICE__FIFO_SYNC_MODE   	32'h0001	// Type=BOOLSTRING; Values=FALSE,TRUE
`define RXTX_BITSLICE__FIFO_SYNC_MODE_SZ	40

`define RXTX_BITSLICE__INIT   	32'h0002	// Type=BINARY; Values=1'b1,1'b0
`define RXTX_BITSLICE__INIT_SZ	1

`define RXTX_BITSLICE__IS_RX_CLK_INVERTED   	32'h0003	// Type=BINARY; Min=1'b0, Max=1'b1
`define RXTX_BITSLICE__IS_RX_CLK_INVERTED_SZ	1

`define RXTX_BITSLICE__IS_RX_RST_DLY_INVERTED   	32'h0004	// Type=BINARY; Min=1'b0, Max=1'b1
`define RXTX_BITSLICE__IS_RX_RST_DLY_INVERTED_SZ	1

`define RXTX_BITSLICE__IS_RX_RST_INVERTED   	32'h0005	// Type=BINARY; Min=1'b0, Max=1'b1
`define RXTX_BITSLICE__IS_RX_RST_INVERTED_SZ	1

`define RXTX_BITSLICE__IS_TX_CLK_INVERTED   	32'h0006	// Type=BINARY; Min=1'b0, Max=1'b1
`define RXTX_BITSLICE__IS_TX_CLK_INVERTED_SZ	1

`define RXTX_BITSLICE__IS_TX_RST_DLY_INVERTED   	32'h0007	// Type=BINARY; Min=1'b0, Max=1'b1
`define RXTX_BITSLICE__IS_TX_RST_DLY_INVERTED_SZ	1

`define RXTX_BITSLICE__IS_TX_RST_INVERTED   	32'h0008	// Type=BINARY; Min=1'b0, Max=1'b1
`define RXTX_BITSLICE__IS_TX_RST_INVERTED_SZ	1

`define RXTX_BITSLICE__LOOPBACK   	32'h0009	// Type=BOOLSTRING; Values=FALSE,TRUE
`define RXTX_BITSLICE__LOOPBACK_SZ	40

`define RXTX_BITSLICE__NATIVE_ODELAY_BYPASS   	32'h000a	// Type=BOOLSTRING; Values=FALSE,TRUE
`define RXTX_BITSLICE__NATIVE_ODELAY_BYPASS_SZ	40

`define RXTX_BITSLICE__RX_DATA_TYPE   	32'h000b	// Type=STRING; Values=NONE,CLOCK,DATA,DATA_AND_CLOCK
`define RXTX_BITSLICE__RX_DATA_TYPE_SZ	112

`define RXTX_BITSLICE__RX_DATA_WIDTH   	32'h000c	// Type=DECIMAL; Values=8,4
`define RXTX_BITSLICE__RX_DATA_WIDTH_SZ	32

`define RXTX_BITSLICE__RX_DELAY_FORMAT   	32'h000d	// Type=STRING; Values=TIME,COUNT
`define RXTX_BITSLICE__RX_DELAY_FORMAT_SZ	40

`define RXTX_BITSLICE__RX_DELAY_TYPE   	32'h000e	// Type=STRING; Values=FIXED,VAR_LOAD,VARIABLE
`define RXTX_BITSLICE__RX_DELAY_TYPE_SZ	64

`define RXTX_BITSLICE__RX_DELAY_VALUE   	32'h000f	// Type=DECIMAL; Min=0, Max=1250
`define RXTX_BITSLICE__RX_DELAY_VALUE_SZ	32

`define RXTX_BITSLICE__RX_REFCLK_FREQUENCY   	32'h0010	// Type=FLOAT; Min=200.0, Max=2400.0
`define RXTX_BITSLICE__RX_REFCLK_FREQUENCY_SZ	64

`define RXTX_BITSLICE__RX_UPDATE_MODE   	32'h0011	// Type=STRING; Values=ASYNC,MANUAL,SYNC
`define RXTX_BITSLICE__RX_UPDATE_MODE_SZ	48

`define RXTX_BITSLICE__SIM_VERSION   	32'h0012	// Type=FLOAT; Values=2.0,1.0
`define RXTX_BITSLICE__SIM_VERSION_SZ	64

`define RXTX_BITSLICE__TBYTE_CTL   	32'h0013	// Type=STRING; Values=TBYTE_IN,T
`define RXTX_BITSLICE__TBYTE_CTL_SZ	64

`define RXTX_BITSLICE__TX_DATA_WIDTH   	32'h0014	// Type=DECIMAL; Values=8,4
`define RXTX_BITSLICE__TX_DATA_WIDTH_SZ	32

`define RXTX_BITSLICE__TX_DELAY_FORMAT   	32'h0015	// Type=STRING; Values=TIME,COUNT
`define RXTX_BITSLICE__TX_DELAY_FORMAT_SZ	40

`define RXTX_BITSLICE__TX_DELAY_TYPE   	32'h0016	// Type=STRING; Values=FIXED,VAR_LOAD,VARIABLE
`define RXTX_BITSLICE__TX_DELAY_TYPE_SZ	64

`define RXTX_BITSLICE__TX_DELAY_VALUE   	32'h0017	// Type=DECIMAL; Min=0, Max=1250
`define RXTX_BITSLICE__TX_DELAY_VALUE_SZ	32

`define RXTX_BITSLICE__TX_OUTPUT_PHASE_90   	32'h0018	// Type=BOOLSTRING; Values=FALSE,TRUE
`define RXTX_BITSLICE__TX_OUTPUT_PHASE_90_SZ	40

`define RXTX_BITSLICE__TX_REFCLK_FREQUENCY   	32'h0019	// Type=FLOAT; Min=200.0, Max=2400.0
`define RXTX_BITSLICE__TX_REFCLK_FREQUENCY_SZ	64

`define RXTX_BITSLICE__TX_UPDATE_MODE   	32'h001a	// Type=STRING; Values=ASYNC,MANUAL,SYNC
`define RXTX_BITSLICE__TX_UPDATE_MODE_SZ	48

`endif  // B_RXTX_BITSLICE_DEFINES_VH
