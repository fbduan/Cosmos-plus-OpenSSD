// BLH dynamic attribute configuration look-up table addresses
//
// Build Summary:
//    Built By:     mk_defines_vh 3.0001
//    Built On:     Wed Apr 17 17:24:09 2013
//    Bundle:       DSP48E2
//    Architecture: olympus
//    Snapshot Dir: /tmp/H238lm9sMS
// Environment Variables:
//    XILENV="/build/xfndry/HEAD/env"
//    MYXILENV=""
//

`ifdef B_DSP48E2_DEFINES_VH
`else
`define B_DSP48E2_DEFINES_VH

// Look-up table parameters
//

`define DSP48E2_ADDR_N  46
`define DSP48E2_ADDR_SZ 32
`define DSP48E2_DATA_SZ 120

// Attribute addresses
//

`define DSP48E2__ACASCREG   	32'h0000	// Type=DECIMAL; Values=1,0,2
`define DSP48E2__ACASCREG_SZ	32

`define DSP48E2__ADREG   	32'h0001	// Type=DECIMAL; Values=1,0
`define DSP48E2__ADREG_SZ	32

`define DSP48E2__ALUMODEREG   	32'h0002	// Type=DECIMAL; Values=1,0
`define DSP48E2__ALUMODEREG_SZ	32

`define DSP48E2__AMULTSEL   	32'h0003	// Type=STRING; Values=A,AD
`define DSP48E2__AMULTSEL_SZ	16

`define DSP48E2__AREG   	32'h0004	// Type=DECIMAL; Values=1,0,2
`define DSP48E2__AREG_SZ	32

`define DSP48E2__AUTORESET_PATDET   	32'h0005	// Type=STRING; Values=NO_RESET,RESET_MATCH,RESET_NOT_MATCH
`define DSP48E2__AUTORESET_PATDET_SZ	120

`define DSP48E2__AUTORESET_PRIORITY   	32'h0006	// Type=STRING; Values=RESET,CEP
`define DSP48E2__AUTORESET_PRIORITY_SZ	40

`define DSP48E2__A_INPUT   	32'h0007	// Type=STRING; Values=DIRECT,CASCADE
`define DSP48E2__A_INPUT_SZ	56

`define DSP48E2__BCASCREG   	32'h0008	// Type=DECIMAL; Values=1,0,2
`define DSP48E2__BCASCREG_SZ	32

`define DSP48E2__BMULTSEL   	32'h0009	// Type=STRING; Values=B,AD
`define DSP48E2__BMULTSEL_SZ	16

`define DSP48E2__BREG   	32'h000a	// Type=DECIMAL; Values=1,0,2
`define DSP48E2__BREG_SZ	32

`define DSP48E2__B_INPUT   	32'h000b	// Type=STRING; Values=DIRECT,CASCADE
`define DSP48E2__B_INPUT_SZ	56

`define DSP48E2__CARRYINREG   	32'h000c	// Type=DECIMAL; Values=1,0
`define DSP48E2__CARRYINREG_SZ	32

`define DSP48E2__CARRYINSELREG   	32'h000d	// Type=DECIMAL; Values=1,0
`define DSP48E2__CARRYINSELREG_SZ	32

`define DSP48E2__CREG   	32'h000e	// Type=DECIMAL; Values=1,0
`define DSP48E2__CREG_SZ	32

`define DSP48E2__DREG   	32'h000f	// Type=DECIMAL; Values=1,0
`define DSP48E2__DREG_SZ	32

`define DSP48E2__INMODEREG   	32'h0010	// Type=DECIMAL; Values=1,0
`define DSP48E2__INMODEREG_SZ	32

`define DSP48E2__IS_ALUMODE_INVERTED   	32'h0011	// Type=BINARY; Min=4'b0000, Max=4'b1111
`define DSP48E2__IS_ALUMODE_INVERTED_SZ	4

`define DSP48E2__IS_CARRYIN_INVERTED   	32'h0012	// Type=BINARY; Min=1'b0, Max=1'b1
`define DSP48E2__IS_CARRYIN_INVERTED_SZ	1

`define DSP48E2__IS_CLK_INVERTED   	32'h0013	// Type=BINARY; Min=1'b0, Max=1'b1
`define DSP48E2__IS_CLK_INVERTED_SZ	1

`define DSP48E2__IS_INMODE_INVERTED   	32'h0014	// Type=BINARY; Min=5'b00000, Max=5'b11111
`define DSP48E2__IS_INMODE_INVERTED_SZ	5

`define DSP48E2__IS_OPMODE_INVERTED   	32'h0015	// Type=BINARY; Min=9'b000000000, Max=9'b111111111
`define DSP48E2__IS_OPMODE_INVERTED_SZ	9

`define DSP48E2__IS_RSTALLCARRYIN_INVERTED   	32'h0016	// Type=BINARY; Min=1'b0, Max=1'b1
`define DSP48E2__IS_RSTALLCARRYIN_INVERTED_SZ	1

`define DSP48E2__IS_RSTALUMODE_INVERTED   	32'h0017	// Type=BINARY; Min=1'b0, Max=1'b1
`define DSP48E2__IS_RSTALUMODE_INVERTED_SZ	1

`define DSP48E2__IS_RSTA_INVERTED   	32'h0018	// Type=BINARY; Min=1'b0, Max=1'b1
`define DSP48E2__IS_RSTA_INVERTED_SZ	1

`define DSP48E2__IS_RSTB_INVERTED   	32'h0019	// Type=BINARY; Min=1'b0, Max=1'b1
`define DSP48E2__IS_RSTB_INVERTED_SZ	1

`define DSP48E2__IS_RSTCTRL_INVERTED   	32'h001a	// Type=BINARY; Min=1'b0, Max=1'b1
`define DSP48E2__IS_RSTCTRL_INVERTED_SZ	1

`define DSP48E2__IS_RSTC_INVERTED   	32'h001b	// Type=BINARY; Min=1'b0, Max=1'b1
`define DSP48E2__IS_RSTC_INVERTED_SZ	1

`define DSP48E2__IS_RSTD_INVERTED   	32'h001c	// Type=BINARY; Min=1'b0, Max=1'b1
`define DSP48E2__IS_RSTD_INVERTED_SZ	1

`define DSP48E2__IS_RSTINMODE_INVERTED   	32'h001d	// Type=BINARY; Min=1'b0, Max=1'b1
`define DSP48E2__IS_RSTINMODE_INVERTED_SZ	1

`define DSP48E2__IS_RSTM_INVERTED   	32'h001e	// Type=BINARY; Min=1'b0, Max=1'b1
`define DSP48E2__IS_RSTM_INVERTED_SZ	1

`define DSP48E2__IS_RSTP_INVERTED   	32'h001f	// Type=BINARY; Min=1'b0, Max=1'b1
`define DSP48E2__IS_RSTP_INVERTED_SZ	1

`define DSP48E2__MASK   	32'h0020	// Type=HEX; Min=48'h000000000000, Max=48'hffffffffffff
`define DSP48E2__MASK_SZ	48

`define DSP48E2__MREG   	32'h0021	// Type=DECIMAL; Values=1,0
`define DSP48E2__MREG_SZ	32

`define DSP48E2__OPMODEREG   	32'h0022	// Type=DECIMAL; Values=1,0
`define DSP48E2__OPMODEREG_SZ	32

`define DSP48E2__PATTERN   	32'h0023	// Type=HEX; Min=48'h000000000000, Max=48'hffffffffffff
`define DSP48E2__PATTERN_SZ	48

`define DSP48E2__PREADDINSEL   	32'h0024	// Type=STRING; Values=A,B
`define DSP48E2__PREADDINSEL_SZ	8

`define DSP48E2__PREG   	32'h0025	// Type=DECIMAL; Values=1,0
`define DSP48E2__PREG_SZ	32

`define DSP48E2__RND   	32'h0026	// Type=HEX; Min=48'h000000000000, Max=48'hffffffffffff
`define DSP48E2__RND_SZ	48

`define DSP48E2__SEL_MASK   	32'h0027	// Type=STRING; Values=MASK,C,ROUNDING_MODE1,ROUNDING_MODE2
`define DSP48E2__SEL_MASK_SZ	112

`define DSP48E2__SEL_PATTERN   	32'h0028	// Type=STRING; Values=PATTERN,C
`define DSP48E2__SEL_PATTERN_SZ	56

`define DSP48E2__USE_MULT   	32'h0029	// Type=STRING; Values=MULTIPLY,DYNAMIC,NONE
`define DSP48E2__USE_MULT_SZ	64

`define DSP48E2__USE_PATTERN_DETECT   	32'h002a	// Type=STRING; Values=NO_PATDET,PATDET
`define DSP48E2__USE_PATTERN_DETECT_SZ	72

`define DSP48E2__USE_SIMD   	32'h002b	// Type=STRING; Values=ONE48,FOUR12,TWO24
`define DSP48E2__USE_SIMD_SZ	48

`define DSP48E2__USE_WIDEXOR   	32'h002c	// Type=BOOLSTRING; Values=FALSE,TRUE
`define DSP48E2__USE_WIDEXOR_SZ	40

`define DSP48E2__XORSIMD   	32'h002d	// Type=STRING; Values=XOR24_48_96,XOR12
`define DSP48E2__XORSIMD_SZ	88

`endif  // B_DSP48E2_DEFINES_VH
