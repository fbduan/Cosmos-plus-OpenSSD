// BLH dynamic attribute configuration look-up table addresses
//
// Build Summary:
//    Built By:     mk_defines_vh 3.0001
//    Built On:     Wed Apr 17 17:29:28 2013
//    Bundle:       SYSMONE1
//    Architecture: olympus
//    Snapshot Dir: /tmp/6Y_m6JBBaV
// Environment Variables:
//    XILENV="/build/xfndry/HEAD/env"
//    MYXILENV=""
//

`ifdef B_SYSMONE1_DEFINES_VH
`else
`define B_SYSMONE1_DEFINES_VH

// Look-up table parameters
//

`define SYSMONE1_ADDR_N  66
`define SYSMONE1_ADDR_SZ 32
`define SYSMONE1_DATA_SZ 16

// Attribute addresses
//

`define SYSMONE1__INIT_40   	32'h0000	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_40_SZ	16

`define SYSMONE1__INIT_41   	32'h0001	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_41_SZ	16

`define SYSMONE1__INIT_42   	32'h0002	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_42_SZ	16

`define SYSMONE1__INIT_43   	32'h0003	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_43_SZ	16

`define SYSMONE1__INIT_44   	32'h0004	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_44_SZ	16

`define SYSMONE1__INIT_45   	32'h0005	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_45_SZ	16

`define SYSMONE1__INIT_46   	32'h0006	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_46_SZ	16

`define SYSMONE1__INIT_47   	32'h0007	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_47_SZ	16

`define SYSMONE1__INIT_48   	32'h0008	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_48_SZ	16

`define SYSMONE1__INIT_49   	32'h0009	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_49_SZ	16

`define SYSMONE1__INIT_4A   	32'h000a	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_4A_SZ	16

`define SYSMONE1__INIT_4B   	32'h000b	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_4B_SZ	16

`define SYSMONE1__INIT_4C   	32'h000c	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_4C_SZ	16

`define SYSMONE1__INIT_4D   	32'h000d	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_4D_SZ	16

`define SYSMONE1__INIT_4E   	32'h000e	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_4E_SZ	16

`define SYSMONE1__INIT_4F   	32'h000f	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_4F_SZ	16

`define SYSMONE1__INIT_50   	32'h0010	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_50_SZ	16

`define SYSMONE1__INIT_51   	32'h0011	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_51_SZ	16

`define SYSMONE1__INIT_52   	32'h0012	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_52_SZ	16

`define SYSMONE1__INIT_53   	32'h0013	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_53_SZ	16

`define SYSMONE1__INIT_54   	32'h0014	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_54_SZ	16

`define SYSMONE1__INIT_55   	32'h0015	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_55_SZ	16

`define SYSMONE1__INIT_56   	32'h0016	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_56_SZ	16

`define SYSMONE1__INIT_57   	32'h0017	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_57_SZ	16

`define SYSMONE1__INIT_58   	32'h0018	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_58_SZ	16

`define SYSMONE1__INIT_59   	32'h0019	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_59_SZ	16

`define SYSMONE1__INIT_5A   	32'h001a	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_5A_SZ	16

`define SYSMONE1__INIT_5B   	32'h001b	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_5B_SZ	16

`define SYSMONE1__INIT_5C   	32'h001c	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_5C_SZ	16

`define SYSMONE1__INIT_5D   	32'h001d	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_5D_SZ	16

`define SYSMONE1__INIT_5E   	32'h001e	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_5E_SZ	16

`define SYSMONE1__INIT_5F   	32'h001f	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_5F_SZ	16

`define SYSMONE1__INIT_60   	32'h0020	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_60_SZ	16

`define SYSMONE1__INIT_61   	32'h0021	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_61_SZ	16

`define SYSMONE1__INIT_62   	32'h0022	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_62_SZ	16

`define SYSMONE1__INIT_63   	32'h0023	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_63_SZ	16

`define SYSMONE1__INIT_64   	32'h0024	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_64_SZ	16

`define SYSMONE1__INIT_65   	32'h0025	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_65_SZ	16

`define SYSMONE1__INIT_66   	32'h0026	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_66_SZ	16

`define SYSMONE1__INIT_67   	32'h0027	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_67_SZ	16

`define SYSMONE1__INIT_68   	32'h0028	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_68_SZ	16

`define SYSMONE1__INIT_69   	32'h0029	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_69_SZ	16

`define SYSMONE1__INIT_6A   	32'h002a	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_6A_SZ	16

`define SYSMONE1__INIT_6B   	32'h002b	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_6B_SZ	16

`define SYSMONE1__INIT_6C   	32'h002c	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_6C_SZ	16

`define SYSMONE1__INIT_6D   	32'h002d	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_6D_SZ	16

`define SYSMONE1__INIT_6E   	32'h002e	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_6E_SZ	16

`define SYSMONE1__INIT_6F   	32'h002f	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_6F_SZ	16

`define SYSMONE1__INIT_70   	32'h0030	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_70_SZ	16

`define SYSMONE1__INIT_71   	32'h0031	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_71_SZ	16

`define SYSMONE1__INIT_72   	32'h0032	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_72_SZ	16

`define SYSMONE1__INIT_73   	32'h0033	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_73_SZ	16

`define SYSMONE1__INIT_74   	32'h0034	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_74_SZ	16

`define SYSMONE1__INIT_75   	32'h0035	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_75_SZ	16

`define SYSMONE1__INIT_76   	32'h0036	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_76_SZ	16

`define SYSMONE1__INIT_77   	32'h0037	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_77_SZ	16

`define SYSMONE1__INIT_78   	32'h0038	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_78_SZ	16

`define SYSMONE1__INIT_79   	32'h0039	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_79_SZ	16

`define SYSMONE1__INIT_7A   	32'h003a	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_7A_SZ	16

`define SYSMONE1__INIT_7B   	32'h003b	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_7B_SZ	16

`define SYSMONE1__INIT_7C   	32'h003c	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_7C_SZ	16

`define SYSMONE1__INIT_7D   	32'h003d	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_7D_SZ	16

`define SYSMONE1__INIT_7E   	32'h003e	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_7E_SZ	16

`define SYSMONE1__INIT_7F   	32'h003f	// Type=HEX; Min=16'h0000, Max=16'hffff
`define SYSMONE1__INIT_7F_SZ	16

`define SYSMONE1__IS_CONVSTCLK_INVERTED   	32'h0040	// Type=BINARY; Min=1'b0, Max=1'b1
`define SYSMONE1__IS_CONVSTCLK_INVERTED_SZ	1

`define SYSMONE1__IS_DCLK_INVERTED   	32'h0041	// Type=BINARY; Min=1'b0, Max=1'b1
`define SYSMONE1__IS_DCLK_INVERTED_SZ	1

`endif  // B_SYSMONE1_DEFINES_VH
