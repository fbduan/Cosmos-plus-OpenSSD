// BLH dynamic attribute configuration look-up table addresses
//
// Build Summary:
//    Built By:     mk_defines_vh 3.0001
//    Built On:     Wed Apr 17 17:24:09 2013
//    Bundle:       DSP48E2
//    Architecture: olympus
//    Snapshot Dir: /tmp/H238lm9sMS
// Environment Variables:
//    XILENV="/build/xfndry/HEAD/env"
//    MYXILENV=""
//

`ifdef B_DSP_PREADD_DEFINES_VH
`else
`define B_DSP_PREADD_DEFINES_VH

// Look-up table parameters
//

`define DSP_PREADD_ADDR_N  0
`define DSP_PREADD_ADDR_SZ 32
`define DSP_PREADD_DATA_SZ 

// Attribute addresses
//

// ( No software attribute in this block )

`endif  // B_DSP_PREADD_DEFINES_VH
