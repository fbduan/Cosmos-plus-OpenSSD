
    u_psnf.single_read(4, 32'h43C0_0000, tmp_rdata[31:0]);
    u_psnf.single_read(4, 32'h43C0_0004, tmp_rdata[31:0]);
    u_psnf.single_read(4, 32'h43C0_0008, tmp_rdata[31:0]);
    u_psnf.single_read(4, 32'h43C0_000C, tmp_rdata[31:0]);

    u_psnf.single_read(4, 32'h43C1_0010, tmp_rdata[31:0]);
    u_psnf.single_read(4, 32'h43C1_0014, tmp_rdata[31:0]);
    u_psnf.single_read(4, 32'h43C1_0018, tmp_rdata[31:0]);
    u_psnf.single_read(4, 32'h43C1_001C, tmp_rdata[31:0]);

