`include "B_DSP_PREADD_DATA_defines.vh"

reg [`DSP_PREADD_DATA_DATA_SZ-1:0] ATTR [0:`DSP_PREADD_DATA_ADDR_N-1];
reg ADREG_REG = ADREG;
reg [8*2:1] AMULTSEL_REG = AMULTSEL;
reg [8*2:1] BMULTSEL_REG = BMULTSEL;
reg DREG_REG = DREG;
reg INMODEREG_REG = INMODEREG;
reg [0:0] IS_CLK_INVERTED_REG = IS_CLK_INVERTED;
reg [4:0] IS_INMODE_INVERTED_REG = IS_INMODE_INVERTED;
reg [0:0] IS_RSTD_INVERTED_REG = IS_RSTD_INVERTED;
reg [0:0] IS_RSTINMODE_INVERTED_REG = IS_RSTINMODE_INVERTED;
reg [8*1:1] PREADDINSEL_REG = PREADDINSEL;
reg [8*8:1] USE_MULT_REG = USE_MULT;

initial begin
  ATTR[`DSP_PREADD_DATA__ADREG] = ADREG;
  ATTR[`DSP_PREADD_DATA__AMULTSEL] = AMULTSEL;
  ATTR[`DSP_PREADD_DATA__BMULTSEL] = BMULTSEL;
  ATTR[`DSP_PREADD_DATA__DREG] = DREG;
  ATTR[`DSP_PREADD_DATA__INMODEREG] = INMODEREG;
  ATTR[`DSP_PREADD_DATA__IS_CLK_INVERTED] = IS_CLK_INVERTED;
  ATTR[`DSP_PREADD_DATA__IS_INMODE_INVERTED] = IS_INMODE_INVERTED;
  ATTR[`DSP_PREADD_DATA__IS_RSTD_INVERTED] = IS_RSTD_INVERTED;
  ATTR[`DSP_PREADD_DATA__IS_RSTINMODE_INVERTED] = IS_RSTINMODE_INVERTED;
  ATTR[`DSP_PREADD_DATA__PREADDINSEL] = PREADDINSEL;
  ATTR[`DSP_PREADD_DATA__USE_MULT] = USE_MULT;
end

always @(trig_attr) begin
  ADREG_REG = ATTR[`DSP_PREADD_DATA__ADREG];
  AMULTSEL_REG = ATTR[`DSP_PREADD_DATA__AMULTSEL];
  BMULTSEL_REG = ATTR[`DSP_PREADD_DATA__BMULTSEL];
  DREG_REG = ATTR[`DSP_PREADD_DATA__DREG];
  INMODEREG_REG = ATTR[`DSP_PREADD_DATA__INMODEREG];
  IS_CLK_INVERTED_REG = ATTR[`DSP_PREADD_DATA__IS_CLK_INVERTED];
  IS_INMODE_INVERTED_REG = ATTR[`DSP_PREADD_DATA__IS_INMODE_INVERTED];
  IS_RSTD_INVERTED_REG = ATTR[`DSP_PREADD_DATA__IS_RSTD_INVERTED];
  IS_RSTINMODE_INVERTED_REG = ATTR[`DSP_PREADD_DATA__IS_RSTINMODE_INVERTED];
  PREADDINSEL_REG = ATTR[`DSP_PREADD_DATA__PREADDINSEL];
  USE_MULT_REG = ATTR[`DSP_PREADD_DATA__USE_MULT];
end

// procedures to override, read attribute values

task write_attr;
  input  [`DSP_PREADD_DATA_ADDR_SZ-1:0] addr;
  input  [`DSP_PREADD_DATA_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`DSP_PREADD_DATA_DATA_SZ-1:0] read_attr;
  input  [`DSP_PREADD_DATA_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
    trig_attr = ~trig_attr;
  end
endtask
