// BLH dynamic attribute configuration look-up table addresses
//
// Build Summary:
//    Built By:     mk_defines_vh 3.0001
//    Built On:     Wed May 21 17:07:22 2014
//    Bundle:       XIPHY
//    Architecture: olympus
//    Snapshot Dir: /tmp/MgzBFkdK57
// Environment Variables:
//    XILENV="/build/xfndry/HEAD/env"
//    MYXILENV=""
//

`ifdef B_RX_BITSLICE_DEFINES_VH
`else
`define B_RX_BITSLICE_DEFINES_VH

// Look-up table parameters
//

`define RX_BITSLICE_ADDR_N  17
`define RX_BITSLICE_ADDR_SZ 32
`define RX_BITSLICE_DATA_SZ 112

// Attribute addresses
//

`define RX_BITSLICE__CASCADE   	32'h0000	// Type=BOOLSTRING; Values=FALSE,TRUE
`define RX_BITSLICE__CASCADE_SZ	40

`define RX_BITSLICE__DATA_TYPE   	32'h0001	// Type=STRING; Values=NONE,CLOCK,DATA,DATA_AND_CLOCK
`define RX_BITSLICE__DATA_TYPE_SZ	112

`define RX_BITSLICE__DATA_WIDTH   	32'h0002	// Type=DECIMAL; Values=8,4
`define RX_BITSLICE__DATA_WIDTH_SZ	32

`define RX_BITSLICE__DELAY_FORMAT   	32'h0003	// Type=STRING; Values=TIME,COUNT
`define RX_BITSLICE__DELAY_FORMAT_SZ	40

`define RX_BITSLICE__DELAY_TYPE   	32'h0004	// Type=STRING; Values=FIXED,VAR_LOAD,VARIABLE
`define RX_BITSLICE__DELAY_TYPE_SZ	64

`define RX_BITSLICE__DELAY_VALUE   	32'h0005	// Type=DECIMAL; Min=0, Max=1250
`define RX_BITSLICE__DELAY_VALUE_SZ	32

`define RX_BITSLICE__DELAY_VALUE_EXT   	32'h0006	// Type=DECIMAL; Min=0, Max=1250
`define RX_BITSLICE__DELAY_VALUE_EXT_SZ	32

`define RX_BITSLICE__FIFO_SYNC_MODE   	32'h0007	// Type=BOOLSTRING; Values=FALSE,TRUE
`define RX_BITSLICE__FIFO_SYNC_MODE_SZ	40

`define RX_BITSLICE__IS_CLK_EXT_INVERTED   	32'h0008	// Type=BINARY; Min=1'b0, Max=1'b1
`define RX_BITSLICE__IS_CLK_EXT_INVERTED_SZ	1

`define RX_BITSLICE__IS_CLK_INVERTED   	32'h0009	// Type=BINARY; Min=1'b0, Max=1'b1
`define RX_BITSLICE__IS_CLK_INVERTED_SZ	1

`define RX_BITSLICE__IS_RST_DLY_EXT_INVERTED   	32'h000a	// Type=BINARY; Min=1'b0, Max=1'b1
`define RX_BITSLICE__IS_RST_DLY_EXT_INVERTED_SZ	1

`define RX_BITSLICE__IS_RST_DLY_INVERTED   	32'h000b	// Type=BINARY; Min=1'b0, Max=1'b1
`define RX_BITSLICE__IS_RST_DLY_INVERTED_SZ	1

`define RX_BITSLICE__IS_RST_INVERTED   	32'h000c	// Type=BINARY; Min=1'b0, Max=1'b1
`define RX_BITSLICE__IS_RST_INVERTED_SZ	1

`define RX_BITSLICE__REFCLK_FREQUENCY   	32'h000d	// Type=FLOAT; Min=200.0, Max=2400.0
`define RX_BITSLICE__REFCLK_FREQUENCY_SZ	64

`define RX_BITSLICE__SIM_VERSION   	32'h000e	// Type=FLOAT; Values=2.0,1.0
`define RX_BITSLICE__SIM_VERSION_SZ	64

`define RX_BITSLICE__UPDATE_MODE   	32'h000f	// Type=STRING; Values=ASYNC,MANUAL,SYNC
`define RX_BITSLICE__UPDATE_MODE_SZ	48

`define RX_BITSLICE__UPDATE_MODE_EXT   	32'h0010	// Type=STRING; Values=ASYNC,MANUAL,SYNC
`define RX_BITSLICE__UPDATE_MODE_EXT_SZ	48

`endif  // B_RX_BITSLICE_DEFINES_VH
