`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
bNIbShH2EA0CHyFd3tcKzqAAHVrbIPwWhMG9NsC+dQUSMA6xt4c379IBpTIXbcWcRu47Z+xjBDyZ
pmPIKJwXiw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
aHvYZyL6jZFeED4yBNrYXGt5D78L6XKvfv3d1wuLye6gycFxQz5GvWsSx0S6xMB9xfjAd58Otvbz
klFCQAqOIJ1v9j3fyjGrdYiRUTQuApDhC+FsIz/c7IXqHLMU7bYHwJKasO9SrDTWvXQ7ih9U0p2k
1AKMnh+qiHrYpQorG5A=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RiEdSHs/Bt5umPP6K79selbyluJtARUHU0yj5nYfHoqZIAm8WpvDCQm54C/KO7nPLeyv8jHIHHlo
ALGpGGe0PjfMvHDpFSP2vV238cyunFX8V0T9k8bl6wjYh6At9VhihdwfU2o+IX5VBj8SP9UjNVm7
vVF4zMGwAkPIQLbID37yUDY79ZMmCkWbDezMLjj3KJUww291O1rtjgyC9U405d49Oz2JWy3P7QMn
8qdrMZbOorlxSjkf+hkEIpgWhS+pbRjZ8wYGv6o7pRDkDsG3+S5QG9lWf289rXA2RQvNu+gKmbHa
+29rBsgGnvv//KXcwxU1LPRwDeg4UvorpCIeXA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
1kXEElfRhCg/jAKI1qgX87/xWqRpS0e1DlrBHXO8aH5H5hRB8yNxfJpWnAEYapsnx3bdBnU1AAyT
aS1HwJVWR+nZKer5YXEg9XX/LwYQGdvNDMOsfvUNry+U7z6Kbe/UEvv6lt1y8KsQyYySOWeC/GkY
gvuKcUlrP9I2nyTJMAM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mYglWFHrB9KUMFOAglZNRnS7Lnvi5gZL2XwL13GIjD89oHQqVk29jGx2KCeeLHh/cuuqyyaX8cnu
wVXmf6095a3qNER/BkizDns2ON7gXlfqDwAiwRQlnbHJVhuv339KnW9GIEeggUZhg16lG/xuic29
kcyTsJU92tL+0bqVkxdCDfWly3o+vB011FmTnOJvdxGOerq/smn5f+CNTSqTx6aWySd4focWp3FP
1IRx8Cjqp34czZQNDbnzZ90IVxyJuFmmDpW8roK21NFNjW7dbg4hrFdS8qcX75ES6c0+1Ad9MDUf
dJImpXUL0bDTxErqK6kqA1RFpvNA/Wd7osKy7g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1000800)
`protect data_block
UZbNrxS4mSBhmAa3/X3oJE8VPopSOVaRAZ1G55q4QhF/Pq3b8DXy7V0jgbB0Qc1XV2La65Tuam7K
kgQ/ynUaNFKOyVfIahKe8lSwARKniUJ5eUyzcI/m4U9xJOzorGEi+mYSQ1oOcolg/y2l4d8U6zPL
3HsbhUXAd9EcWd1mfNpYubRDRs1ZCsspjQdYTCKPacHjXnvzqYwEJgYugbemw169HmkVYD89NBmg
jhqYCDYDTQyNcnLSpK6+yb6T6dajiqCXYIHK0V+VKaAmRiiGkdND3RDq8QQ9J8DbiAjr5kSh8Gml
rErCJxFz8+vXzY2utXY6pyzzZkiFZIai+z3qL2iXlnVlTK1OcvGL9KVl1nR1KeCdyqGcVKVyIzg7
QpkuJlXlIZQo7trF54jL1zgSgtwa+kumx1Hdd7Z7Y2eruLVBEgKmZM5ee13qGVIOvRrGipYn3EsK
LTkO1u+CfMjpn/WssF2VFR//7TkjjLXBZAR7xLj+N1b8dv0t8HibiRwsCyC/vJThztnABbktalPA
ysh72WP3hXCLVjJJumXxAEN/FXnucDt0YHY+0czM7DGZWCckEzuV9mJOcvmuZix1Ioj4kyUV2USu
U5YAEdnpIuS3BkRkvP2f+xtGLaBk/J/nNDVTVl1GkSKVbzRikHeU/A8LR6z2bamhOo3ot2M0bXOT
mJpKfkEvrjJ7HlnBZZuN6tHSzQhsZfetPpMDmZijFbMt0EPY6qYF6JKR/N+R0py8PwaCqOGnwDpm
/2ZCuFZuNY0ZMB8qtJO4Nq5foa1zOOuRk3UnVoI3oB8e64fmWzBNOLtnAkkxnHXuzA12IAKoE4PQ
PoFibVTYRaRx1hn3osW6QUrvB1FJU+igxOq7iJS1rUhnqHZ/IprU7kChoTg2I3uiZZicmKhZgO4J
gRqH6KcUNdcPl8NexIK95q8mY1PXyhDfobuhAvAJR76f4eoRNrHoSxdnISDyBTdSvH4lMUd6EeF+
NMUsnJk9r5ETmgg1QE2KFlGAdjUQd2BOx6OtlAcVcZ3w6et8wocAbwczUe+VzLy3EatDOmnFUPWA
grmd0ev50I3nGUgG/NYp10lYPs4pQ4KJeoK8hwt2RMxnE6YcWXMhObUuljl4NrADy1Wug0RfLGXs
LVRP8nI093pVHFiyxU7atpJf+3K6ULPzZ6T4qT5T9ASEF+E66PLU+kgFDECKOlp02irSSwJ1VT3l
d0UY8HpcQxeNUQV2nbw0note2efYWytJZAHgf+rh+P9+kjSS3i5nW4eyXhHzGLsBTnuRKI+hjKXG
k3CnvBy5u5azjPgyelMf/hagZzVIvDPRY3PW0y2bPKkImyFs5eMAA+DcnZVYalcvR9+N6Sw7PpRs
K5YWYFAVIqM9sWQ1I6N2ZP6T+iRv2aOs/D8XuVTrPzToHE3iiswNpg7m40eqnOhA8K5rjYonqg02
SETB7Mz5AdelBiIcFP37KUzaOBfwiO5JStaqx6kLEs7V6w7ol3I+ERhx4eNzuMl5M9L0J+qOuXBx
O0arFcwEFDe9MaVeEukLZyHCAr+XM0gOAMYAXbfZ/xeuuR4M1nGkzymGSBDl8vKBimU7y1YCWicn
iaxcMQGTkmr95Y9eLWNfAilEWFvVN4i3rhqsX7yf/8MhZMslVuTfcJ5XaSuuXJY7ezbs6CnP0p3/
VdcKiYRNaOlhcfdF3boLas+WggGS7YQi3CXUup9Vb6gWqhvNpef9yjPOXaDwJq4r0Ub7/is2VvTa
o6B9QV10vvTAod69293ec1wqfhZacpqBJPtDgWyaCCsPpx5W2CjJLwqRw6yDW/f1noxfQGD365rB
yebZpzb+0MuvrjVjgackDyiKP3KcerN3bFSTaxaQodIxOZCgkvBcCyCMh3O5/BgeTzXYelRAzZ7T
ZuUHkuM5qYLL0OfKZ7kEZLwd3wn5tvKIOhhViPccc16faO7OyQzcCIyNpD0dFcoW8X6wBgij2D/c
2UNU+Uoi3pr8IuzPSO4KIxfagGOh+/B3V9A+v796giE2TKYANhHsZxXoHp59FsH1fgLBWiGILi03
2tSNmKC1XpezFFhtMBqX3pVSaW8NuaozgndPS/RvOvurU0CSfpU+jJ3htAbE8jUVKSqddzMCD7fJ
fJt0xjHULFwRzWvzjecUbac2EbGdlYn188VRnC4TK7G3Er+TjJ4QGLRHxXWJJuFV/XUrELnrlA8u
urPqHY7q1wccKCf+lLbVWZ3pmli1Aogxw0k+ys4FQQy6lPZf0Z4tLFJLqHefPrFdcqklsKmK/r09
ev7nYyFBpBXqFIDGVGh7a0nRGoOlUJz+z/Xmx8G4zlMPqa5G1B6avh3NFUJpSY5kONhkzhgebXrg
sgA5HPBJTE+LYcFyI0KQy7DmcFolpl3H27OmSXYgNXLBBBhrdJ7/twtjqVGcpi60R21BDn97N5mf
h6ZBaIJSbu2RCENs0wLdFETj5VyftuBfZeJZ9wfBzQVKHxqknimG6hA5RdzIwaVzcTmFdU0o3koY
mxASi9pC1t+yszqFTbAJfOYx7RCt1jwGvj26b6M/spYv9XdtL8chSoVd/XhE0pxAI+8BuQbh9RiD
k0KCes22gcHWG2fizyselwequtS+S1Lc65FtuHW0q4gO0MYhj0AHojz/oHLg3wtBb54lm2bKx3J3
djUoJItm33e2A+u/Qt6B4wHPPnqbyLjB3sh4sKHCIjaaRK7JjciHuooPwBGDrKkxjKaxsYlF3rRu
0kUe5USVkKaYSGg00qkAknpb0TO9iHKCmenKJz33fUDvQcdmZIqQE+vjXNCEtzd2L2a1fKfis2NX
9eqMCYP1SlBF751VD0UEemQIcGj5kuOZE5bbUtTPaoDgmxXOmoJuqaiKJQINHpyWGQ6oJpkMy/GB
4Psfo4ISIFncvegsSceVSqJ9qGLrwAYZzd0O5XA1vrbImz7lZW0JGvO0MXBPmyBnyafFuZmkXFFG
PnDRavsdCI3kjX6b0RUzggNvKAV3tUZlJaKgis6dEQU2smpa5stc5VJPPyaHlsUDWZnUOUJBm3qo
TSDTNcLTYetDfVzImdUaYPYajXx/BMqVQluZJEPwbjG86Pc/amMFX93Xiz8vSXW1JoC3X8xsv1JH
RDrrJDEDNgpn8zgfBUWPmIGe9a/r/daO/O8yQxl8w87r7ZeNSh3UTYj8cFeswm17Wy0kSzlTVOjp
BDSouHL8YAyf0+dD0UpO/0Qm4HG5DyVT1kzjXqonr5CsiX2PwtLbyFLJ4yz6faPzzgneaa5SVYHo
k1uoSgcAKGf+A39cYlWTt1BUXZzb11yVN2rBgYkrkUgiYSCrBVckHrh5Y96wSBxtfCBDmr5ySFrH
cVvLnkZiu25CQEpkuje5R4Hugn0mSSh2CJjBlOxcU1xg1wb5xoSJb5lO1f1aYpOTSmKo6jVnm6ij
hr/ADSTFPzCskYkurYvrPxyEaq6ftaIxcuozzsw/igRrUkEVxF3pOSprZlH0w1ovoa09G1lOG3Wu
hIevZOCANKi4O3vXHTCeds+SMPBLNPU27V3TMJZK3Heh3XeIJAGpwV/SX97oOnQH97y1sGgzI0WX
nbfq4aiugSgeo+bEhQxaS//gn/6dN5HY2Ukpnv6BjeycDBla2ILOepv7AO5ld40dOpJGMaNFCDKM
/tN/ixR34XxlzgE8X3Vuecnv9fVLMfdTLUYlETQNRAaOWU0Z4pnkAIUXz4/oagBdwAMJ95dr8NdN
q2DFO8072ktxbs/S7lmg242KZswcp8PJOdSap+2EUHOSfxoL++eXxH6Vwe/fYXjRnpuT4GXK3GtN
X0O4YBan3Yci1/1Oi+07jtl1bipxf9X1vZjgBt50kIMw7YiReOmpzV9qn7PZzHvkxr4xkWwlfVI6
HrGfbLwArMOmhMZwSiIIlN+gGNM9beHZ22/6eTBvFSCbI0I2K77H7QoD4tGkAlNj98bA7mK5jyvR
Os4gCGONsGFeKMdZ5zdYuf4Qgo/j5JcywHJzPl7GlhXitX1UwMKbR3Vnl+Vnwi2EL3h/Qly89xej
kvc0bKjq745xxi0W8mmKodAGKTmcsTuIaO6g9c0MjCHvRfI9/QzqYMIXClglcJxMApfEgSWxIfgF
TTtSh/Gzq4pH8oOu8OsU1lXU4etprIg9DH5ij1RCM9rNoiK20cuOE73rdcL/utWqBWqOAiZQN4oZ
Xqa+iiJ4biJfF0um1zu0Oz0WhTCyJSeA/cuBxq4faouZ3l9++UBAGo2ULrED5MzBtZUiCAMhWBJd
Fv7g46+rZ/Wo6w8ZDrbGOwyIEDojrb2tJp8OeeMYD6ykvg7mLOxstduknPTkKKT8VM/DstbQ6npc
tqpBy0lY0wuzDZHVbu3vPF/aDlBnf3k4EuQ3Mis/FgfeOpcOT6yk1m5uyyzR7aBTdafrEDXFjoar
RgrYOBhI2edsBWHwEkD3R8OGxtMHCvAILwDLmugKvQyL4e8anJ4lp/vovfA7CmeEHv4sJs4NG9WC
7KDd9y3Hkpvf7Lpq1cWyjGUlZ0SzgKxUBzRyjX3kYsUCTnSvQpWkYqlYD/CeAcsE/qcpKghdjfwA
XuyWOvYKEjxncf3nLHGf36huyllzkJxUi1+4ZvsRHd1w4X3wtkidIdQHmSOCiqKMhG5X9Q+UJRIj
NkUiTHLYN4+mxKAGdZwCNNQ8HL6n+DpVQ5sxPKjGvyC8tNYOP9XOZYoo74eTJS9l7QxwYAxuD1ag
I/8rikwb8frm3iW9bch/RIDHF5ruJEWceer3f3CzTb/oxXLXFQen9F4V5GT97aF68RZ4S1BH24+a
7NXwa1YiCBYkIlizVRyba5K5FIFWo08HXy78yllSu6yLMYFZGYTZQbv1TBa4YpKcQgfewKgYK3l3
3bO9HDseMe8TILSN6zuJjkmM13617yU3pGvhL0u/Tp1ySiwSRwjXhI0GeQBHMoyqV3orR1a/nU79
rEbJc6o1TZh/cqb8iUHQNaksON8iRLmayV3G387A8dOs4w7LhrgtaQ1ahwhVAhsvlVNE1RLBe5Q8
8dH0SFjXqBjusEMuNfmRptGo+GPt4ymcDoJ3U0C6D4ueQfZiLn9WgVFq32KhIpRe1YEcRKQqFRUj
ItdeJ537vad8qz2z0AQGf7Ov0be2Zfzua2g568GKKNjyB8GY2gCW1WM8Q5aEk37B+uudUSnvzzTe
TRraxxHQSnHP7XokXRR/8L/0nxjMFzpDrUqCb2QXML0j3diOZAeckqM0znJDZ/saPW+hiUc5QaIi
ghoHmdXsTqm91uYKyNnf3ykwi+PQhD1Id5AvJKBl0D0/YwmnxuL//9DtOnh44QACv625AWX674I7
ysGUa87N92hUVeObS3JWchZncHh/CNDhJBVesWnZmIT/KqQ9+cDpLkjFC0JseWmVVL3JVitrXpPB
4YOTQfpwaAZZnrcfPll3RytjVuU7Iz98/Y7bwZvHL6iNFPfFFmZvLwEAT7Ezq73VqS5cVFwlHXTF
JBrNXQsMLL8z1NSsaycq1tY1jvguo1RYIMnE0LqPU9E9SgBdc9TmsqLF20HZYw8Tfrz00NE1lCBT
whu7Y8AoFsHgtHLEERW0hp9sk47Jb52xiaB68V8MW3SLUV9R4+A33JPYqUTJzylT7EoExymOkuS5
Iq9tahBs6DIndBegsZDNE90vEwm+hjj+2hblv477ZZgw8q+XenfK1p94zXmYGQlSKShsMPt6xAFW
1T67vL4mbOiE7aMCZeSncFVduvHrvSM4phpqKVDVJZIOvYcZJNIuEVYw4Fx9pSGM6zmJGolsqExI
QS1REkobvlBAIdI9wUVNzu8wPL7jBTbuCfxJqKSrkVajnW4587i9JBGPKVL4YgzZATm0yXNm62Js
njnxKtjs3B7TTeFcTeqTDbdXYwW7kkVqymAGGPyqkZNf9qeB7KkDezMdqaKT0b2d+f6p0WBCk9sU
Rshhe7AZROUYSHx6ENs+uZK9uyc/W09GZx3zkbQ5QK4MLg1xINWAss6juT6VaYD2UtwpRWpu34he
ON11xWO/hvSyPVtz0DeBfiBSFt2GgVnrKvj+kZNpRc/jgv9xT5TwzbXUDZDE2gZK0Z7UokX+wv/L
ZhBxTskO2qSW0CoEnPY0aP+cH7gOGGX1f5lRi+DPNDI55wYMQV7tBSIN9Cynqtv4+piipJN/3noP
Py2tPdUah+kSg34nTXvqD6auVQJgCNF9SEZP8t/+faSrYdcOsRyg7gDSslZReI1CZeGAhwts6kMW
y8XVq9crYAOYmCXsUkRFSEGclpC9Rp4F4TkJ7u2U4rutpW/S3ZCPoMkrQbPrSLGu5GTFqfrptoxG
0Rf7BKoCXfSG6KZapR8BAEwuFOUJVTEDiPgpLrVr2+sewdabgdr63kqZosOefXqYk4QTtnpWC6DP
46N5ppPWD77G8D3OsBfrYdd0mcytsNq1+AZ8V6FWuEgopjJ0yo29Ksp3m6y1Jtl9Kn15LSmC7FZ/
y8fb5wjNia9GaNPwFDyPL2YMW8CQUAtfRmU09Uqf+KU+Wi/9L+LoobCfZ8BGu80KnDFkYbAWVzyZ
v+QjEUsKAloSgonoQiGngRr2pMDobCHkHiUXzeqoiKTn7bVLLPbNsTZB35taV5nVWfQ76fxn7gi8
Tkt+usOQEVs4G4r5WOS/aqlogi6axPNwjujvoV0WeBnuE8Dgy4PwKz0AJjM2ZUjVLxDH5iwOka60
pQFdLvyDtgLJD4G8RuEtbtJZGkLtibgfxnZaa/E1ZocqyQ02wmtU3adqYOMEg469J5ehTZqxEbZP
cdSmZZTUE66jnWzFfpy8WCU08Hk+wINsS3llDufhpfCFkv2E6Y0fbqCb21jPQ2cu0DOWEp0qUlaG
larKuwE1MH7DvP4QwLZ8HarNPsk5p1VvGLCPQsbyvRDTlP0XNQW0gIxV/YP8FNlTnXJUH8vStJFz
G0ib9to/zXEEF8ouBBr+zBrx2BkPea96gSKPVo90e7d9HXaLS0dD0NaVfUaKlm2ZNmBdY+b01tzQ
ADImhStdVLZdE3zNZlrmFQOt3O+j9/euOPo4p/ZUSkUX9q2MRgtauhTOs9qmOi0IQhekyRgAkmQq
GGxVXKuHxtg48+zIravd1sHN+HAaxg5FznpEAmqrAsQBRqCtGMEOBW1/eI5QrGPgQYlZHalyv8bq
K38eTBEbuYGttUhKwlWXv4hPA2Jz/ZW/kCRXLaCaB+HmZSNX30MrlCSo17IMh/kwrDo0nzayHaJe
RuAAKITb7nVwLayqd6zyh7YIk5mMMF4I26Y1PhVG1UtpLXYlrWQ/OgFX4SJNerD2v1ijm18cD7As
4/dLX3Ng8NKustou+6MwsLwrvajJ0oV8sIEcWuMsljI/sUWodXjxDzEA6/iyK6Liojh/zo9uVedj
UgcVcc9w83TcvtWuiTG11ohJ4biVuy4LANirSblcjSy4c9uav47NuRMMYzx5s5VWlm/CkQJc8JOP
GgdM/xw4FUevfaXfYO7d9y18ro+mjBSalptdELfRjRwOiTf/p6D1KqzMjCBJd/V2BlcqKI1ndz7/
AQfUjLLTmTk3/LyYs3Mq+X2RMJ2EpFgi16Q6DgCrmlRc8W1loAvDnnUjNW5Vr80LrlgpR/fGfPI1
30dGDgbZpw7qKXXrTFwTmTvTxunPDJCEGbI7AiUS9NKvv5gyjHAzXVYPUqiWyT1NH8e77UOz4NMs
W9FhGCtr0QjGbmjKfU7Dvw1Ch9PGov7g8BYGws+nQAF5uDmw2BwZ0L93VbV8VhkzgPQKGr3rsBgm
75Xiv1OctxH+YctaTnRD9xH48+eiXTZw7pIJqis6PQdEVez9AmQKdLefdiw6e/BZlAJmaYICiJAm
vddVBx4vsMjUkRtCkrhVUOxNCcwma8RPTZ9XSnmp9g2uWM5dpSknq3Z060cdMIUK5tYWAIndbAuq
4mNr3R+d5yPNx4+jmUXYExqvNlUbq1EENsLZmat79jcyKPeFN+R1QZebQZBLGsTQpa3Yt7xHRMIb
2HHu6TPKER1ZqkDaAAxsN8TXsYtYT+whDEYWhb526T4CyOH9MD2vdPnHRFDsIn8qqBPkS5NpY+EL
qODkRJeS6G98WV9qvccfKly93Pbk4X06On7hagPP0C7uYATX+LORc/9PN1VmIr1L+wq3jRmYdB7Q
vT45v+ZNwU8yXR/P6LgCZ1UuMgfsKNLlz9PhSeKv7awLt00ZL7/kmtqQ/ZzJ5Fuu/WRQSYqT0gmT
zQsEd/dDdHyWGW1c7+bXsEoubMQQLXSa1AZwZvSfObfoplzvdAFBjkBfrsRlCa8O/I+N6khgCUNg
eqHGonIox4xjoJxDJiGNJDNVuWpFakbi7JQeXBQRKS0UH6d74/CtFQlWY53Hbl+6zVFSanfpFFnO
aorvgVVEd0997xgKaV/68platA4p6T7WTalSQYGb0qM6Fg5DfCQaGlvJ2NwbvfeQFd4FB9TNBzSB
vsTy5ZE3tNgXShWZqQj76omlDP0dnQxT/mJFw999n8ygf9LwF6CiIPSPr9EzSbI7+Pq54E5GmfEd
jWR0M+Jvj2PTzeUFN5/hBn5PFjdUF/WEjG2O052vC/bqlHa5FHYaDgaIFpngJ9rSnmU2axLYkyUp
6G1Ur3VuxmA7jrtR+scR01pIa3IVkGFu9qVllmygGWTx2FzfjlwVCojYWH5+YGLq/tcg8zw+DLGs
y6NALquI7RuJL2Wmd4TD26wawSnLdeb0B5WwC5Qy1zezp31hjA9Pje09EZvS5ktbymuVqFHELS0/
DqnZOayzQFqNz2pbIMPtOUMq6NOx8piBjlXBpVCreQfymk7ycfBEL2BWkkLDSUxBUB7nkDtV3hjS
ZJjaYyhu2kfOOxTUlAoM899y4R7oQJ4JPvJ7FokAZB4C9BzxHabNznPVlsnG7ga6lqFW+SjkN6/O
Gg9BVr4yk7QWWiFKnNiipH6Xeo95CyDvsyCbC6JYiREWCbrs6+DjOjSUZa8yWHZcIbggeYkAuc3f
q6qf9b8G0coow1EnabMmPIWZjkwhm+t/l3IVF3NbqPucYlMgbBKoh0+3CwvbzINksb1jdaIx1ctA
gIIxStEZDee80lvkUYux4ppby8x7Z/GrtPte2jKtRH68yq9wWk+yKM4NxPqfnwPIaiQNA8IwITSF
LJZhVkdbA6altL/t1DcGZtZUOMSgo9CDmjYQhXPV/qHMlch5jSun50YwzKR60Vd7DHUZBGr5cBJm
GJHIVA4b3GBlOgxI3HdileWscRUtf98oufJsihQXVXeb3CCOYOLKydysMgkAd1ydtyMeKjEYnbZ8
UZdrDfODGTKJYnZitiDlMsxxnWy7cyiC93PF6aDYcrPPeZnwfpOf9kIcCVQNWpUWszKXgfOc9OKW
MLe02ahuvtIQ4HbFm4Hb1zU3i97VIYfH/Ch/przsttjp9r/Hh4no8ZbmWL+GCZhIS/AHSQK84g9g
6baHJa8QBlWmqDO9B4DaoUxJ2qqnsiKpFjNPLLCUYZBdP4X+NM7aoNJ6/MdgBkr/nOu6zmqxQKtN
bAKa1+WmVuVDc7UHhVQBB1Cc2aRlMa0VkohX5AtE2m9xBiPGcuofsXjm4hBlp1tZ8PWMVMrjNv6I
u8WhPLsM7GLzVL0cBMAHgCTTzUIfALeADoeoofOAXZteeK1dgF8hvsH4PykItzpJRMzw//wY3Q7O
JtOT6sOCTk/6Y+kuM4lbWEfsWcXO7pBnsnmCSpDdo78ZpFoGrMXss95clHjpPEuO3qUereH2i9YJ
Z/YrFq9m7CmbsOPmFUdJJFp36scGqjvddhs57FdAMKyeM9GR0+7a1EUd0XyIIrQlIqPM05vkTy3U
Fv2xkdFNEt9pjD2jld2KsDPM1r7dKHH7Ida7brFcKKV8t/LTYXgmBBT5HbXNkCdcbpl7cxc/cdlE
gH2WoRd1VeMq6lNXg5IuUBFOj98XM4/zORMrnFQQ/zNRvrRpJoLVmpCNUZPZNlE6jpXCczZ1K2pl
7LjMxGdiFkSTbLs/f2KuBpganwK0seR0cH89y5WcsWdSvahRVr5a5nifkkDxmGT9s2z4zE6oA4c8
kQTU61L2fmnQQMWdJAx5Ov5yBiyT+Qr7PlFltxTlIkITRoj7mn2wwwD0ewLlIhx9YUAnfZV7VB25
IdjpDvREjzuWaWWuC8fXejAw+jlKLQBNj/M4ZIBqXgmImNS+O5v7/N9NTJhtweWMQpPzhLxMPYbP
5BcxCHSHXGM8lsubGcyQWWUJDJ1omz5fPTXPAHB5ljom4BoQHk6ZbLwnNikHEJD3hmkUuPiqDUr6
9iqoyY/yaI5n/lySG4+gxkHUYHoSumQAJNroTPgjYzLou1kK9k/LYZATAVLR9+wRNxwIEJxHRuiI
+tBG4SIrWztCWgCuXMmEILAOfp369bCwciyRkipFEOHUumVr088AnUmCh8EYx+8kSApHYjvEgoUH
d401E5XeXzSjgSItAG0RNHOXtfmwLC4iioZbNvI0KJyAoFmbTQtQ7f31UH0R8ne2qcpdSO1+v+Xh
zeNz1oZy1wPCu2vnMhzOrxgpth9cNJc4aJqTAZEIADH972jbk1tyDD2PG7Tu+K/YWZzhIUgctQ15
cFMAYKK6ody7H88IcK1ZNSpPqSODvGQfVtLvSHdqSPnaI1jQXhzlSEPK9etL+okT6XZg9otZicUL
G/bCjHXcosohvGCi6eAdrG3GoS1jgu7xF+0oxmrgKAXRpM+ikesghNGvDCRTIBz/SmDkYWlSCiIc
dQvfQr5JJNLKVmoiW6PruJDFL2Va+LcxbtqSYzJZWS3zcIhQKk9DFkIJGe9POM/C1FRyNSccYSQt
qokWrl/vrKlSCZGWXTv7UES0ASWYIW9PHGxMP9mg8BFIY+r+09n5RPdxucLUWjtOqF9sTWa5tbJj
tl89XRBavt4XwCMgMmmLDK7vOXrkLRxwJQB/3l3gxEaOjTEC49GETtoOZjw8QwgVOdpxSX4rnQ54
C8QKbmAdmiZmPSsaXZg6f9n+zMWfnkfRAMEKdRXy385Wrp8zS4pCBM+GNisQukb9O67bnE3bLbDc
4M7a0AMswlZnbG2vBrEyzW73wA0dX/6Pq6CgMeZLRJn78EcoLweLi/saVCCicG+XQu75HewTKD80
gI3kSLtVzwbP51VP4SOIOiFgHFSUP+l/qgloDuaFKuqWt3UGgoFVZHgbZwYXVIDcNENweXqRTbzA
vQZdIsU2mEE+GMPqPwDWOck+1rkiMphPIjcEbEYrCGIoo4IVJu2AanvLqyZN1i8TBVFoN4TPOPrf
8F6plMwq7XhGCAnzJuooTq1B1wCY214YbViFEkCRW4se/tG30MFqDXXepAWJUPj6h9772q5eUfoM
jd0Y0q/sTPPtKPu25GnRK283mEq/HBtCBiKjtmCBy/tOXGtAwivIpDUWYdsOs7260SDKdcoJWMQa
VyllgcOQNn6VXRKenhCrfHR/Np451mUEqf3Xl4pUOz+jHIhPzCDEOm3Ucz+VX9veAED8b1xbXhfJ
G9kgxgWEZf6/QeUBO/0Dfe4T2UEgPs7UiVbQbMqNh0E2NbBkuQVCWAO2lnItb7waSk5TnB2rkuwq
Ud4Tt0rtSbXLCc2lJf6+U3Oqi/C6TZEsj5Svh1+gAJKrCDr94FtvDetr5u4KAUfo6EE+0IhacivS
69XHOJjSMWFTDgK+SPGjk0qxN/k1MytFmb1FXXQ0Q1pVuUOm9ue79kRWyqGopydABm/BfiNNaa5K
Qs5cWq39EasknytJDqmbSNoRfnZTyHTGbbvGaabLiR77cH/DhxwWLpBMxlWOX13fVRz+05lH8lfq
fMMKBtTzWxFQRsPdZBR/AqL/6vvA11mkw3zvanrrLANNcWb7pCQevyHwgxacRj99CYqUsNRlArqm
1XWcBkFm2HPeorLs/SomGZBnFTtABJIkGxoOja+GTwRL283Av6V26AFCBIK6609M987zrsE39oen
tyTd4trYH7AC6SYqOBn8qdZlmZcnP1/jVmgD4DtjerxvhdhCxHQyljH6gcfsgw/DYkRkK1VPR1Kg
P7eYVpRD6LpCuTkIQ35wtKbKPEdNDRfl/OFcSRPPGcEwh6uujvALmgPkuHzpwdrBH4DSrwoEjaBw
1+yhJQNJo5L0GRANVmtxsgdjjRS0pC0EoFfyUeWq7kJJdumiSvbVVrdsEabCFSRVEQ6hZTNwxGcn
mTKFpAU/QmLfSIqktN5FHTpXORFegTdW084uwJIgD6SEOg6Optno9UZ+Lxp9iBbnVsII/CgVMbsB
5xvG45ZCqaihQmjXuWtj6W8YArTSSNnLAXrgy8HuVPfe12L790iGG7lNGrwaYhE3h0kDnrEXJW3t
MmKH+ZIIBctsykn0jnBSBpypV0SlfBcGFqETH8zZeUiWuhfWHrX4JaIo7Xyf4/C3dLYE2/GeRyZS
LF3DDxYEycng6teJp1OSLa+RSzyJil8KZ3l28BBvh5WlW7O+agytUvO8WMl/xBHDtwYSMSDMhv4W
pBpU3oT1F7U07PCVJOYbnhxgebgwp+BkAnjACb2/j70Q4ffjU8gIGHZ8zVd7URu0dPclEh0ffC0g
fWOhX1NN4Ljqqf4bi8/jIQYaEEEjjJU7l8vKaP/02wI9ADw3SMBG7MBz9fouvuH81WRKB4n4Pc/8
7zbdt1Ap/YclkM0KkkBlHmtYhYKU8hXTJt+RnmjpzscnYnWCkrWHY5sFjZB6CL8IHRqYH/W5oyJO
i8N/CJAj4Vb57ibztO3HqlI5a8c1wTWaaeYAiiLGokJvA1CXHtok4xIm5xOM44lI7ISQPLCARlu4
jeDSv1UcPbPW2NPrBAzqjzr/c45mqt/H8cTdRk2M+IVoZfVaV6v84U/BxfvbnJiojtZUnsZ5CwBw
jrhWxZGdmQIKiQbZGCXC61oyZur/1wrBv2k+sfCaXw95XO3LmHdazVQeOENiG694LqidRv8LWaYf
6DUNE7+SFykUHDTkVwODQQuxl7GHB9eJQIV8Oqk3zsg+thM11lO51xZhFdfXGjgCpc4tu/d5v6km
avAeSN2eK53PJfPEcRSpVr1YNWK0+VfPGfJnAEC1/FiLdHGvEpizMG+U0gStbde9qvpI4470JyiF
2S4U+tiGHDcfi7tkAVKmflsJgSbfz1uU7bEDvnMMGIjSRp2Ra2M0wTV/7n4pp7AQVwuq8qJYAKG2
Amig0EKT2yUEhGWCstur7x1VSntwrD5ZAqB3WI8Hyfz235v2Inmkyr++w/cuCVaYK4OehV6zYe6G
hQ7JQl6qmTnGhYHS0bwBQghNMbg113NbYdP55cokxDDheSL2J2XxLvUHd4Cr0LTnoRrtNdwOdECO
dZHEFgTPCMX8C9mXjwC8gx9zeJGRL+ID1ve6X92qjfos4g7mfH9JdIzpk8INmKe3PYy8eSFLt7Cb
L+dGz2/ycU9uxggFcqWK2/WKNmOBrmfMOjnfWv+FW8oyT/2PuuzimBttkIkb2HKb7n3nurBHMw1k
BrRwZ3CBMWUkcfL8n2tXcEzK6cvMDw1a1znTzM315u+jatXUIpAlhuyhBzks8obl5E9pLWP9wfc0
gy5umly1nQEoYrdqts95SRzRWIFuRw4p3XnUhyYJG04hi8Ej5Hl1mWfwbh/QMpcveE3eP4lH1WYp
pG2SdI7bwj1QH1cbQiLuMfe4dxkd1iiQ/mp8TgzQa3zVjoFphSBekq6t0IWQf2GGnMJqH6Vq2LdX
ogy0OlCI1eGVemivT2X1Hf/07ZOkgfmL2oQzChJTK0Y8pVXI8W7nR9gKRUd2BgvxTLcJd0KiPFDA
+lYFOqS5s0XBLQIbWjenXoYxTKPSZ7Tyrhwe4REkGMpmpmWN3qPoYzMhzI54/Z77+Gx3a+fCUAV6
Lsmll1iAF0uWm0M6dEU9jHMEjSgu4Sy2yMp0bPhK6stQAuyJHFZqN3F5NZOsDplXyZuTzPXJ3i8v
wjefk2AtGoDE841+Mjb8MhqqKkY5vlhZMmQTG9vIz0Mb8gRLRLBb1vZYpNNfUE4eN0V8JLN4140K
KCXymfpZx1zjSPDtV/Tpq5lqwtGdJ9Mc3yUCQanmfNrUgqGle1zC3wbmM7KH9ciLt1+EhnXZg/Ba
Lda7xdKj9u4lvkOREE73hsLMucO6UqMA/wMz2QphPK/B02KmnAVPtHWT9s4cfOe9ltu4sAY8xaJE
eLGqG2dtQf+/eTJsQw6cvCsR6/sLgHbCDLFSdj4cL9Q8b9WMSX3OeM8ClhxIFgj5DxU9MbgNxwAa
lc1vb1ZPxZuPUERPewR+eEoOa6wqd65Sd+0TEjmIA8B/Or3D8S7w3PldTxpkP5C9mC5ca4rcbzqf
oYT4qP3Sz2xnBGJLLJ4/PquVawNjYo55Lt63a445bwyCWZYE56eBf6j7trCal0I4gw1Ww2wthlM8
szcLZavo28xsFuQ2gLvwI8GQN2kDElRIwZYN9V13lhNbZbJOqA6wgpHZzjVip8Jbr8f8Rzqil+/p
zsrW8atoQ6BMCIcT+t2X7oM+T71belrlcFSaucmBfH1VXwPif9Re3kghzSs75aUm60UVc+Xb6krp
1++uIp/CycxV9A0SgE7jfbA56DO6dIt6xVVsAxmGyILf9VCSdOIlC/sm2+UqtGTn2IimE4CTrA36
xe5pNKee3JhCO5poFyJT4xMehkVTtdjBRp5xOhK+qdsZBpUUzzdcRcJsgsP4fqeosmuF4QrqrkVS
D0T57rMebqBXr+K9QJVCScIN0Oqx/2k/uvxAo6Yggb25bGuLEBddmcUNZ7fWQhoJ6TnRL/u0F+UO
p44a2Y2Tg2T5UvRuAdA72/WqzALFsO6rpY7gG7N+QYoBSqWCNLzN9+zY/jGOOijpKiKAfvEofmHC
gTaIRNrbbjOlCEhpo7rPg0NIM8L/ZFCrq698sziVDSU2cTs0uTMY4pomLza2XKxqrToLRJcUZkzA
OPxLRwwfcP5snigL8Rk8dzxZUkz44XNgCAbdACQdn1Qp9FaVKPJ7kKLPjl8WeCjhdfNIqsz42poH
Swl+TdwLqWCwzzh/ANZc1+8cxVk9lYpIzc3T4Hr3zBYxBR0TMe9SRHgxIV/pM1PIg9gGrl7tB4zE
MHvmqkwxnhN3O972cSGH4GJYqPBeHWqjacf/YpBcY+hMhiIu0u8cscgPzAviA+FgVctzJA9LkWTO
gHFtV7YeDa5GJOnSApMYlCVaoo7+Tvxe9GvpdYU8FCLCaf12fyA2tPEzVpYo4uNKVHtYn5QuN2jJ
Nd81yIDVmWlghb3+/tEd7Koqm+2mAlxw9g7lOyqa1AP/vpxg94nfJ8aDTiUJQsynnLDrZNj8zg1r
HLXbNNWYYgMxXCsDoNw+hsIzvxrQHP3dnRUGzkTLEPnqZsjxk0QE4DcqXt26NZ+UMViM0jQilgi/
14k2ynL+deWureEpWUD4w7C7WLtn/En4XuMFceM4zUmuxVmhzZMkYHvq2cSmSTXBHQ+OmjSfYbb2
oB4XlR44PsOFyPvyD6/b2d8IWJCOsYO0rSKvKRvhoVpD1NsGxALnRnOhFoozKLSGxC1lHHUmjAdN
37Aan5M16T4rAwBdrKyWDHpJ+m8xQP1fK8vs8vJ6m9Sm32r6d3OgR4efwCUCSN4hNcjOfZNODKum
ZfRMxrWkiDA0Y3OyupmbrI3fdtqiNHcSq4hSCFJWlCzyVJRhCjwYs8hoCoXFw+T5IkHfaXT1pr4Z
LSfRQpsaPF9XiFb8xTa3Vzpt/+QZSWjGi9oPML2WkBuBEdjfULTXis6wHxAR0qe2ZkN5KwNb6Vxa
W5WI2BolFAL6T4CkpmTeuqXs/nhJqNZ08dqR8bBALIfEhjcN+W689+cartS2D+ILOIk2BONmpKFG
Wrig1x3ev7YCRRPiW1Hr0a+O4cRUMFbi0QiNXmWOoEBGoGjjU29FWi0etBRAK29JLh+0ZU0OtbbX
j9qvXK32b5OjXsO1E4/CDtoXHCbUEwagCNXoN9JkU15VVRMTaG1IQPlliUjggeP6BC6bVZmMglzQ
5N9EoIVXpxkXqmWYDXwH7UdmYWsmYE7qkDB6t1Kx7btsppzxNZ4Mna3CJcEhe1UyRD+/tVbMiD7d
JD2Q38yXQV/oRIz1mi//dHU/1zwC5b3i2wFpTlk38jFEx/YgZ5rlHyp0Vxpkk9Y9+vXJp/HBRxO6
0OVfFB3563RJsdjbbV4k69/pRuaV6w1YBjieDTwnOHaJYMMruJsGdvac7bOEfpfi7X/pQYn4m2TY
fetUGx2fBvnoNuzOKCRdbmH0sbXt3p19V0z7KgDcbTZtyDvwzQkSvFHDaZbfGtkmfGjikYLYUnJN
dSu/UmexMwOBrOLtE6Y4SLrLLcMRpNlp4DlgYszVoQ619zWqBvrTkKfj5VWEH9S2UDW3P+lJXn4P
6WzJzFwFDft5H4IQe6EZpDaYoIwotDyDndUKS1S4ltCTBDlh1EBtTg3kgsgkP5NA80+lDHDFhtr1
aCO0V8fm/vDxqlieCL64mwpf+kkJTe+ZfRrbafwX3Tw63WvY2VomKSQGA+Q9EJUhWD9++HbcinTR
k/7YhYrVH2yrnWqFXmjf+vVfI5/qk5fXLgiXFUJvRPhlMTuUbpKOtBlF0pk7UxENdgqhYg2NobtR
Sm2xrrL/qF5K5/QN1Y4YxB5y59/eFOs6V+IaZimCvv2q1HJ4vK5ZM1naOiKirgp/tJQ7ZY0ikJhb
CHubM/KTj880iDZ8ry3WZto9so86vo7lcBMrWs8hgU2//M/MqA7x877a77J8pDBU9jS6HTVEVwb7
IETqoZojR0ojOJlEpUUw+2u0LqvCvq3h8bN5cqhuf2ejyqLOcY3ENuV+G5arWtov2KXOQNptUPZr
QHFET4zqB4ypVzZuTQ5+RLHyL3WK4FkeCyb0GWb3Xkzza/ukhuZwSHoOTpx6Ch849Wci6g9cU6fs
62wktmwYX3xCqDn/04rJCt39iEkgcACYl+hiUp/MDNA8rkSvGZcyLH039BzP8EWFME16iduNl8Wf
9iRPuUSLqP0IocIRZhCjoRKNUwRkJ0ZKbgCWINhYavbMA//2Sx7kGZnP59ZLA7Zq/q0/lwg5b6uH
1DWk74nXD+y1Ib4/PpJZQcacayU5iw4JgXAqvhvrutxLPgNL9oECyYZq764cBqCrSbuwnR71rysZ
8lvsLJm/wirIcHO+LEFYdRoGiiPa6iP0X00S/0HzqnfInL3TCKpsZrc5rBeigJsaN2BizYt7yJb5
u8pWzoXT1M6WXMzmpijLdCfmSBMH8oA5rBnbL/utFXz2QpcxqUZy0wRPOeKBhuVmlt0+lNgV/4+/
7HN6br22ov7Enhu6cSeW1WzBue11AuBlSp/7UWbqmExl0XQxRA4339xFv63DeGUY2NfOHnvZcPGt
nAf6it9eD+MFvnrvOfk0WPxYTzS+8EnGkvbBR3Y+IMopqbI+sSePXcGT4/ieFy8f/g7O41QiRA4/
S0YxgjeMVh8YKGdQrLwpyzd94OMoPZZL2B/0lUDO2lsozRAlrSBNoC2VIU4l7zk0lDgq3zqH8jC/
ZeS20KiskDTNy7em4koCD3fRZ2yW7eMj5W1BoG5MpR+T8n6e/iHWjtudvF5QwQkM/58ITaSYuvDz
zODChWjgwXXjnGVh4nDUS2eiPnhUHDEr4fSaFrsirKye1tC3wcaCnY6ZsJRPckJVqz5YB0W+JX2U
CDvlvw+nFQckWLzlrGhzfDZsverikdfSgNPfQ1r3EbWja4f8Vs9AX5TKVjNOnCS6LPygG/LRnUP6
fV4w+FNqTi5LPIVp83LyCMDaGXQTSkuPY2rOQti1SmVNh3UBTOaeA4o/C0IQSdMpXu1me8eDjGHL
DbFIWfOaWxL5OLBhHmYBx6DQr9MFYgq9sH2byJRiCE3PtkfGE7yBrh6gUyb3wa1O4WsXaM9Fywqr
qJiUiz0u2kz3M7TGiRa9zWM6B6j40cJrrKCrWTTwV9ih5BHW4L0QtXCk8oq/kvwT/0gRmezcujGf
imm2eKGlKS3CvRp/+o1dBDVCIbVTz2Hc+LH/zzAL+bKJ6AC7hDq80Al8S/I4WWmwwbmMX6jX6GVl
hnbaKf14Pgwl6q3WqwwG4fIfwWHPl1PTbcM7lPdP/5Z1ePHEsjAOQNl2d9C+OJxbdUNv7s7CuWrF
zgs1emNhcxGi5fsWsg3HhRMd//fIoqa21lIIO5iDVYE7EUJk+xqJ9laCz5giPkd4nQT2TRisquM+
ejDOmvnFkscSOUOE4QQR9RywWQZGHL6ibJ/EVVAdWBy4AeEqv56c92oEeOf6+m1fmzEit7+Sqj+x
pzcm0C+1o/rRBarMglyU+gZ0RJqCQ+pMv7K6zEz2vzCHxlo2S3eHjGJJi1YGSsFeinlhXVg+lHyh
VrxgLDZGJh6duHCBsbsT017qke9fJbbbi9k+2oPKQ/+oOZ+goYxpyDbxKOT54cc4MO28FvfnZe7/
rsQdsH0g4VEDnR39aL7za12neQeMpx0+/Sz/OYEHnxmdyN5fYIZvvptbdheBA3OZeOpzTgWhiDKN
JJl7MfjVIo+00kzIUAfBWIv5j9/+KHVNxPRYrAPMrjmJ7H9XA5WAIY3M8TRuVc1bYbEsRk0YHNB0
mN3LyFKCPpMOVC3KGSuZw9/G+qxiE4g/30XVRBLESa+egSYlKBIFvOuT2dw/PzJAyvYtizaGZnhg
bj2Covfi1MosxqDkm0aj0ORXr2LNi4x+PKlP0uztAuHUCO86HDt33bFh6cKuq+ikcNtCmD13qo4l
5cOAWPD/WSPrEYUmaQSyO/hHR2CxN6xYSVOmNlINzKqvKXI/+I1RfzlvIgiV8UlCY0n1bj7pBqOA
Lx1vml7jmnOyg4z/j38cWK1Dg49+8fR6UyaUAvdXgZ8xL0/LmvkWFgpcrUVNruNXcdAj5guaxEpa
4xBzGn7I5faS6/eANoGIMeqlaLnqxT0YGBz2psvAVLcrqzwFwixlJiEsEiRARjJ4VqF/dlro9xZb
al2gPQE549U6AM3N66y8j+JqHKlxgZxbotcIpLSA6Cq26H6DFagC8syZE/cXmpsjiaGzh1nz80Oa
porvYi/H2TZmvWNSHE519xDpGuXTMEZ2IdcMhALtqiPQHjAr1J3tKvq+qh/NHsJwyVkOtluGaAmb
C6yVbs+iSzF4WJKuBXa0lId5una0WOaHKYmMl/ISZRT0gsI8/LDKZcvpNrs1+06T6Yus5mZp/xBO
or7HaOw1Uz41HlGz7z5O0quWeYnFTdFij0KtRcI5lR6OJre7IMXU0/GvzQF90FuGUM40XghNx0nv
RKIIDeYN8lGiKjgTqDuizO/uETL1xjU7yc2fLIw2KiCRf5AJmgucBceu2d9wdpYLuPa8mR0/aExR
gLFD7y2vNdzoGflwgUFctnzfCZq5O55rWnNQy9hrehXd2Pba2Z0ksjNOCfDN9ZHDdWZtd9TUaUbG
O8EhI9wjMhlkmNx3J9QauPTMWkYqo+ZRPYNDNuFHUnv62e5bke+7dsPzaY99n91L0gvAl1YQ941n
tqSWABeUrokJTLXBmPzNh2LCrFdBovIq4cgqRWPOw5uUJbWNWXqjvZUoZIVtyDX9mOawopU9TKxl
nriePp465yzI7O0VIi3UUcIj3QhswOcI2zHy+ELxIU7C/2HuHqSk4R77DfycO2iQ7Oz769+M/NRQ
lLYZlZs0lt7U7RogBaeVKH/bfuvMuzyaadXSJPRF97BQ/PU9eLYLMWVo9bhyz+LfjCC/jhDA6R67
L3TxzAoMFr/UK3MXLVC4xrkjpyU1H95W/RzEVOLMdu8+P6Cq2eAmTd5J2qNhkmyqv0uhdTdlYOnH
ASul/rCKd+0YOuis6iCaOF1TJFwvidb6BS2xCxR8s9Gp6lH4Pmjzv7G5EwRbF6AIniD6eZnLsWUY
y4ed4yiaBqIj8Eq/0Yp0wRPpOfkNbakvPzgmxyRvHy1dFrHwYvJh5MPrt3GrTZiQx47YsR+BYunF
Oz7aI7jyvkmx48qE2Aa+w17lDRO4YKGmpzgbY6+ue4o6PPltO20gvdKxZr8eZ7kaNlkQjKUbCqNb
gZWkO9IgpqtgMJCYPpEO3wf+nCyp/cWP3u+RoVPF7519Xtam5D+YBcq6WqSQuL53UyEryxwAZTeG
65Ty9TXpvGIvStSnr76ggngoc1Q15v/K344sMc5e58WxVQMFGgHAfv8V+5KK1exGybyAjtYmNYLV
VvPhEMq2UkxkCRQt3OofjRrGr1RLYPJQpYNp01uuf/irYQ+BiaIfoFuBRgGvdlLhmcw5zg/5cElz
fUbABhdF680XdnXnX791ZnX0gW37hXziHEj1GTAaNpORc11pDCLvc2e9WttwSxDtfZeZAxFCH7J/
qB9UOM8j0LqNUIOCaJV9Ez5XwKOuMo2N1JALz6xk7POh3fZDQ7HaHj7PFczgjNyJjjQkh5gtQGrZ
hiCCpUMP91BlhpMLdfm/69g2377aibdDv/Z79sxmHG7hM2yKJI0WYa5TTit5L8somnGGbZnOpY6B
j078Dwevvl+lnb4yNzutDrXLoQyrm6pQ7xWgctVXWHSklYE1la2D2HNkrm8J5/Y7lIOdVnze7N4W
NaPWyUvRVx30xVzFoptr/GOu34Ax7VxwJQbHlA1DHtfWAoC+8ze2HQMKWTTxuL6hm60eBE/gOyK7
r9bTuHGif/NV4mMZRSQ9IRnowpQjTMSIKpOG+6DbFI9q7SpecZARdnWwr15ju5KKg59FUcekKfDW
j/Kj3jJVQ3bllx5xO2c6pP9cMml0/koN8acE34w9kGDhcz5x29F21UD4Y21sY2u2Wj1bA0P+6Jxl
fOeGK+Zk2AIviYseZosZEZ3jT0Byt8n9MzunkRzSEtRcLZYYzF8DPD77YXf5HSYNxqNUAMhZswWi
6zS2zBimg51IQ6/CfiyJskNhd7kxj6uDHCXyTQQoTgtpkFN/BmyCUB/aygyo5iYFd5LST5AEX1rX
X1J5h7sAKeTwwY+YfZo6vdfuwbolsv8LDUdHSGtmauxZEUz1sNV4h98k2bkrCxOOEXUKzaqj8ytp
OcN9T8LQ355X0FGspDEdpxzkQNOj32Eyb5Cp3V3nrwYcxTRGDwHqqex6HSNo4RXeWN43TEAi6g1z
zLc+RI/EjkcUcbi0gbnJGRA1toXiTfZD/oxlFBZyTWuF2m7kLhHLE4UzZF3bz7iv24Q6Wxg3HRbs
E7qX9FzIo6yYhWgzRazI+UpMJGcAVbz+hR1fQDbMFO5reGo9Y8X2lnxBBWCzPLlJ6vIElV6NrE8B
JE70iMM+FuZSzFUWblWLyzQXhHUWBy6KijKgbb2/bJ0g8Kd+8EJyqTgN90EH8ST1K/hU9JNQmUXq
usvGpOY5aswfCOPUnsGYsFRBuUCBYsIySjseTFWKC9EYc1XeCjQzK7hI/qXcwO7j1Qlkf2xg5pBb
2G8IVQhYUnbok+wNO3bCggGqOc0kIn611DS3K4ccWYYWr2Uf7jomkGmWWXHvM/SJw5xczZpW5iEy
oEG17Ff+qXiPHqwVmZobpPaFZqGYWuC5rPcgA5NXDJd42iw02mHoAAphwzUN5V19zpUhNNA4gQjP
rwgug5ecakQbAfhxUNPL/POmFkh4/bqhpM7HMPBVQIQKkewyl2rZGC6m8Wxn7cupPIv60sZ1MwjR
eRyK8Xa4phWADwU6kzULmLRUcJly2HHxLpEAxhR6j4viK08nFHXsfCLj2djLEH34coMKNDjpNHXB
i3todpxbNo5Thk+40Z4npvTmNPRYWSMxl64MwwL2ePdK5nDm6RaEDQMhUX6y1EWi/dGB/VVZ4l00
IqsEx50/+OAOdEOK7bXKSlNjNcsBxqoNdQQZ+Dgjed1v7+K+n5MJsIdvjQEFsM/mJmNxSSZNAOJK
0quo6Gp734V9cf3HmsGiVkM0oZXo9835QzyrSw15D/07mkskpG5O+rKtnHREn8tQr/Wf5+4nxWdc
sWPbTcERt4iJcKjDxlg6wTBxdOcuL3PntbKT5z3qTZLbhwH1NAhGL5HJ7uhPufpGUdGi0iU/6dFg
k/RQSqKxutLuLyJgJZ8Txh8jSBMWtAhKq5XeB4MpTlxjhvNSx5YnEbLWOuKPby8fwbqMLQBsEIHk
KRwtP7RSA7pGmiQ3d5UoXj8wwAfdguCLxK8+7Mg87scRzwbZys3ew43451AzD68UJ68iK3sIDo7M
6ZC3L/5DPkjbszYZZVEZkQ04KtP+YLbWDUHR4cCYtgQPCDBGz5kIH/GY2Ojs4qP6ny33Q/hILIDn
4I+WJAJ6NFPhYCQyp6nFQXKht10QOQS7Y3q/6EIC7R6ih0WnkgfE8iTzi0nJB2SHk9VEfO1HUgA2
+Ll3O6ABXJo3DU7OvahilIayK7FhpfbOo9YT7cYIATa2bk7bq7LiDK8+ehom7a1LBuBms+4y5K/D
lugOYSnlBa63xC6lXT0bNYcK/C8X/uV4/NRQOtMDgxB5P8UYkdGfN6Z6aUhRcNmmJLYdaIWuTlVK
avi6yaFWg/8GuQYEPsbR0wDZuKodaC4Z9yj1X6NSUexW+9CbsryJvJTEvwbNHFbZswZULe+pAP9e
oNxen1FdW6ZrKAXaczXQv9+Y4ax6Yu0DikJb+/H0oItYHj4nj8wKCmk66Uae+D+xvdkdQ/74Ox+v
kocjn0/viC2nVRUyLVECIsx3S8FCJ1CxhKK9bTp3lYgR9o66AbiQBSDR2jMnNTacXEdFLbSY8lni
OblsoObTL2n2h3XY7a+JldiJjK94thZeULxMHQlr5nLESVBY4K4OT9D0KeJCxscKF12zkXsELVER
lJ6xlOt41AXelBrde5j9VQl3BtOHMXMKwH8FuY5HFZEEMb4cy7L3FuQuLkWDg41Mk9M8TaFxXsBS
+vqP60Zf/PQDokCgt7Q/BURFbF4KNhoynHZv5jHUyqoBHcPoxXu/qbFJruDUVD8QUYtxGEMGJBmk
NcY7Ud+rZ0trFxGYEc5Q9H0eFTl5behz5iePM1k0PLgP7Su8mL2W7txdjN52Yg2PPBdnKJDsVIPk
HQJgWt82MWIjUvCZrEbur1LJgT4xtozFYfw7vmAQL/JDCsrl3rso80UJeyxUs452mTIJs6d07mLf
ZrFacWpu6C3/Fspg7Dq/GlaV9cNl8nmy66ExJbSyTG72dQ+VVoVmDghKI7LS8g+TPNs8144kBNCJ
uV1VtRZ55YNkB6L9xidTlXzW0hh61jgT+VtI2JAJ1tI7Zge+refEgqeV7xtqspN+Pjn0fnSepsHH
2fzpGIrgeEQQEoRRC4EBE9mBVQ6UYvjBX4LkUKoXI6pgxGSa5pIib1DLeC4+ljkaurkB3ukOyxYs
G7cdwMNgiJ+6sF1D2kOEhB4NZPrbAIUpNjisPP8l45iGKXD/QlVA61/ucehfbkGngmR2f468Ovf+
XoJ/QiPI9GfjF5irzk9iap0uGvsHdUO4UJ+OJn7KbDfCcod5XBdfteKphWnb+bGWDQP6mn/OkhfZ
6B/4hC2mc9CQbmiAW0zMd1ZnqqN7JF9dO+qEFPM7mphklvkKlVLdyWGb+ZWLUvFpifMqJYz1RvJs
oVIMJoSP4zjpZEzkZ89Q8y244eEany1czJOm5CLw0wrtj4BFN3jYyo79vtwfsv2UG1XYss0zQz37
oO3s9NWHuySbO3Xdk1OWsYU+S49auilMCa6V0yCytomzbeQHHkMZnQXUZ15PJKa2MvTx7IlLORoG
MZcxpG0TDIpkUqUndDRrr88btAc68O22ELhQl2m/bcwt2ml6qhWcXgqvDSvjC+mO8FSxyBEGWPXs
pcZHNDrL1zhxDrKsNHuY0rn0/qWFUMByN7WYl/Csy43dB0qzBOp8D3A4m9WBpVdklk6ZAFGMKIQs
nwmEBjvQTmONjFXtvcxqVDro3qWV4fm4SyWWgJk1kdykjdVDarZqgJRRmg+c5BoSaFnXg4L+tzBN
ZUBXM1pIrAXSfnCEjSHRL43C4Uf2q+KQCOhfgZTTI11JVwoAq3fI2uHnY4oL9YOFPBA9gYWxkTIB
HdnbdBn7neckSNb1uwY6UpmZhHlq8GXgUpNsBWAFdUSUg5o3uU4zpiRTQ44Qj8D21FXkWXVVIlvC
UzdvbC26p1ae4FnS2MzDD+RtFdvyhVguR1rSEZTqn6rQiRpxfmKjVsgAu0YZ6QxiqOq6hQJDQCyc
o6hoE6a4pct+prW87Tel7ush9A+PMaa36AzqjtuHKgkzhHSltEnoZGVfd4gVYGhLORW2LCu6KSUS
IHdGCFsivO1DiOi86w+vqJQ3hiKhQasXmJ8kixF3bLj7cQd38REOzynJ7yhTxNkNdWexvH8TOQ33
vrQAE1qdfvqsUliELWJo8v9A4LYoFAJChK1OZeqYSPK1NPiMXQSiB8cSwJ/1Of4F9bIYl+4k4Fe2
VtaF2xBG2Z1y9KRnlgTa3A99fQJnpp4QMIAT2Z6LIuwqscql71YxD4Jdbb54mvMKUxt0VLwgZWC/
FQrl7nXZs7dUE0yJ+sQq04Am7DkW3u2c1R4yb4JjSt1oLQT35MqwFAibiqfMMbjFqBZirBspWgYd
PukpZUIAcb8HdQxnsuqzaEtecCRaRKkuggLi8sy0TSJi3QZ6A7ee4RZEEc3NCk9Kz6WERhrF7tQj
e+H+LPD2APeIE/yF7BVeXAmkdGeW6aF8OxCoiUXMbVPB+LAF5xbOwz1EtD68FGkoh9zkA/Eoz1OR
pFdTYretopT9TBFf1QPLlWSrmt6igCxGBkULyoDYScnFNUFcD7wLb/Jrwyc/3iC1IqF/nbZXn1jm
zOD1ralII20tjPAiyBlx4gOJegJa9EkFFE1WSTY8ZSH2slnALf3zZIgdREKVtVCN9zOvt59Ql7Zv
dGBRCiV2u5CCxKTzOL4rkdYjfgahb7H5ajCVByj52LEy1xtJgWsMhSK3NONQYVC7TswluYPl5LJH
iWPj9A6ACNytF3KZxFyRKFyPMD93MbsP74uu4BPE3dVvjw+ZcIDDXJ3ZsG0KBa4x+TkwtAcQi1+I
1XwStblNtcNFQbq38W2KCCW4811VV2Jh0NaS/IAg/8ugz/pBPHMlSRNphVqMTTbxoAD4slWkvcpE
G8E4FHCoinTuVaWGLG+hWdW0jlDQazGfpX9YZwW8K3LmHOJ3bKRtv8vv3FIEvChZ6sjy9AL0RipB
9353amJWr3+Erfn7fKc2ZeQmAn9mUjgjHTwCDASiUmsQtxhfmozQ0tf+Il7I3zE839utrjzOGGe9
SuG0tZmSMJGeLkyHTnUrAdxcsh03/oxgBqNx7zaLeeyNjyN3AGlYmF2CbSawJYxUPJNwf45TMJCL
N3BODXWkqLLdUhPU3U5ePYTUKiblReMdJO1JJZoDysD4CNIIJ+BoBIZHMAOs49nEHXny/nZ4Xxm6
XqmcTJtKQW54SG3HJ+xJzLCsD7Ouoyrr3FRI7/XyOOieCHIFiOQ7k9jwR8Mgmpq2jp9hckHiMNZQ
ziDnb69gw/W4yg5b5Nb4VnBaYc27diS0EEY6kN5WZgTldTiI4aqpXPM0rn3kAFWxVY6FBnnDpWBw
r2/xF2RhGHYsztvSN4jzsb/rIziDOHW4g0qLQP9tYMI+wByblCbN3UAQvcDC1vvqG+xUKfiYddFQ
T+WFUhevrxqNao4v0/+XxQ8PiSeOrUobIXH0SoT5jRHv44jIB/6q1hcSCi5IoacxQF6nBGAAkr2Z
WD1zgNYdtdIaPIFf25ov8e0iPndRwSdfrEqM5N76eXfcKi21Xbs2SbFJwJBz4ykee+TzylVNEJLd
m7sNE5XJ6ZHcId7GhEMuWexKXzNEcCbXacZ8sg4avBO592MA2di2F51mtpHfndhPAUPZBglarYQP
NvhVGqLnFggjhZeMTrFVCDOrRYTSUv3HPw8LXeis0ftdquSfda6G6W4Zx1WkCL79/zHoGdDPaimW
S1LyzmWTYrikc/02P8g9ICURgdoFkC6R/uf+5ExUahPWVWGYLDcW9z7Mcvh3uKXwtLEBsJfYKCtv
eo8SUlxATdyRGc1vaM8LKaWcZeJAcd4xT1kVhZzhVogcwLJpxo/e03GzTEVaTuPXPLUzs4fKmHCx
Yow7gd5mk8ryvoJ2GIdfjbWLXj+LLdIQ5hKyRCp/S9FZMrCKve3DeJUkd5miWIEjJldko61iqFL3
1cfVJ9+rhs6RciCJG96JDkp2W14knZK6LWcWwWyr8SQRiin5c2teVFB9jV6vfYALEjeY0BnB0Wei
kbtGLsOyAZRR0wjeGEGnwBYbVkQ1ZCXoVvzvUGJvL3bF9F5WhRVLOxAJxnTq9URF46GtU2znzAcD
z16Rlie241xjwUXdSRSWJyV3mrLdEVKo9to0feRj6LHKCzv83p78Mf5Zn39UOmGGK0MjDkXH17t5
i6wuH/WHToo/MWStt2M+BSMejffSzBxM7MRydSHt/O64FOAnEG5O00llOsBU22ZvOUBfWC+y/saS
bHfvUE7/4tsqXdFpJT6Wkry/brzk2bc9FnE2ZSKChaiUBiuWv3zqLDAsxoCjQ+z18yqSr8Li7Jog
iqUVdyTWB8KREs8ZnjxCKR0InISJGl15/lFTDqdNOfhCmUfJHn+FsUd+rmr/VLxEO9dLhAQpXM2J
xcvkQpLuY9k1jvQOdCb//tWrON4AdvsDodv1plp3lT5hjnTNAM1aRwx0s1MJMYARvH3+sWOkAbnP
92nO5EWVLErshRiEz0nYh/T6aYOk2ugyc6sS9+tFVxpDRDea0c7kmp6vbjrbOXVmwzqipwT1BpmK
z7jHYQvyg3wPc42dQhWaLvAbqwTBWRu2rVBmNybzo/UjWVG32zRdlijZlmC+Uzmx72c8D2Nr3o61
0zLiwuRFnn8WzJwGz599x5GQvTjwahnb9WsMw+NN9JQ/CwQ3GLHtke6qzEEN7QGXW60mVDqfbDRp
bsWf3Qa4ELLbTo+Qjcr3EQt6Ih+K/Oo73jsRl47O0ATefN8A4UEChshwdYPfNN41wgTvB4HbiY0D
6pcpE5MUUU9ScetQuxcsYNg/XLzmDG1K8Vjpw2+plyX7rpoyJImwmFAU3rmu040bc1+pUuaQtYOw
uNB7zwvvxVSVbJdTd8k9GdANB/ex4s7Jm1OP9dpwTiTGYHMdOR0Aa8Kw8wmALnqchw+/Vr/VJEVD
41yC5BsCAFliWNatn/EBwymfr3gHkINOzHVPLWYe0Wc1WcKyQGmqi/0wwseME6Cper1R/n2d9+nm
pNXFrZuo0Epgf1nvTN75OUfyBzz+MZGZKAS4j75iEgyvfhssfw2Ec/Zjc8cigPkoQBHCeCLzIzHX
IFJ3U3NI6hUj9RunwcHJV+CX4Iyo1cTtuOWNFxuBmoAZU/iQHizhsha9R4iuhDIUNBIR2jT7J6zJ
vSaaNX4UHdjyl9P4aC0uGSG1qsCx380Vgb/wZooJuTfTooMWHk5tH8e1HfrcBXkLnoa3XHstBAf4
t5A7NuAV4VXKW0s4EYIJy3PykHzL9Zr2y3YaXX0qush1j18PUH1pOhPFYUFtGPQLvO1e8ey5jMQs
eJMsXWyeFFIdg6olnrHjFsAqhrEv8X2tU9bfdPgq+WBXO3lZ92uG/jnKi05NpmJUgZiO+q5Tt5Hs
LVN1rJoE46ZARcsYk0eQI94poAWR2XDHn27fhL5w6/afU189tWwGAHDIWYB0ifVvexyadcq/EFMh
t+zXkTmUy8njvFI29iawF9Px4Pa58rbvz+kxamMYPNoTiQQxTyCIoQMo1V2wQ2NS9DbYyjsR9Yc6
iaFyPWjOuBNuCqwFQa5GpSuGmAFxVKjseS8txcjVQbAvYC7M0jVwz7/C/ZsijeUvr5JAj3f0eQTO
oEHzNS4M4TfG+I5OT6tp90c6fjCuOkxiIfev/wb8MkIU2B7lWjsOJ0l0m4osvCJLp9HwZ73vzBrk
eAYhodpSn2nvmFOIkrxMJMdSFDrk4MygcgJbWnND8RImVghy0pDRWg6qZr3dM5WCWS7qTQKCLz8F
xMjqP20L7+QpwHjpuKf5kTpqBDSttCzQXwOqfjmI9FXAOuGOdPSbYWZRX3qS7ruYI6xEiwdpWt8F
d6MDnYKrD4tqM4KqyxxYLq2O1xVa9LMgo987yd7gieIGG6ED66IfJCZ6e5P2PX7e38PaFt5oLwSq
IXrmiQsXzfRn6+mj8WOBc5CA5PRVRU/5IpKDSCHfq8zVN8SEiPSKUBMeDBFmEQ56C2L+NU8LEkXf
NyNHB5h+UyvotFL0xPWG6t+YsQsWd7YBmfcRRn3TcmSJNTJGDeu+gHZ2wLpHDNoe04YRdUtnDhX6
xpbRlrg7O1Bq2PvGCnOyEH/yF5dizcoyW6oYNX9jA3p8e9v+NPEOPwxJww3zWEb1+QVS/KZhR0Ug
IGKcBefVQMVNzV0n8R5rUj9xiGFYUVWDG+Pyywzlq+fwGbJpN7AUyAlExa/ctNbiBClHJhZTMkzH
2DnneM+ajXIrmcLhd0uIU+NVzuPaqFKk9lC7O1MmYvyXH3Lknc6Fpz9YOMEvfuA44R8T3OEMqvhE
8c1cEXMUXfLeE3/X4bp7Ir77HB1mNorodSY8I5ldD2LxdipwR3rhiZe0Q23y3WqZ/171B36pSL4/
iFEr1BLABuOL56V9vWdLt61Zi2HGOCO3YXAtSS2HzPD8eFWHRyDWidQta++jW9/zf4Rj3Hn3tP6j
/fp/Sz9Xdz9nxXOcdGa/jHOLYKo2ForDd6a8+IoZEkaeOVa3vfjW1mNqC2jCfO96D5ArP4rIesax
pZo4Rk7twdBxIrSbrFqNhSvouzA+mRU84QX7fJ2/4aONgG8I3d1KcfViw9hk5Rg7EnuN3wzCMGXU
rXGlwnBczce0cm0japHAQ1XcBQ/0D2zJdNB0kGIJn0TcepM11vKAeYed45moAuowIJu3ZfecAqFI
SlyOMZx58C8REMDItyPavraFQi5Uc/+eYhQP2iUUGVKH97bwzmuI3xL847fDivmzB1HUxMadfkOg
H/jNYsBkHT0kRObMxzlX9NgpcLvTvkc3Bx4jpcDz9+SUpRg/CkATDzQeVuDuGUPmCnGf5dW2imKd
FefonhDKKU7mjDYf1uogpzYxNYJiUWNBJ6mbNT3s1jmLw5KH4F94ud1hdOj1+lLAsCGZPn1WH7EV
kFW4RdnPiWcgB94no7USeGWzkGRm4w9gj3u+bc37rJyKNsTRK+b0YtJbKnjFCTqaFUB3l8IbGAPZ
tSsLv+iReEUElkVP+Q2jXXG2uMTpRF71ps9eJRfCTCsf8+Z3ToBRfCUDm1SU37zHi3yGkSSI+x7v
08iZCJILTb5s5Ed6wbamWSOdXI+J4trX4MCl2Mn142gw/68Cu5dx2QaYXxE5ztyxkkHYsl81AptH
2VgSu10BxsL8EVkd5JDAsW5xFyuXSxcbZ82OYyez9kqhmoYynEdL2f+ScF3DKQ6VuFncl9ur3vzE
hAeBC//mSc5Y4YEDR7tbLSKmwzS6oWwLBJCcNsx9k/OkD27BsMnaHnU2NAIDB5TskEfIbmK5zP4H
EdUJFu5CdI4EiLM/0t66OK7AmuSNyFPyeWQSZZex8EuJjxxfxDFXppkNnkzN+kPomHg38F2Qp2wv
XIFMphbUMVYXqePpPQ7NOQ6nieMNV0XcTjxpCtSwF2Jl3bTBcblOTDaDXc0+AmPTnDHvRyz44VPl
nYFfofKKzeBE/SbKgWS0Q2I7gCLz1Gvq/fd9RG6vHi2Co1U9GX4z8B5PjS/Jy4Zodk2VM8SpqAM3
5rNjiCylAiWzSHxzzDNqKH4kROF2rRgzvQnbznVm9Ep7AroaeujZHtTBlEd5POwlRdmKf9A8vVyz
JINHPQ6kmmSS1bbpGPHtea2IqT97Mi1O9XTV2dJDUQRv8Ps0XBh4dGCjogbrW8gghyFXGxR4m2cE
i95QGeUgZQvt874nhWBdvdNZ44K0E0c1eB/ERoFkgElc9l4RmZf6XRvSSP62UfEIDKCQp2PZ+KUs
eJdcMb9UXeqSQlZpY1sl9WW6+mmaQQeskvGCWbX25UELYPKIS6S0ow9cXNs817z2e7m4b+OG1TAX
xoO+hs+98bh+E4MJujf5Y+Y0vj7sDmBDgfifoazNkCwnSW7nmXDZJNKq+B4lcVmRPXaMd8OAb3Sw
9Dq6PIBLO9rn7Me8MRVnNP4cuybCuUY983QdjS8Lhp36QgO3eZBWpCN1F5ZskhD6tW8LuGq0Zxlj
VMpm3mjrxYudrkKElRZAhXxkGhgm3nQvAPMX0Y6ewhE50+jAvVIpLIkR633Z1xhJPm+i0R2Dbt5B
/xWfDAqOSxpao5r+Lf5HG6RT4Bfq0gk2v+HOuGssVjrxD6AZDUju2BBUnUmtZ3P7NUoj8zScER4+
Z91edOxl12Q8c2GuhyuoU0ZCwKbUUls6vF9yOk/0bP8VeaDYM7sh38EWzWroii+bE3qokgP5mtW+
vrSAcXaLdcwDA7NNoR1JcBJHRX1rm9uW/kiuIEDAWrsZHvuR2Fz5iiUt6bg9bAyOLblyX+HMeXRD
cNLzoYsXUivwZlm08H/YTNz2/+3lIJSFOWkv3ye2OIc5tN0J0ptBqlY67/ah6Anu7KR61rzQxcNO
vnRmkmliMCxeeYIzNvPE5x0WRZL41JleGeiDrzP/jovgKK00eWZBPe139DSze/nIQazQeDO4u8to
it8RdEHVQedOlDARwvk9gW5Fsfp31ZOwD2kNTD9QN3oHzbgupsE7jfJZI51d/9zVgU849tA4cJf5
iYAkOFsNxP2j/UghF0t8cQ8RI4n1rnqobgMSNaJP6uYTlfVa2Byt196WHtgH5bHe8DHHfvGaNaez
uMv2DAI5FyrIhDHcR0o6h57PXgv0m1vifTb7UGr+v6UuAe215J/ugZAtGSRE6tuFTeAKpmO7nn2j
SXZ3mG+khiAs/b9ZZ9N9JqCZVrni9WUu8RAamxyRUioS/3XEG+L7SN7EZhqlQwwMuhLEsVn4kBIs
oIPDKh24qbczdPup20vp5feCyjvvXtQsoDY/RsfAPK49s5ZETr9r0xkdfdvjLMVyBnQUzd3uF7Ek
P5L7mfgpHqlOG/LYtK/WAcjkl1cNLDY0MgqYcxG3H+ZDnXKM5/bCvOjwHvkJOzKg5Zq2eOb1nid1
Bv9wt/Aa1vuVe61akozmTDGJRVykZhw3RfWnJ2i49whTfwomXv9mn/LihGGrvMet0V98AgoHMoCe
7RmnuK9mut9EOjBvul2PTOo+JeiHA7ZToSBD5iMJPRAOrDBmLMncAubIG6DDi+y+pZrcOZxwvNcm
sV+y9WiMdsXF7WvRCUkU+g4V1ofgyOtBdMoDE4OelkvBJW50pA1NaGQrlSeucHF8zEMEN9LNLpRZ
B2PZBntlbAT4SclcdOV/LyzuNDNonR8QkFdKrzZBO4MvkpYHfvGvcI6FGUAC/1OYCZJynAtk98gs
6Vq59CjXu8crHJRvHTJLKyL+zAlEORFGOIHDnXdPB5nVxfRIMOJTQeWxILF7+6gpvwc8nW/BMfik
RTSF7tNLGFds+ZqbzSsQ966thxLuUTLIg1RmJ7DrigQNQFPQPuAzhBIktD3Q1dWtshWiha6as9u2
Om8RJc68y7podP4JZl15JgQancz0LKqgiTiuWFpoH3jwEX1k6+A9FUiwbuL7/eF4momUUwfjoyp6
YzVzVK6hmJjp1kla7zpf4JLUcRZFn2WzIdmbx/ITG8LBlzeoWGCkneCL0JXpBUQH4Jk6YXvgZpUU
54+P0KyP+fguocJjznM9bVC8tiwP7M4k/6RubCxjdYoyeH0CdTxQ7Odo9VtuMQSRVeFESfbBnssY
7aROxZXOVcxg0GronnhZBO/itU4hHitwK+ccikunGi0BQQ2o+gy1b0xm0YMqElDdbbCTMjT2Hw3/
QnZ53qgB8iZTo8Z0ZKkgrrv2u63axjqGcPMHgWF/xvX9HXyrhMWg6TBkJ52+5OZk198WD7opiXlx
RteusJS6yMc232zSiriGGm7YSTOYS8fYKyC/7WZ8+LTzTg9CetS2jZAxKLAsBWKHCdk11SILePNc
rBfz6Y4LaMAEre16DvkBqLps4XN5SVuLJmGJNHr+FdFqbQ/yUjdlSchnxWo6HT8GPQo8q4gdOltE
aTUx38biYXL4SwA+eL5aB5p5SR5Sgs1Nu01ASSDPmXbxtKLqB5jTTzBFOY5MbbtVSUY/tSPYCAKm
QrlU+Gp21Ri/0h6ljlnG5Emi1Jugc7DkAc9cbdUNTDfTTFGFrKklAAgA5nhy6FdhK56e6AAX6kUi
Q7uYnUtdowVHJxYdyzfJ/5SHwv0aLXZbQWoR/CWvoXnfrXigmK8lQQ9IlFrBec8g9fB1KLn4MX65
LWrsaEw6OKmqznmNq72UtWTjWtEMOpRFfpt39C/oYMObQC5l4gXbzAe14Q7YnXti08MU+Hz3/ATB
zjR1QaMc8xuMm4vF+hj8f90zRRInrRrQtFw9ktbc8vHdT+vxSzNoaYP4X7RxsC6q6nNW9jYcSNQX
gQrk6YOJK6fHH8jABkdmt5NAQ+ybLhL1MvYG+NQLP+wP4SiyU7a8vaX4ZkrjSZjTMrNfyr0m9OAn
EWja/IzvPDjtIjHuVv+ES8LVPRysj4bXRK2BZyqUT6407E/ROONdji91cLoXsYSkmLAM+5T6xMya
BsHfmQJClf/A/BopBVm7qLzNONQWeIiTDBmFuhnAX7VdJhbacAXlTAOAH0R1+p2uWWRFHvQjwLYC
oEeMHpnmRCPmoFIZ1CJRrUVSW/IlLC9LhfkoXGydEdhAfGbWaSsGXRo6N4hRPiQbncycg6wAvh+S
UGbZwC6AERKULlfiqr5keI4NaUokk0F5oDZglxIv6Z4W3I53B11HHAgVL/e8gyNjKWBrS839k2Bi
sWGeqdcxCfFDPXUmZFtusuf5axryQr/CVyQJ4UxAGhkVEtYRcGn8Tmhlu6k6YGWyAojeUNfCeLPs
IMT0oDwAz/7zGHQcVcL7e67pPrNnHt95j9XLmgdRYhZ6rcYFJ1ERkoH9Q5UEBbZTKBNFMS9d2HNR
stpUOOC0z1JPARd+j7doOIJvfE/ihODqbzdewN0wuWYTD7PBhLG+Rezt5FWPvxffGQC8X58gd6HZ
ehJp8+TDDDAK6bCaWy36gjL30PyTBFncY97UaKL/Pbx/Bp8sM7xjfegwHA1clMxSAscnVyRuiuOO
Cf8kidrmt8VtJRzTobM9wZ/TBGs+7nwNsKI06bHFQMABqUAxX/bk4sIW69sdKEw7V5hMLOnbP7sL
jj9GGN6NHEyw8AWIO7ms0x+/BsUdLz49ABODVMMa0TFO8U9cIUlTUGf6VpWhMaMMHNwOfst2pQML
+vU7Wy7d77vfvXx4HGf4n6KC8pMi5UH9Ao9Ju900JMSuwbNE0bUaEyunTL5GBCLQacJEcSySWrx0
qSC+NByZOVICBxVTzudZBkw6GpWtpNbRGkcOzJLqk6CvSjItB/hYHy3dBIGIRN9OYmb4zjTYBNyy
UIjT0EhEOuVJJ/9yQjTCpci2EZ8jkjIeePFgfzqThL6fBmakgS0urwJU0EYQBR9npbO7rSmenh/u
7ORLxZLyNDWerjJExogF1fVdtk5WDPOoFSBBOHZx4bw7R1aBpizTfvS+/T7x+1Z+/x0q8lUrovTK
/G1jh3wg3K8b6/ugkGPnI/N+pjHKqQqEl5hua2mpAhVtIKDZROJdQK36NULBU9dx2bYQp4yxZ8aO
mM7m+OR70JriKy5fdQWSnjEyCO2B08AB/jA0bKqBUn+Jt8wIYtlIpkGrPmUAQirSrDtwbPfezEaQ
7NGIIqA/Xd9ZYxU3v+fEXDCUMqHvNYBBya8gDy7kv0Op+nAxvSQkhLfFByXLKxuP8h4/uXXmGjck
wJLcd5Ulys3VWq9P7FiKI74IlAib4a6+N2FNpdFKcNkrTUX9bVGS1MAoyIZ2q7pWiNWkXZkw0GaJ
gMBhFVuxCUConOzplDNxvOEJk46YHA8yqyqaxZx/3mBlwYNK998vPIbONKDHC1pBgS/ecMPKGER8
AoSKkMpMFnq3u8935dAOP1wtI+3zHxYS6hQmJl3M6MrxfByEX9GyAEaTk62YBkKoxXAAV8JQgOYM
Lv14DSjP+2eXx97xBBrYMBcEcwkrXshjNSpceDmOy+gG2J/37yrklgDSfONepMf3xbZ5wnlhdhaB
gFcWv5dnIWbT3BrYlOlQMfop9Ad9ZnChoBzKTGlQsQrCFi/rnOyssAIvJ2s4AJhJ2A5CTu6rMvtz
5tcKIaLxRf9r9UAif45zJvDNIs1oXuI2OAunu/p/cTmliX3fkI9mkDSKWsIDQZB4wkfUyUuL0g83
omgWstVwgMM/CZ+TMUyKCURoF0wfP6mj6bU3r3EmTgZvKwHx5RwGKBNzP6PkGwv122QtxTSvg24Z
4Z2DPB0vNm6NbAnO8GpIeSZ+7JF0iUi1ypjfGvyEBxwDA9LszoQOR+eVfbQWGkAI2ruRmji3gig8
BuyAgX2QfxooHEZjtGj3Qq+G/wSbbNiWyiZMDqbcj0RhCc1j2+KSb/ScEUNHEioW14ZA9Io3qypb
cOpI6JUF4GWxzqAy5BvRDoTny3UuDUPk6E01aFYQidJhglVU7s2yy8PnqaXs+rIc0UEzgWC9qdsp
pJGO+qX6/tZRC18jyvezgj7oCuAItaVUAjTAPlzv1UC3DsTpJuRts2KzvZoNUZFBgkclKJaYmi6a
HuANtAM62ktv3EfO3eqkhhnpRsxc2VppKcmQGOovnNkOaz6og2sq5Gl804OrtZPGlWIIy2cOT9if
mVxaeYZfaeIqdrO/Ad/VMv8pHH4ta8NrSTg5dya52iNLkIMP+Pdaehy6hyc+5QZmBAPQFyGn6IqA
TMiGmSv0NRIOrVMe0velnsngRd1mcCOersR1CeLc8OxiSNPXiCZdZ2vt98GYopOhKIDfoSGsFqcw
iSJHkWWTEfjo/i9F6BoJBSu245YsdOdgqP+odFqd0GyeiCrCRlv1s75g9feKnX9GMfv95yeABw8W
Fv103NHLl+Zvje34eUVrQ9LRfSneQl+m7/djzYwUcDr8BW+Bh93O2O90Rqu6FhlOr4DPk4DtU3Ns
HlNg52MyAivdbR4kXXB+dQGwaLOXPHmdpHCAQFaAYbS5B7mBJJKoYsvZu5Hl1HEH+UDRyiN2nSJ6
+Fr7n2QJ5bxiRs4UiElnAejzW5IG3+O+ZqrjiekiC5YHhPWJh1+tFz58k7D8ejLHSQimAMfIssHL
creuJMEMjF6DUaRCA7YDnf/x+kKAT0gXt6DyfhgjQM+5Yd+jvSXpOpAYjrL6FBjauqP/h2dkmIbN
pb0AbvYHBHvhyc0DvDGk6rAvWa8G9OXAkog0JeA6jGfmWOZyReJ7cxypP87Vvr80/ItK8/X5ZSeO
o26VkiZLxLUWR1M+9TgaUk2egGaB9wYK6M9K6n06zdYvwjjBCtC7PHN32/gG9wyCrYf1qoMpnqmE
nSI+KWJ0TBFNRqcN04B+tTz01UA7mbEahqMaXBUy8qBgva+H/qLNfQo5CQzEufmUSYjT6x5jVdZS
fP6eyUCSi0I+cEx+iR0u1B3ApQk6uPnL3hDO5QhI2OMCHfeCSbvTTdzsXgGJ5Gl5SnMudT76HZ7u
Yz2YV1Mhx39e9Ax79AfBvDapsn7iMKnnT2BWoA1f8qcpgon3wL6Adn3c29tHObG0h4E2TXBDR4ft
z93edIthR2bG51ClUXV3a0vG7KkjiHSmcJ+mLGg5UzGYRi9GKzhIoZVvcyJabq3C/+p7EyK+iry3
NVwJeQgUWDvHtwMp2z6Yta5NtiNPE2ipDcKAm4DWDx93VwOiJ/NJjmxnmyz2Kc9CMGs1vWf2z6xn
FXokOLBVB9dStf2V9sNAkBJTqn8dMcD4ntLDbaSh6iVpnnIenH0rlXNZcRr7B8vXRhMeZqDm5BSg
KcbW9YtYPl6WrmppPO4aLgl3Xjx4xWhMYVgJJdutWhIFjh/mpFMhc1sTqX27tPacXz1aDzb4C3zp
1OkBQgl9sigWeS/3cy1XHYqWianeCd/tkg3ZekheaFXLYJGwjlubGSr+H0FfEl0L+4rxANTuvTHr
6kNKLYsXU0xtH/s5myeC2LMatgQ38gki4b77OnqOXJeFOYy4SeUzfe0RXMOgxJAOCQn1m6pC2+NO
qZu6pdIAEIpr6nZJFDvplY337q/sY4LbpgDYHDk13aqEDKiv6PfDmv22HuqKVMgS/Xc9hwXdyvc4
vMP58nMCx5vb+9O/ahJ3YndYn51HlL1zp+OKH71TyGg2gF7GCl294YEZmgSrFQfTyNK8M9zqMCGi
igbGq/e/p04j7bv8n9LH0XJ3pBbgZO1kJcl+ZOjQUNcrGM2fSXsZw5nBXmHDpJ3EBolS4ifFYn+z
Mln2EpBB9Aic5CgwNUxxQuKxT8vgHs4BZkYJIQh89c18TUpna2AxcSiiqHKjOPhThoUwe7vqj+5E
PlyQLdkq4dzM1WmEUmuUSNV1UePjZiM8udqQb8AaTRddZZgb7AU2U3OIxk7uUhzosQOtk3EqmZUN
0fKfCP1Mq8s/GmEhCecpD+Ry8mxAette+iFPhVAmcBVVHxx3ka7EUldMR7hzoObUrSPlzcj67jXf
qrKzglFb7w3eu9vhswXAcUn/0ri6hilAcTOCFDRUTcHjfO4ebV2IhaqYHBv49HHMwtf42CKiMRcn
lQ2E6Bz9WcGjJebjKRakN+lGKq/dvgtirf+51454Es6eGM+r2Il+HF4aDsbMCoe90MWAvHH6QuyX
BesXMmSYaLoTgGYjcmzc1AiPrf3Lzbe3LSYDRvsrgzt8hvk0NFLLeumD8+NpybH/7mUu20y1qeOq
6WsNDI1P1LMW5bQ5SX0cBcV3HajonNKlTT6uUwxCu2ipzgkKpv8ltkmLVNrgJcaS97MWg5ssWKaX
UwtfolWFG+fx5XIxmGbf0CYEvb+8xtLr51ScoBrAsZ3bC8rWL4KfXMdLp9F6wq2tHOW2RaqBq2RT
8FUY2XTKmaoJFj+EQhRMX4O9yvhtYip5LXpsVGUsx5EObNT0bBnTJOLyCvP0rYOAt94vX61ON37J
5GBahTEOWAiw+F4wyU9lgfJfW7/IxbOgC98uUsafKUbdyRUaAo/XCYHOxGKysTckQk6/IhxTa87H
rkcvIDz9vP7FWzAoR57QwkepUUfa1h7zQ806nc9NW03QFUu/MdmHl8X3v8gI4GA6RB3SXPB30XYG
eG2MiN7OtgsDTgKUu2NaAgL0L6jJ7XhRRwgB2drnDFMEWEv0GFb2vugJOt61GQRWOxdVP5K2bfN1
PAtmUfGzaIxTU+BuX5m6gckeplBtXhN88u8zJN2SClfQFgDye711WUl1bHDtrTLvvTK2eJFedfPf
qg0Z6Nwt09IQkgg6KzpARA/GmaALHxqPn2hwBV+YOOmbl2NpvyF3lm71/nzmHKOUPBPk+LpKd8oZ
2i3i0v0ly8OjA45OE/hiO+/r94GJz4wwuY/R/qTheZ1DIEEqBoYVfbnI49f/3MLYUBHLy0jBXwtU
6PhSHFTMbzCkEdRZUfHb6tRwHGSfa4hcZiIPGfqzjZlUJ7Hdowph4vjM2UBoB0Y61527vaZ9NKs4
5xooGlKh9uNqXvN+NAzG++pfgyR2u+fuAlpYlNuefrU8d0wfe4LiAg5WlfAWpohKRIDEHLRcdXlA
d32iG3mCcwlqQT3eaHTCyw5DbrlhLbTaG2N+LwPoj2OYQrtHf/f2uxd5Jr5ts6s6c7TR1y4egGS1
RPULlQwT7sb+0BctNtSOh0snqJUUlcMInoO+vTFWXksINZJdXpTaPfkBhAYmn93yENtxjTWz70vB
JhzmcZXlVwLeXX3Nq7785sBTArBbvYIlCKeEsLa6VZy8tz2/A0PMnswdsIqyl3WTQyQ5/mJ2mGWI
Tm4PoxzcufjxKdyZ+FQAyUdKI+4QUtLH/8e3HPVwfq2WH93ZLvS+O4E0jEV5Ao13WUhY2OSmf8Aq
dIiCZhGe7PP8pBpzlHX7RTUzz3ygyfG3W133z2tdStxrNcLVVzscpvX7chnsk0hjM7mAovD6R6oR
A7NJia7+aYhBfyxyrar+wGFJvesqKuXVBiUO73QLlWRaLSaHW22CkjZCf7CK504KhR7tgiI98Rv3
uL3szP85pfFKxp5DNoa982wPcdrSzlz8gDOVqK4zQ8Z3L8jaXG4fcoeNZ2AZzzTHiIZkzsSykzmU
DsY7EO9x+gMqvLaxZgaHDWKre8zY8b1ETQe0VL85Brce9heLpWbxWCYoOw80T0nzhkawg8dfvOVK
+7v9oG+A3ll4mXjsv3lLOWjZEMpJ7Srq6ZXTLvrniiL8/0MeraSHSEPQDP5rVio7vAXfgDttOrsk
IipwgTfEaTu437Vh94DD/hrTvs3nutZNG6X3EM+yL5Dqf6KlYEqs3tPeJlU8aZeODt3yXZ2n7ury
gcKLqPAJmPDR0CeStKZc8ZCBWbqUa5ExLqxf7ledX84dyaRM/DVAWIuKhRwwDMko/FPMsdPbSzkf
6Xi3Ou93KEpat/v6Ur3hANX4t8hF3fOra0niqwMpesqOhgYZEQbO08rTsw3IH6BOkdDTIB7s2O9Q
Dfh8Dorl3CDM5nQ2HLOYYgbBwsJl4y4jPgf6nV6M6SJrG36++3OvZ37MRUfGeO2m2H1DbBIXn4mT
O+dWS7YKf96bvleBeVeQ08SKNuGUxMq9n1uMtSHd0YeEull1paCNzppwM7XNY8wRvT/P/wbsmu3f
vYu5O58qFdu5qBLW9I9uhw6z2eU9LbC2D8vrlTTBPImgi8HRGh91vmLX2pdTj/Zb3X9uHIpB8zuK
ybV/HzpHkI94Vs+418VxNRbWQkOfYyZ3SFJlQCJWh+4Pe9f2Cwd3rdlCZAL44pthF8aDl5nkg0FM
P6JhxfBzGmx4tHAh68NvEgJzjqGkq0+ZppL9edwvfpSCd/zKVvHP1BQbosTt3sWc1XpKNInfgErV
E7l8fKU2vYFkRHwcV2M5JuAV9291xJ8PjXzQ80ZvdsHQU4rHZdu/tD/BkQ820jL64ybj5op7C0bJ
iRF/YTyqnpVYiE/GWsOZGRm8QBUFdfgmF5N7OAn4qyXMaYEaU9W+m6czl2SkUXCKQ5mbTA5rWDw+
S43t2lNJZBuubnRLy39FFzbXC561R7SA4ggA4U8rKQDPf8mI0USkcSf1FzWD/xo/R9IM2QPHWQ1u
TdwoXvPfxlaj0y/f5+sq7A5ru9nTrqu/yG2HfHRdqzMty3NT9nvGmp0zYDI8gjBjCbrNphg7NKrD
AYWLCb+RVinPsDBrC+1SxDcNN3JNZgVHiTLUevajzqj4J0Glz3un7v/b76NV1BUouamg1c1lc4aI
7rxTrnrmggxYtOrmCP9v03vvYZjIhaya2d+GVI/cJkQCvPBkYLbnnR0SJRSIXAV3s7Au2QZmp5oI
eCXCiLGPaC9wZJKiOeuOBGoBc8rArRsAFzEnU0tNiidDDjwoNi9b10+SEnv+Ara3O9SZ1UippeBD
l9d119jrzdSvcShS1eoQadutBq75gQb4amEpFdUF6LVxxDemqaZZ5EvdfW05Mo9e9UMYDlz89zWS
f5i6tx9pKF7UvUt7UKRCJH8RGWvGoaRIJjRR0Dtk6wUk9a4b8PVill6EIJXT+Tswg+FQmhBo10FF
5cJRabKIsrxYQIraynKkFRlDF3HbN7X7arW6nJs9ZCzxbAqt9rIScikSzWzd8O9H0ocLJEx8wjt9
YRqVcrkLBvXMSOeGbaQDKOJ7mvV4kmvm/+jlRfs1dTGCEtdBX4DivBLCR6g5jT3ny8fnCu2xEmDl
qbYnV0dWvAb6N5EjKZsHZoGFg/zgVeF0fE9hlDK2EqIMgzZpWpfsnVlvreHBtEaQMgXnTB1Y7OF1
V+mSsp077L6V5N7s2livfImuKyUqF7wMzN3Ozy1e0AyYUgtfdp51F2Z++zTLmLbwqrDzEVGxfiDj
G6KS8iEVjN+Sdp6X9KubBrdyqUrftTlcHnrimE7bVgdGjaGbrVZhlQOe3j/ZUtKihe5aT+kImEos
5qU0L8WXwU7KNz4S5QofKXQvW5Jd3Ki8Ef1YXdh3kYe8AoBKWx1/d/3zobLYiDBVcEb94wIYYIIh
ACa+AAYNDV8nkVhp8A1lOSGu7NXqZucim5nfZuqQfkLyPi1zCFJocF+0SfQH2Aud4ev6CEFUK7hL
YRxUfks1qf6ioDCp6TxZ+rxA80N5so41hrfOGx6fh+Eaic1K9U3gA0GlKSOA8RvJkHG8cM+BaExE
DROhcYaR1ScV4bNHvU4FYsQUtqX4w5nzr6Gdi5c44hWaPsCBf2++H1hBAynDd51qrUsL2Tpj88xK
syR/fAZ/kSNTjG8ltmeXFwHSgkx7rbaNgnLHyV1R+slnGzMj517r3QMebnk37lZp5G7Bg7Y6mkSD
oZtfbTOVNzhf6ov7VwkH/cvnlz0ed9Jy1H0EPUa3ETCYtmFcocXw0oiNswge/paTKAYr6C60/Qmh
GSiRf1NoDkTuljH5FD4IBytZIz/XLQ1Ml4MIyL3owhqMhTpMjNpT0c2WDAG07+upXOerYCp7syrj
aIA++sOPiOGNtDFkXwe1heV6eCudfjEVipFZ3UKIkn997dQ446tZmkYRFac+iGKFGFNHt8Cnxp3D
/UQQreWPWEOXtb/NLqORfCSYVcfWOfkRIT5pn0ZU21oIH/EjOjYZsT4gXhqqjU77Rrb1mGBv0b7h
IiS7M5HbpaDx3gw16uIVbreUumCIfdPCti4Q22LvS2DOl9Wc14xknJIENbch5+GDhtAUMI1z/vvT
3AzSXqBnAht+r+3Rp+k+6GxHaOwkf7cOjv1qABFjtm892gr8HvybDBN4HPFP5gTRg/nIGySUsF2h
E1LeP+65VaPbtWG1NxYXmesfGiUHi6XhyNlo/Lp5Hq2WJ2XwGVsTfRPI24RP/inOOvChC5Bf3rhw
KpsYJOXZ0HWKm0qDKhs4SUfRqdz5mW74l0jXsIuc2Y0JtnO0bclOG2RojzZYoOzScB75hrOaRy/o
K32amSyCFbeoUqIivxw6VRml08SWubnZDkd7zfYpONAWVWf10KIdueNq51nL1p9G1Gh/AtdNocNw
sslii002DCGLzCRFdfLqLKnpwVCXWgex0cH/8mrx8KnKc4S3OxOe+x0A3kIFkUwDKqbcqPB0AjcD
EAVAM0zQrUo6IoHh5hQH560rYEPQsyZ1L9wTxnEo5NyKLC8PekumG6vaTyQGx5kf6Vpd74mQ/b5a
EDviHcaeQgm5PuTzpjDtraUbL0GJKRBy0ze+TDJZ1n/Q8ZS5ViL2GgiPRC9xvQRJeKJT3CAVF2IG
dl/+EXccyJ/ViBzo6QqVvNJ1c/gao4lS1TSdIgyfQfNnbmZIN5c0j5tP7xJtturo3eBSYnEjKMYc
n8J187I5ksKTeLzOMwdrhV5N8MaMnaygWnHKjHA3liypnTEpFBp8MIzwT9BHKGEhUvyRWDTm+gee
Q8LVhNvC6LvNGUK5KeXWyvlkSUcfpsnq5MuTGIKsOQJsLWfE9r4sQd4g2x9LDHGpCmJZfXAV+pXm
RzxPYIXHpQPhbItXSiQMACHfEs98AiWBeRF34z87xY4BPk+8/JJFtbfGfeC0Vc+je4BpXYx1mlK0
JokTHd9iSlESpfBaF5Scgat8kKok4yu39o0IYx0tXoVuw/sZgGe6B6PS6JVsbJp+KLPdTw4UYZm0
QmHfOCsLcrBHu25dTTCLjEAAntuatILb+w6fbyqQCky88Wo/4sjTbMTKMZLnaJNtaNAGx6GR1uNg
gBLE+kGi+vwOXjUe4Suvxg8N/RdnkOQfafxmZtJaX2VRH/5jMJyJgE57OQ7oyJ10zopCIaKFyp1s
59uIZUBp2zTt/reqeRFrEKvEVEqcSNsI/99+glCwXRdpOJhKs8tVQPS8ux2X0DWYdDF5D6PXnxyN
aS7EfVFrWmOc9GM3CiFCyAX6g/HQTyvFmfFjiTWDr95FTqaXF+KB762RwRM6MTv7VjVnvggW8gVU
eGs0UamvBkXBch7eddZ48i9LeMZjfuRZhOCPc2fQslFiEP5oER4DpgMPLzOJweLbY94nnIAzzU29
fsM+nlFC8EeP+OszhLf1Yc3rms0CC1BrWtYooVgPpFGuiG6Ov4kgYGYCfsxTZCCx1g7+iyFKC1Q2
WSAkA2TjyHdH2Vb2ZU+6FlDiCF8ZVNjkVE3a9YFEIL/OsRbOX2QwkGAjHashTrj1AcxT+kh1ownq
o65QLKkmQ04ZljLUG7Zrf4AQp8lE9BpZKuyUybfRrAGvgj22DM/W3jJPP4HNcxUNHPJewvjCsFIz
MAxkoHeVfxK8jYG+CNJkzklFOFB2EKQMsReG3OmSftsEVbGP/DE+UThrDYHje3l91IykPy4Cu+C0
+LYdnUcw/nQyUyBMbzRMqeljvBrtvPXT9mw9EXhby8n75+8psJG5ITWsmNr5NLDyoXAowwQ6ZLE+
sqLpJFal+MmD0EEiSMdTOowj7fhOyRwHxLxNyhhfFTxXsmORNwrMZqaCzfyawIkpdhUUQBAMBNMn
4XMGp22rR3joJgr89x62WYhec6S+2ymBFHOmvz/ez6WhW4uorz4rdVfAt3oMj9hxGcb7Me9tOPpT
mo/Wn7iEAai6SMqpPVDJxcWPpjyllDx2hX24OQpoT8yeF4yfw5/Ynv89YtNwAokKcwe5Vh/E6u4x
hFBzRmNIfljep5FhRipCIeE6UOB+T90xaCguZ3MCAn9xItGGefZL+qE705PbNoxJMaAzA9f0L6WD
Z7fBxs+MsOEp5jFBHHIiSohX8h9SPc4NNHJdnVGQAFfesomRK9+AVt4YfenOdEaX01ex/rG7LSjd
A7LTgf+C6T7eE2+qvdR+284o6yagY49w6DazN77wI3fn+J9YeGJGXWuMg6d+UfL6SgKFuk1pMZek
YwL0C7vmN5KlkTRxet/7OP1VNwGsUbSonjHknospr0RE8zKyCjfHtBKzmZisv72mH840rtrKpCFo
bRwbSA+zp2qcgsbWEBbMezFyoEJq8++rcmIAvJHgbKu5idUoxbjOnZ7hiiMwqUFl/IwW2zRgHD0/
uFEJJk5lUfFy+GUwKoDRZKXvEEm9PTiCuXmGmd5OwR0aVulUN1JpCtiDGAgkynhJcGcByLtaGoPC
JiQfx5PRqm4E+3c1CjJhDq2C/YRRnf1Jy37pWaxAN5R22lOi7ouoIvzapV2t7uGEKn8Qe2wGprz+
ikPrF/mBfCCgH3RO0BSRm2AqXnh6dr2tTbZkms8UKpStoSOTrh+i7fe8flsu5k8wbGwjhfDS81nS
gHLkkgpZO23z2FwiSk3TqIVD8r+390BvquYMQb8JI/EMDKCo93U0yGdLBfW85xIoB2o46zjEAgew
CX0oZkSnhc/OtnotkaQRw2UVDWSVzRrCIQ8WOuxsFpTOc0NznTbVQNJZTwxgpvfFZUFKl31JJCyD
1WFhLTVK/GqMn4pBLURBbhA8XyMpx4WKuUsKJnQUrW+xZ8zOuIIlrXGc2cdJzoBKVMUBIfFJuZ+f
fZqzXDCpXKwg7TctjF5NlREUtZLzTk2NE00xwaOvHqQZvAI3Uqi47kuPLHrIjO/1aSmgaPTOtYa8
sp6M8LLdflZNId+U7jzt7kha7z4glfGaMyQIB9NkIoSiyChOkHSpim5h3K6vqEaXD4s9KAy1ojZ8
NRi2QF9rCI3oYh+n5YXYt5r6SDqD1szqdrMVRqAi7eeBAmj1Pgl0urD+q0PqEKYSCVsf0/ird3JS
XUA3qAiJ3kD2NUPENxA8WBYwcaBH56flxft5jTamrH5AFNAw6uADiQkQsvLCBT2XRi6BpDfboPSb
tDTZqGKjgh90fdiB7LBf6zKrX682JDG0mbgMhOVrwHw7/cm2nmegXoOQHBRJgvfi66QxPnjl286M
HBrZTYX76EaDIk+HFbed7u6AZBmSFx0Xh49WgXHEOAoYDUE1raKFjG9h52zj6vp8Fk1bfG1m+an6
p/KBfFHWIUBAt6UaJEmmirBdgRt7N8xZXJYb6bK84Tnjv1qWalFUk1dbQr0DTuEfLwekFJIERuHG
rm09pmVPV3i5glNoTXI21UVRJ/kYn6AiQcbeHpWkqQ0HypJ806E1/kZv3vslrwlalf/dfDKMTZqM
rQCQnXPJqJi7rwBasMLMcE/LoJi46+ca6n+nWiXfAY+kE/LTeA0rQyvCuv5a9sPDUAKCSQWz0uG7
vIpu5ZCiFPqPhFolUPhYsYUSkhwrGeKvgnGFoBRWGoI+B1Xxaf+ZGdH9Qoq6BBVuDq/bbu4x1MZ/
g9WVRmpoom8KxHram3cv/dDJZ8VeEcMnQ52gRYN8vrmym74IZhnGEXm2fyEi/xpb50H/xmKNw3z/
+G48rJKUOafAU+/FmpWdOs2YMjN46N4IN0phfOz8/u+hpMa51CQh8xjJIt6Abjxo8e5fKLFnmFbh
3hWmuS1OFHI2N28RVH+Hx+/T8gH368qRqxhcXrwbw67bJ+x6rd+dChE8cm5HTnV7DanZKBNe0ZB3
81U8A0Ynz7+UbOlZIlDlTGl1T0oBXQ8J1J1SLUc8pAKirBbQXfsbnFOlj9YFBAr04MWxY7fu6dgg
Bzqc1VwaK2dUuuXvfF8FswOt47dn3R90l4Y4uaGdsLQbrXXpGynQ2mh3LFmmDHb+k/4OxOySwqXo
P6sxbRthLazuRyiJgY1/FXyjMPqi1So/io29yDp9LUnOUO90p6XL6Nb8BY1A+J0J0QxBvUGDynn7
RSq1dTkp8Odf4dCPzX4XOezrWHAQ+1FlXtw8PTfmUJnuUhbL+ceSaPRR2KlA75jOcGvunTY3XSpv
uOTmvFHY+Aj+52divH4ZrZ2E0rygqEDhKsWfKO3TLh7M6tIITbbjSrmDYR4KGb2MWgIY3loTWYU8
UMNtyJGuBznz6JQJoVY4AhHXQPtck7Fu0Ewd6FGTKsdEkw6CbDw75YcoC7Su4z9oOwG17W21H9jg
XzXEaRlUQPOiErswkiJ5y5YdmqDoFcm8eBqaPzM88+pRg10cjHzngeDgYMXx7X3tBGu26CWTXaDT
Q2mwO6cLDzKxY/vrP9+p8usmDeVktBHZvyW2IjeqsdFOx3tEvQWMx/qPYUhfqerZ/uc8bhTTtGpF
U9YvlNob8krMd6ZwV3P6pDWpkmg7zAlQBjLgG9CRVcCBfjzdPBDkc54VsD3ptcZcFCCmltUUFWCG
sdBtEAxR8545oznq+hPZWYgWd2AbMf3bJ2ROdukMPjFvyPDavfbn9OZOimrdETAQPZtb/ZycsCfp
wRrAjUId5wyEDoWky9CGyL342I7r578DNgPBTaeak6KuUS+76PaRHTUfr6e0BgJ4+AnWb/YRNwWT
5F+RVocHu/JvUt6pHIv/PoltNNetycbwvKO61rQtsygycsQwFX7FXcDk4lGMh/H/pJsld6EJZpds
AbNSXcNYvYNpNDrsLsIAs//j9FErUx81K5U6o2/QrPMYrVmYO47Om9OBpkHqXofNFcexM8gzXR0y
bfrlmNDPZCWCOhLkv3zDdKBZaQ0gihmJU2GC+L5mzXE/xjOmVWpE9cOrQdiuIJbXvPIJhPce6M0q
7gzvh3bno0gCuOjg7FYTui/8CaXW7+Y3xgCGUGnKsiLfJwJ343NKKTw31oidE5ZxcRSmYkmiFY/o
ItciUJg7Q++LnQzF4Km8rPBE+o5uUzMjdxs1lhqmSqhcSzBrLjYIRGBZeDKs3CyIOq6TifBZKROa
H1MJixJnifuFzxPrifC8m5zXpyM96JxDz7w+LzeTk6B3bCWWceePlHwiWYngPDcOlOmtEjovCW7E
OakiqZKfSuuJOw28P1BGjAVLf/pJlswHIUglV/Q6RdC/vNACmBwCtnSyRfBq0N4rcBs4qhyaLY37
p9LjSkNBUXHxh4TicskOpNoredncSEIk9IEeYDTmaUfFbetdCsOreGgcdQ6V3sIhyA/GvAOyPg62
M2kMt77hBsn8u2KllmKOT71eV+V2cASntcCXnX4jB48TvA/7SohpK/FvndIDO0J9nA+alSoW9iWV
eZO+OrJdimGOuE+XxkCplMXcj0JIj79BNSuZy009RW9XxOgek6CqX5nitiFyceilvj4ir0po0de/
kURDPcEVi9ZARHCO7s1syRKzsxZ+C3YOPNymnDp+KeyP8XScMLwTTBH/CCJg35Ppcst4lJvOUPnz
AIh8roIQ/nQIkZlPo720eAevsi7jU86Bo1FW0wrkOmEjb0UBTagGH+Y3EixJGp2YCIpjAgUdhSb4
G2nPSS13OSS4iTyJHH5a/YOL4VuH1L8a+79MhQTyU38Vv0L7QK91yH5AJ5P8phQaVDh9VGotHyNP
uzwnCHoEgnIx07nvQK83sNlI3F5qIY/kiYkdqcNQVe+SPxksANP5uCKMExvSqMiVAFO7x9yaQacp
ZVEF+vUoJTGlHVbBsOlqpyrkjmJec39J2T+xWzuay7y2tr8rzNV6X+iPymMhPC/xIOlmr5djqU3E
CD9FwnWEJBxJHK4FWs2BGCjwr+aS90T+ooIjG8xO+W5eFBsGgGn4+PMg99oxgxBk7N73zeD7xIsy
S0OT6U1tKOc06wvsx51HjpITYt707uOkGebPUKRQYpvu+QoUG7AEuBGyCyWprOJy0a34vkiRnHVY
KXTPklbTbcGzMBaYxG38Gz1W612aOyl/5CiE5NcVSqnSi58RLdnboX74NWseaPDC16WJjIQw+dKK
gn7jIdL3FDosqrz+Qjs57JS+H6Lz2HxnUWUeVaDYNX72nqbcQ7nAfqMMDKe6zEjipBUDD/NvJcok
btKkQ/wpprYhkfZ1fKbbZ5VMqX2ivFspFDbVcjcapFI0cHKiYDxlmFudyQJs0M0IgpVHaKyrLXAj
9hWtp6pGs7IMAkWV3o9jvxb5/D22nEMID+/xSRgKfCIdzSsRC1sYG4MAkgJqU8Q1YV045C1P334V
3QZrBE+KVqiFIQugvFBFdppgkvrHfhVjmnuy3i3UqcXtDSEAjoXq+RUHAMo8q+nCWGjK1nmLYNNM
dxfwM3Fu8caRChC/1BTfbQ/uuEysv7zALSYQEQY2xeck35QFesB2pGkd4FzidtLvjlX4SyYsEAEw
df2OaHnHInNG6dzgtlAd9EJvOOX01ZDuYgCXKUUVEUuewCR58E0k/9xVhG+Rs2UC9ZGH6IvimiJO
IipaLasVvlc4pzznmtFtegodxm83uFXm1uaiWEmlz5t1VZfgr43F1GM3uqrqMNmdPpdQpn0qT1L9
G3zCnjOCj0aWzBUkew4z5cXybB8MWOupJgxQLMe7RoSYBgCq0ZdDssn7m0Tyxoq/XI+SWB4nIAfp
vQP7vZDny8LQOcx/auVvgp5QeUihLXBgP1+Gz/rvao0MmLFF3uU0t2UzxVyZUmTksBsHRzkoEuOQ
MgEcIXWrm4pAaZFUW9Zk1uF79DVShblbhLrfdDvJwy+s+p/61nJCICSBGACo3Fa3FxCpkizK84oH
vSGAxQUiaKC978VJk8kyc7DxbLtId3va6vtMLlhXpwiNufN4Zh1WbXulf+r6+uVH05EHW3+DeGCV
2qc/s61oEXSL4oB8ND7/l0yPNc5tHmfLPlV8Rsdbj66YQv+x+RINdiESlGrfxRws0PPuMH6a1GPt
NEaTPWnesvXJA3vCy7ZhVdt/mOusybcRObqTbYlk8ODlKjDnSi0PScbXheQLRjx583vbGWo9epdm
I3QMJ/kWn5UpAe8Chfg8gzzhZI45vxAF+GU9uG9VyWmVIvUVu/XHZd4UXz/ALCdvdRpQgI6MgtNX
AY+KPnf9YoC11eso66EqQs4WYGwUTGtNGkgM5lJG3+ant8cgZ2jmw2DnnUpWkzNiVt4KfYcckQhP
0HgjlMbr+q9Bwj+R6vPnFQdYVBb4EAuAq3VkbMG7E2Fvi6Olz2xZx02Bbz017/WvubBwxAtq01F/
nvmZ/yBIIdNH5m7Uj4COGtPfl0VaRG9eJls3H00PTg3+NwrfTxYHSPKOnk/wZbtS6p7l7eYxLWa7
ygtpZM/mPj4398nf+67JJ4VWzNMWLhVSn09LiOety2xhe2WHY5Jy2MY2jVJdIe2QvqdtZCDxtEyz
ih8tvSt9Yd2R0RPM+v0Tj+8jWDRedLlV19djVvOWFdvX9ik/iuSnHK+M+QDs0PPiHg0DdVNJ7qeJ
jvtMSHm195/4eY9lZWhV0vgx6ZLJ8QFk8koaRnQ29Qdp8r7X3qBBSPOEG03bX/BJ61n/DqxrhltV
d1AxFqjwxS1z/fyShrzmJTS/JcX1IdiWJ9RIolmE7mhc9DFUQFt4E1RQUhaO5bHRXSBj4Q1SE82E
WYUd4NVsd4+STsv7BZ0wfVsGB+wt/MzMliQbcOMjz5s46guVJbgCu5BxOUfGLcADtEBznNATJaak
7vlfLz04ftH1y49NH5FdMJBV0SluGvEoJLFQQQyRSH89HUA7Und83PHPj6SNCGtyjBvqUdoONwlv
1zxGnlQLiElx5VxTlk74jH+/n4OR8xopU9orSJaiptF4CcOen8THOC1o65+BUdD/kdcgQwCMR0IF
IpbEid7xzAFBp0mZNG8px3Q76OV34YL/q5dmmbZ8HsYy6o15wlqu2KptpJnyC/y8xmynb79tAYfM
QYkPILJMumNt8NH8fgCk627cr3pJKAHYaSVlnwJUNnTzCmD1JNKUy+eN9Q8x54eiIPCxgArDRQEj
5QE0k99NnPKFv9CqsDeNMKZFuRRm+Js4R17b1n4Kt9L4FG/vRlB4xYy+AukWBHxlSDolqPCaoex6
H5uHoH+Adn0MwX7nZyH8o/7ionA2aJOnfRTYzubYqkX32ChHPJeIM98VWnH0RdIE8XOLgg/rMWD8
vaxbo1dRAsxQxVIS15tEJw/IE1/lEMoI3bLQUWki50WM2glMet9CT5xyhZGTBXLgIo9Mec47NeeJ
Qj6BCn7D1doH2FOFYxeVMH4kFJgp6T9b8EgbsY1mi3FDD8E8NCFbXsevQO5EJc+ONmzZk/SOh7P+
hKXeXtLUEaMWrtmu9A98hjNfKMwHPG+24WCqNHhbYeecRIld86Jgc6s27FTO4qW3WW4UUpOyyQmT
wZlcKlySJtUiSouP91v9Th9I2l/E2LuOEfLklz+yqbbBzXRcUHIpyAl8tM2lDozcwenEOITMz/kT
uyQTgY+hKuqIj65NbyNYwZ5vvlHB4o45MKWR2FFSwK+1E98hJ8a4b47TkinlG4ifyVCAo54UZ3Kw
l+KBiXX68RgCNVPNNgtE5Vgv4Xq1hY2vGImj+epWKnX6rv4yuuWVxaRzTG7frNhWBPZP4KJqPI01
nj2XHDXaZ18uTEhNo7TrHzZ2JWsET9Kzu/w5tdfIZ4trRrViWXFsZZHPklL/rrii5UgVJqvsWHAd
rHT2/vT6Y3FVYNcL4dAhvdih5z8U1hWwd5iVzpY1slDjkXizIQFlzEVq/xtbn1LJsYUmJ6o4zb9t
AMv+oSWM9iTVZ9WNGtGhp/uHfz8W/VH3KW6OxzVxhdDwXOjSY3rHpI2zSPlZgd6E5NcBFwj1POGd
9SabhpJQykgGQ0mT88c3pPqFhrcZFFuOLRXyu5+Oqvl9TT0BxK10bNuvRcNWo/Kv5qrs/O4j0Y3b
BngNlOq/6t75dMaxR8czaD4z89LaPXphS0voFaiQaISHIQ5KTUu9ux5KQQY/vzpd/JM5UMGrEmVE
qmX+qMqA8OsUGeKYVnBGe5YL9mDO8AFVLIf93UuDUds1lDc0IMZFQ5cAVC1iayeIMg9sHsastCtr
keBliv/1X5kMSNU7CeCStxxpyncH/boYk5eCl21LASPg3zlx/YFyXoLov+ch6zk49uwN042pfA0D
UVTup3ma5+cfw4bP/fykM32GSqQfa3Ofn9Ca8KMFm0XEqHKuTTgPq3fRH9N4w22+SLHeCUiJfhIx
2VYgr2sqGHMF9djf5rEo8I+wGmrEPB/GGe1Fya1eKPueVQw7JQQHHdvEB8Nqr93s7hdUeZ0XCEoy
P1twlwKnBuadgFtiM2hmNcEFby1Hf8cHlW77PppqyFSspwvKg7Zvg9megYUUXxLaXyBi74kSJDGd
XeT/f47q5BlWBA7jyT7Ha6eMf93HE87IaFrMALhryu6QTrWQEa6v14BOgYPDK1j0WZcXNX28DD/F
BMloowCwoQAtPnrJvC9k79hR2G7lgPRU7SIPKhLZ3oeeHsU63Mof6nQMYgPWopWuV1QlANafHTUu
DxVzqC3J8HwW8Fz7AHryHbZkyOZXqoFV37nHukHNYE8zZ6Vn8SPC3rI7ATSV0e9F1HDir7RswQot
eUukm0GLjNybejBJyw2Xx1rlSAYKg9Kz7szEJKErb9pDVHM2pF6qO0NoFIk+Nbs1VG3yba3T1CID
+rhmq52N/SktqYFpwZSaOauDHgFyRPNBDiH0xwB9INeZD4MmUEsKe97Bn1ZDeSedqRFHTMrBhStJ
+RwI5xk4XrjqWF7qouOeCVcG/+Y+VKx1diL5JkgUrqaV35Qt8tTAKzQieqB6KIQyl6lnaKM5FJCx
KRF0gJjEsWVdKybdftQr2oVRZz/D+HDSfJEUqRsvvHTaGUV5XlR+07hx5OU4xb/B7LjoBFTKjDoX
Ck0deNWlhLoGdOT4QoaEcg8yqyWpU/BJt1fR/YCIR1k/S9j9M5dDamQu3GAwFAJcvgDjx6gKCxqq
KT/xVDjHiDFyt/Tec+VAdAxKD0g22EcFVn18N3gO9Ix3XeVopXlxULSVxC5C9oOYb1ZG3gzwyJe8
zye57KOv8A84ZxLN8DZjKVVPnfaHDY+MkEiQeWu+vHTctRot+C7EnK4Pfeqe4lUUSN/E55iLg67d
OmrjWFniROogmQdvRhFKNVNakG8R6fVmm21RX83QPDOkGkfaEBxagl26LWyo6cV8iuUWGfg0Aqq9
0enj+HJJhnj9d3Ql17cTd6fTuII7dEU+wLr+g5JrtiiauTWGimzzA8MamOC9UqfGiaK5bDrbzH4D
ncfvRgsgoWxOvI3JsL2MsYMvmkcbkaUixluO2WbLGpeymkwX2IZysDeS+fLC6KjkxUm2fYXpQmry
Z2djwnEoQDilhnK6/4SO2HVV69Wwma922fjzRmhgxX0dhebdijc0wxK+WsyPj4XZF9RjIFt+hyJr
VE0QF7CwxtcijKQpNRIk/WaL7uqN7jtuP5jsUg6NVBkdgMO4S1f4RuSrbzXy9DzNOBArvTTNLhEt
E62LRPznnTGWcYuRgPRw6tMmnHqxY0CYF/Xin4p62fjWQM1QEUZLsyJAfvBHlHkqzR5Wuce6RXAF
U2ieJjMrD6a42Val2fg7nEZYXAPew/IiocUcyXndUr5OHtfUOTyaUHxBQ30EGLomKuE5mJM5K++W
AKaMq449WB4uFw9GnYFlrPegtxNO7+xzzRRta0moWwq6H+P0osZWYzsyV5gLssCO1Qsp7UiPK0zw
cudM0ZTvkOPBG4ZRMIUYKpQPHxDrFVyLPNGyy6uobv8Kqn4AZxGf4XhW4Zs71SLeV1imM7Yru8E2
11jHUL2aL3gj2xTRxbvVfpdNkydWS+czlc/sWsrbzyD1GlKNChnkn3onByturyLhA/9jPEMxI45o
hOE21zUqeXPjihwbLXxi9iI99cSFCFc06hv6ztXPG7FNZOUiCDqP5g9VebtdwKwWO1I7eELvCuf0
hTYJFHnPuqMivk5zZGsOPBlFTqmfypJuCaDeNHbga8aM85AuJvVFpxrA1UodszmB3hiqZq8uvJyk
rJc2WzblqMKbe0fHHvTBexmf/gFNnbpjsRTNLwhHyGiMWc+EHrufSVfiqCju3jQBDch6py7OkBb9
m/g647jhMpf8lixZOaxsHQ6R2VTokidJCAJWfs6Yyr1BnxugoBAdGnERFFei+aelgcOTwbm2dH75
SeQIAOYnTsGC6YzQxArEaYdD2hcMcZS2JJDcAyYBB+NOMa9JiK6tRMyYWwMGYcG2RmNjHHRXqEjN
eJi5KFFfHtzpef2gmaEP3h0JB8JkK2adwN8dSJz0pV8CRUtjSE7CB6w/b79euSXGCVq4PyGg1q91
nJtHp1r0BuYyH4dQD2J36Ns+ZnyNCNUQ399RtVh0CwENftI46OUXknugfwQOf51/6gJwikbcNvxO
wYQ4Pri1xQacXP4VvlKXzqczbZ75f+RSlhURDSOETDXpNBPvWO1K00HYLtvg5Uo/r17ftdkxKzru
1f3A2M0nEAf2WmWxVh+XRBXfTyp+d08hSyoucNWhlPUAm76RRkh75WL0kVVjlOEfOVcIPGJE8T/l
3sh+HWr94R8m4GdIbi/muI2yr7fWp+heWTGJ9o/7dSFpsbRkAhpCc+STvSYw4DypIYsS4JKLDUTZ
fE0v0yOl9+P24/6OVaL1ad0XTyowtHa56Z5VbErraTo87rQtwaAMS8DzTtkpUCKuDBiGB415UBao
HurI12w11YRDi6cCXxeHT6RyvUjwsP8MpN/6fv0E8NRRgzZ2NY9188VLo1xNdyTiaHWZtiaLtabq
pONy+ckyfL8+p/FGDR2zTUUKD1Cj0s7BWfnSq1mtOkmIPsmcZTXN1gK+11Sf4ekYE4ZV/GTF9nXV
TN0gp7euhlHzsiWcwfwgiF1GgQx+WkYUbXIPPw6QPPt6R0kbWyq7L6CBTAO6RVwqoIhqur7dlycb
Deb1HhYq6aPSUopbn/kM3s7N+FhMYnemjduhORRcCJ4ZndZOhMgDv71nP4waof9I3goXBOBIgMmn
5AtzFQMVlyrp8R+V+Wyd+rdvcQWwghaKgfmlBstpCtO/A+oJb+wK5kZZB0DeiNX82dkNIMdc92Cf
9clqAhZmUOge3Qgah6V4Di8jAuqvu92WZsBLvWnuZJZKZ1akwbg4bR5JY8Fa6PSsfanP6rGRNiAB
PWHWuzEUKF6kmc3x6iyih2PPYzi2qQGirMiA/BGgzCWEkuEqhTsv5C65QfcFpkXto7RTILKIkumE
RaZJ8jgep8aJfqHrZ/cEvHBnBO9jvCmpTVY9iZfO3LmRZwcqi242eNh0MGnoyUbDzHKVYz8R1rdi
pPUVtcFECBkpj2SIhyKppFjQtPzgqmAGyWU+64AFib0wt1uwo0MMYuGeTH9GzEpfVR8gPH+K4OLz
xIYQSS55bbsMoV47EyAploaeCrE+kNQebfT/PP6FzvGUganEj9HrtPPUPpRhMf4aWaCtkGaZVTJE
0GLQFm+NQeIsS2sxDvAkWhc4T8XB5x7M1638Z9x1ZGl3Yck9C8DXSTFY3KBXlwTEGJb9T7fGEngK
9ecWgSn9yCqTY1o8+246Di15mGYIvg5VD9xhCk7Dev5c0wAAFnch+UfdOu6mDoIvZ5cpD9qlxxTx
D7pdf/zARqD4azvDyTAosC6AkMFu64gzj+3wGL9zr+Ve7nym66mFU+PygSoonE6C71ji03Tb1Bcs
oeHkdHDBMiH902h+bXrUDxM8aJm7o6Ji4EqSha593tPfYA5bzbxuDUjaXfUhARy8i4NdK7WBsSrs
jCexAZiY96OMDLz+3mBb5TLfsBywofz7gnvaPWp3826ExI4Z3kIQzr1v63A/IRTWa2VyosQwfc4f
NGFxs2R3T1soSr+T7qWUn7CaRRHYBDCEROrRyvpBY3rqOiADgZ3VNe1JPLbrXNtL5boMnnr6jsBK
aGgOEx0OQJQKrA85z0JO9x7m8LoNuNt20jpPF3rPMviOzPTqO1HbQm68mCIpiB0bQKoil1xPgGQ4
bmBWvl1t/frLzvcquuoDGny1BwSQbBamAoEzFJVXWm2xfCEzGBE4dJXFPYM/A0/Xnhw0gCyk6msH
LN780hmdPQl/mry3AvtnnKOwUBiesCZc6Z39WtURDmc8jmDUz7PAV8atDbbfnjXyMsnuDXShSOdf
JLS1ckSwLc3uKlzAATgs8JeOhKX7pCM2cOa3dUnQlPLrs3EbiOotMnL5DAkYjA8tmu9PV7QN4ZTv
O0yCI7wriBU3WkDBISNSFBndvfmpqJyp7MVN6OB/ZKqGQavtCuMEC36QSlYRu5hURUBI6KukNa5/
ePucqIBe51/qQDORF/mn8f8gMk8d0TjrGzLzlDgIVO0fSiP+lomOClCGSD7kz2pw40RjJ/TFibhy
Z0/jyNP/6arW0TrK2DXFU/sXQyMWHi0mfoXTb3n+tGeXHFWwltcTXVhlGUGBMXmlsjjwNKZegBw3
pXG5fHK4SGfs9Upk8yz9JJ7Ip1nRNdQn42DRi7JxAIeNslpT45T8ENlCDfa5HEAUp/uWUDTabL/5
tc613VpCAdg7CPjDcUqeUvLXjooveE9IAge9pzCrg3Jum7Sj2/3FkpvWxhxNx9tsKOKblrFiWAWN
5/rgwJP4FJl0CXh/zPSke6ypGLpTmWIwnmpyq+VsyANSUEBrR6UtqbxghHDQ5Bu4aOGJKbPuduhV
9yrup3l45Jn29JgaBdQJ59TJ2oksb2XEIWKwfe7YK6rDfOj9UbDzQ3fFGOVJY66BTDW1hy+tWQtM
U8SlO30Qmuo6dEZqWLxG6v490G3EibhvQE7X17kGg9jwp+F1rAFsIehwHPRWGfRiEPFMkc6Vt/LV
Dvrc28/enxVw+FkBNZOqZ1yipEKHZ9qxaIyTdwBaXLu9AhoUIRbJnh6nzS2X7p4QtNLIM72tazo0
ej9koFsWFoObPGrGioliiobSpHz7RyMab+T8LGB4lP5W5btcoBmg3WMjm3lgRmtoIGJD+cQ58QjJ
Rke6w8sNqBXTiCdd4ApMQU0EYRMR/IkmdFjXdJsluQlyvr8n7P4rWmiOovEQzuCXL9vJfvtojQTl
yn5a/J7JXwu3s3K5nlguk9PWEwYZ8ZN84EDJRbTNvNwVAX0Fq6tQNu9wai0n51x8UySUeA6gYD8s
rYYemWov9pp2RAYRyHgiolQ116Xld+5AKGAFgFk0mfbBFS9JTDRvtnRGil/fH7ThPxLb17r6NKYR
BGHHKtYI8fqT9n+MVdaQqyoJ2LDurdPZ/IePeOHB6hY6d+7sq6X4WHiQk6TKjJ87mhZvQqCDhN43
ddYG0E+gTChV6nDLD1hiYHnmBRPHXiFyNiICjVs2ovYKjwq1eF9w3fgm5f4V3a4WT6+7z2m1XTH/
tDqfjU9I4HdDgQsUBUaaFTF4/xm6V1EOoJnb2DUhG2qPDHHgzgrViKV3pLaSZx7IOTH7sP/wa1gj
/77DRWiz1bvahvz+DKiH2p6OcsgQ5iCGkvf1GsaBuVFRMGw560JIZvfPKXYx2zmKNbgOpAc5r7ag
bR2Kf6dTcwxvQw9u172D892zP16A8jzO90zx38gFNDYKfrSDl7Zsv3G4lrL5+l1JPqdMNfXARWFB
VQslvBStvZDd0VuQDFxab+POuX9eWrNFuc9hAGLhOznpmg3yiGY+LayEmvGpkAZBf183Aw7Yq4pm
mP8oBNefM6Dzosfm2/Ieoh1QVsaG8cNeNGyHnRWH/BJp1BlV48o8g7wHza2q8urnDqV2/LCP7DJW
hki7kwexIzYGnb0QGvKP5P/jygqNXH2YnhHWJyY3XZdWCHC5+lqfzyaLRRUDwofokL8G9aHLInDq
dUcUpP0UjkgsIJoK+68cKFADq0Gvm8t4av8owesd+Cwl21Dx3DD348vV8prKaRLJ8VfCQMbLMkdn
lA915yt+ObHz0OVXQbK7IgPNeAEAIoFJdCaSNFOdeehwbVCuYCrevi3RDUbedxPnOmWiTt7DHLFb
tgd4Mq6J9gwj+bqh9pOjkvgvtiXh3rYIfCmzaqgWm/mdHgDtPsvkFfQwU8LnC1ClNKBqPG8/THJ2
AcS02O9gtrzzFBBzJPFoWMdbBlqZ/loaa2CNYtGYiIaS7ceCwODi93oO/TrEs9NA/BHWrUJvcBjO
3eZw7jTWhgm5owrJd3Rr9I3paLvssBMe7GbUC/KxmUnCZMxePZF7vkR1udx0/SW55lZfchZnNy33
CBPlXwVBajFss4wd2WAkh8DVP0RptKE4+WkBZFptI2ISIoSdjHiVA3oU0II4vSozjZYhuVHd0M9k
9Sl/nY18dGnOEij00Cn6ZpRRCBcBbJJ4NnroLss2Mejf6CuKjWilQ+UCk9DgyLfM3yzH3onDqpOB
5zXDsdVtLbOelFil3Q3w6PBy2FclBOI5AhZgIX5FcViC1uWaI1ucCyhLmQrBy2WwOUjo5Ir3pk6W
bW1vY126dHiUss5jnc8fYnZlzKof6rvAEhJIm86/M1Q+G57KtYzzMGEjlB7eYb+TSpeNgXv1NrTU
uc3D+fyvWTeC5e3uuuwMNRFLkVrLMrC6KLUuIeRd8/xNFWvTDLGDTWybD1IBYBjAiA3Tqgw0vgTF
6XYOzciFjP4VSGsB13uqB9l8QAP54KSlANNRJiYaNKcBdXj1vqAP2ciYNOzYy3kh01ouSBYUMnzc
FP5J0DSiFfmgw4qCoiT91PPZ7oe8RCyh+qJxqV7bRr0CI3jb4KX6aSwJxioR2v+A377f7nTol8/X
m4pC8fu0aSjuLgpRLrMPZfR20V9TxwbCAqafE5kQid1DK58x65Kr5/CX7JnoU/bE4099G8ESLbo+
sFs12id017BJTTRRjvq827jCxG5lGMoF7ckb3i7mDIGYuYWE6YNJG6hjwrxb70e/LsDvDqQKHlPQ
ul5vCyM5JSFb4cmTnEgE7f8WE3P5eZkYbfYFs8/UdA5tX/yULg0k8UTfxMjDrBngrg5qHTqVxIoI
tLORmOBmZIvLmg1gyk39ilJMSBkhnz28ausAkdK7eFQMokrA3QjMyYHO7OssE+0AoUjFKnklIeZl
+/Z+lDsCHYYV+1QAy8f79WQCx87SKMF+R2IjlqrGt9kTBozQ1Iaoxb2VjOlUW7DevfG+3VCLdR21
GPNl/9g1rF14L/Fl2M/GRCYlzgbQSN2DwO7kLa55vWjF3A2hVSXenlbgacO4KfQhQwmgV8vXBJ23
TGP00945MVoCLrBTV7ny84q8BUG54VGqr4A3CCSdM0y0mYrNbIiHr18GNFSdPo3DAHxu6okFy51O
A++o6/7KcIVbIsGdUo0yycNzk+lFaWC7CzGA+gZ/FwgwBGXXnl1aYwVNUSmmzPrF3pXnKs7vhG3W
cIsYsJGP6J8MCseucIaz0e6Ufb4PttiMIhcq/W1nGE8eK0WdbEIuHaHDf/PxSSyDSveG8xSrgifr
CRa5L0Kue+fdk6OWmYx2HBmE0xPnuW39kz9DYAO11jnSaZMif/LSbgchI73r8q3YNHkPBpqhb1wd
R4Wa/aK55+ltE7lkyflyfWi6LiwfJ1CZPd0+psagvpSidzfik9o7T16t5CdJRIUeOqbI1iaJkP6b
/Tgh9FAwTplSY2Yq0n+BJV7WVrhWPxKjBvD0JLZTSSFuTyvAjGc27nnTeA/ke05EQSeDS5CTMYhW
xXY6AAkavA68dePiE1zI/zht0BpXgvh+sqmYHseXdhVvAz/e8Qr2yPlttT5n+MLjkfj2HwthjeDG
4eVx04oCFDRmlmtCigbxQC+0IXahua5aEzNSbck7m4P6Yj3qtoQCXcMfbfH9ehDJ1tBkWGGBryeh
ZeRXp3tI8gJvVZHqrtD0Ct/M2cLmUIuVANM3ZiuIXQYFLe0r6ICNIl4/a+6f1xfcgtgfhzpWh2KD
32CgS449mF38fVi+C4pU6h1WxLsttnztRrM3G/smGrhOqY1VMgIuTj7graglAxj0F9FuvQNDIzeI
2Lm6pziSDPErWvCAwVivyVwm4yuzOPuMdx5kgxUcwxlskyJnKLZxUX7Mq7NTLptNfcn653UaJWfN
/ASI0b4ljOMloB0XxkZmrZ911AegZP+CVAPZCJJYJ15iMa1mAGBVrBjZnP7XpUMcACQeZuoPyKa/
A34/i8ONCEVarsaTMKzQnqtByC6v52SGlUC1QpCmBMS0jUTqg6uoZpSauh0JZzuuAMoHI+gfdZmD
5gJQfwJq9YysCxRh+l8lpcKtljegEtT1XiUpXJYWbWabThZWOU4NSFqXfIo5QtTij/FNjZ1RcFub
G7WHBqCw7ruQgXHG8ga9iIV8UAPFQdT8WckeQlLFAtfI4Ag4or4MfsFP8CI1ihEst9pYooFN7F9g
Q4V7W/wRE14wsuZyt2XEtqrY5wOQI6Jr+UWpeGIFmi/80ABksW/9mAuEA7rcbnefzFwgz4mqaEjF
C9qd0d9RDCkCk9VbW4g0UeCRpP3DrxKndMzI50HzECiISA8zTII/7BTkRGCfKA9+Azxk2vVBxxdY
9OfAwn6Z3niYvoY0+o3zysRrAjszQIzERbqQ/kaVvyYrtEEjonDVuPCFqrcLzLfVebkJ5BnYlX3Y
YOKY98wf+GBmJmlbZ9whBAS6Fthe2JpaRREBpe4+5XCBlaZNYSy+mh8cmkChaJLit/XDN1nVZs9/
9t3Y/P5vq7lFaIaZ5KpPX/xVebBvD5vjRkgXGh7XPR91Qd715kB4d2SsI1v7vh03r0//x3USLGCO
avKwjenUX3EhIRJcY+cOTaCBT84rYkxDLFvzpnXZ1Srt0+MkTvP4/FpWNVV4Fa1PMULapA5D/O9H
/48/GGObLb8N96MBCyX2fIox4EDKmtB/meNogDGZ7duMEqreQG0De0iQo9C06x3Wliu2Yv4Q9ddL
Xq14UeQINOUtZPukx7mtTdeaQltJERgB7VEvhIryiBHdhqvGs6yT9DREpYId+svmtnelE8RCFmci
43DFMXfdJEFTUWL62aO7xr3KjLAobpF+p+RdfWZH3rdtAWfqLor4uayLwYzJOjaHs/KDmTnKWh57
eCIOX4NFT/uhK8YjaBOL9072h8b/i7CYuHjbtbIchRU20AAV8wN3x+W++havGcncUhzePOKUoWkR
R7vNvzBRyFR8p+po/A4SuON6XqxEmDdfte7mIfv2vYFavu3FpRzPPJTcApVsDH2lfyG7PWKhLhry
iEGOQz48cyMh9WFzTo/HfESOW34Bm2pI99WNILMT9famwJ6oKjcyuDoVGQ0qBtEPV6R0mkN4aF7u
QkWCf9E6x8/81GGGixrFuiYz/o5wT34Hsbf+bJPQguloOAzkYJ1W3yFcfS8cDwPNt3aVbNCVcIRd
FfriTpKqB0ICTdF8YRjOHTArmJeqoOWVJnoRaZ2qOOA1xNd6zvHH0Z+k7bm8X5ktA2Sls3YHkA3B
EdRkqxrjV3sr7Xr2gNQ8ISVy+tkgwP8CYvx/zcsQPp3T5UVYY/yeuc6qyE/m/7pQf3F2hXBAvzgY
vZjh+aKNUgvEpkSxK3BcIxCC6NwKMLXNekhXlRV8lCtHfekO5vYqkXocX2tc8yaAE+gm1CCeJE8Q
9Za34uP7kxYEh+vg2GklCVYyiFh6BpPDJ3bdoFLpfdTRA19rL1Lukkopbv8EhAC1PS4cbe0M5ogT
v5KGUmo/NnGIw6WsHaVCjWb9/sUcRPXNpFRNWyNquq7/YsXoGo6IEfr+k8+z+R7MyJNKFDTyeIgF
B/7+rftYUN+FpGHvt6clIuudDgNB0cdpN2r/mfPwB+G5eiK1EZ58pHG+nUoTNOgFJH4c7qQYKQdn
7ovCRxrQivGZ6XoDpD4hyhFd+CZ0EeYPHqPByQvd+3+G9oDOGta/5qctD76UOFw8zurv6wXk1ROm
5puOsZAvENdqMfYOw+kDcvHm+W+7hWSF9XP/Mqu+d8IvO/agmyTNIHpNzwS7xbdflZV81MiUCIzt
TjflnhUyK8+tIZlZuOddLPLl4aUXAdEuVYQm636m/aIx4kO2TvLHOqIXPVZCprCKChJ6gODJA9k7
CQh+8MJZ2v3YoDFs0KIVRR2lg2TjzvluDuAMAQA0BUGj8yGCJ2yEd+cszbIeB7UgdU/+Iwcfu7rd
c+Ur6nmDyg3cvqGJKfRG3YBfCRhhy9CfsEO4bu6hvl+TBlDeztIqHKaiJ5StGndCllmKbHfGwitP
JfyxqlFScze4jaXxDTIp6eudDRbyZUwKDOfhpLvR88j7OX4oSyjaISoOUYAJSBcdOa92MDiYcKON
43t9yI6ughu4r+i4/hCxLEpqlXgrwB1sw8R2vxxwXbfo66Keu2MmgWApJWENFvWqoP0lfTdp5R/H
wwIbAv1V8ARw/zU3sBy7hm0lNfCYCbHA0B+7ZzZX+fpA2HmRdp3LoVk7vqCQYkrfFSSI90ju/Voy
SL6MaH8GFdqFpawkMPghPhZqMdZ8QVLmjROC4fxRHLv52zez1Fd721P8PxBg7tOLGBNrKzS0IQvc
KjAkzsPtqVsKjhAG7OyO+bFAtAwo/HONpFfrCdgAZcj0/gEawh/NWbfaTIL2LRgwPnJLkfV9Hgx8
o4CsLpqPsXyNq269mIciB/wHfXmpksV55x2vO9NpjMnd4/SzsQyjlo75o0ZAUw/+sOEk2nTUYKg0
DtU9kRNEXpMvqxsA4bzOIZmz6N/pjIGSnkDIDk2LaIrTuWvm3WGb+jkR8zk1Cyc/QV7PfzHspMzO
0GV3OH1XMXSAu9EpFeZdA0/5GTsmYQbt9r2X7psh0HldoU/g67/aE/LeY0V6qrkJXzNCg2+94/xb
KsNYBbagcHGX0Pre0mJ7HnO3/b87PvXU7TPeWxVxb34+SVkqZnY48mNuUfGV5w2o86AGYwo2E6A3
7NPgbF9dkEkaJNjucsptBfp0FTsx31OcPBNUlh3vLkvBP6HKIHGdFFnXe8CTroZQaSlxyefLNpTV
kVUjwZNVZ+1SCjpaObaGaXxBDnINU+0R60oYWjfl8RD5EooHbkZ0A9RY0Zzzes0NKeDpC8sB2Zxc
LCJ3dBIufm24eUGQzFp96rAzehD9jzckWkJT8slxMmRoWOlf15X9oFrVB6KeM19WMIY585/nbTlW
xdfR6F0RVfOsRWayQSyfec2yg5OA5IY36sF3sq2xqO5c0bYVRdz2RKD9DRq10S/QIWkZjKBlGfiH
vUoypytAxqWo3u650rAhl1v7Qi+gLPojWAWlFRvf0nkHBG4ij4A0o/SnHn+s+Z3mcJhvWEIglIno
N8Fu4Rw27MpkLS/jrXU+5Sc0N7BecKu3P8HAy6iWkMA3YYr6NxQKqD6Trad52LdJYwnPD2W8/1cy
EruSsh0GRs87XsdvAkMFRWDaxaTcWvLmSjKpddrgKrAyp+w+vawrQbBX5GegtQQRd/mM8it9NMXB
oVX6IccrvsApQ7cSuw5DWtt6zhNtX3feL/0gP/oBSAto3CbCp01kWnE4OfGCQjrsNs8NtfrltZgi
QSYSIDTu/JOSml6SJC8PYxKUvRAjlGrURxoHzYgX1agRDRv4DWDlhW0zON7c+0/0y+pAlosRf3vY
qexwUhnIeDbLXt1UpXUZ9CsLi3v8TVzEhLr05LYzvBlvZ9O2gsdzDZNJKnDFW7hQpZrzT4+frKYj
Rxm38BMqeus12Yw7Qu4Vo2eBBfQ1rxQa2PEMMD1olT1tUxw+DyBlNNM7dk/ofLPEUgBFKb1ht27z
5ndpUt0iQnULX1RDpRIm1WWljuQWTGGYSyNBUunkuvhZynNRg8WHlnoCg6aIEPLMoALzpCW90rg2
a24YUJG8Ety8Mh8whnKoCjKeBDeWew5CtrVEzGMwBT8jIMHvyf+9Q/aa7YKOlGN/ewFiZZMl5K2O
RIOC+dalVH2XSpNV65ByGmZLGAogzO0LnDJtOg8lTuf+ZZKoWO3BdCmRnW5ZaTgVk/mZydQteJjs
XopS99sHS2lopj8ETJiGK5JiQHsq7To0BF3tGpN4KmfxgG0C37Ved3bVqT3w0WpG+KHmXbOkyb5w
36WwA1k4YvVkZTO/snrzB9xymonOWM9nk/roMIxKJsomEBng2w6nTM7+3D+wH5A8Vni4QaHM2qsg
FxKqYKYJVgQ0S+zG4YaS5dVxj+B3/6bVOWvWKIleIWuZ55lh9yMjWpT0HU96gXQL6sxcYQWwbOgo
bdoTqXki2QbcVKEcSjS7BvvUPsaKuQemJLNn0Xr9MBKtDbWfE5jxbfdrDe8eNR9lIl/PVxVwTp5U
InObk1i06ym7+UcHgtktBZCwDh6L/TF3k3k+7OdxKX6tuEFPLB9IakN4uvVT8jLrymp1qpBPiY3Y
UCNFpDmzEiYmCcIFPSSL2vsPLnSFg5ekqALys1YHEpL+k1xch3yIVbU4vQxdiOcbJ+EHsZxTrCdV
b3jDl4TDVYEn4udu1e91v3Gh++5NLgCLVRdy6xiZDQtaqXt2f7GPBXzHZyeIydtMGBn2v9USQQWL
Agc/sb0iMH0u6GN4pTmTq+rf5WKqYF1FPR3Vy5UfXVzP4n7mIyrC2PJUz2yZm73tiNFseKPmnjn6
J3ptj4W9L4HJMsDm855VImODUWJk1YalDmv684Vmd49Q7dbPFCitAcZKxpQlxa6lECj7KwwIWA50
cByFhVskl9Jy+Qk2sKokCT0VaHTlRH+EkSGH/+8NoQRO0XCSvO40wv5eq9hg7FUUnXQRuoHKvKrh
hP8FaD9o0yItHr5Zb0A3j2wfMakaDvdOLTOUrDAVPCCw4bNRaRcJTxmss59tF/cZIzxzTy//Baay
vKyosflbW+7ee2nIdDs0X5LwLM8N0XDAM0vuc+Oi1sRytR0KQZk5q0eYRFk43V8ECtpJhN3iova6
nGUlHTeNxpJbYSzzucmSdPM0zvtjJVmJ2bsZR47YOf9Tei8ZbiGCck63Oo6ilu9L/3wIJ/buinkS
V52C/lJwdtvtA7opmTDY9GqlTbbiVuS4nPdTL/7at8ejc0gs0luU7pxXr+dcCbP8ulIb1JGWeJKy
m7fW2yiLKAMy6UC2sBp+1OR42IidnZT+ATvlO4Feinu8+ioVTVUuqekexsw42UXINTOSv7rj0ID4
cMTYoxO5Nko5WKYmkY+KZ19ZteQzp81ScmP1Aspgs7mil3P+ABaRrRDe7v4xcWo/OAxK2NE5OLyT
elvCP6SV4Bly0wcpP1/N5JDTWYfxrnxVEUUZkqlm7NH+VksIxK8E5Dv3v5cQjx46AtfRxh0Ny0Wy
p6rFp9LHX8rMDN+5SVwMml5NWgIQgLc/kB1x1D3yaQV1Axb7Tdzn1D9MC/N2VJDE9yvuSrbmneTi
X57g55dT9cEeqUw7YsdJbcIPb1+VJUS/isneuVRXiJQOS429AV9n1NUrvef+I6BG2lE1SbYmET3p
9+nSh6RX1HKPJMDb5/X6W+Yy6dxB30hZN71fePqn8dMgW25RAvcuyClPkrDcZ6iR539ixW4ZpqKS
ELu0SXhklwcgT/roDKL+f4EMJUZvl0XnFkFEBywhu3vKykNLIQbXzGCd/qMYvzMK3uNzl18Wdq8j
NhHbV+PXJOqVZhtzc/AMDJRxhAjXjX784uU30z/yle8O3RMDmhxi5bT1QMyqjUhtQfJf3Ejl1cRx
qdvv5b0Yxv0EMxY1uKgnCBmlT1EyvHUNaKXPg5kGVa7/JPWUFBjBKzS5bVmYJyzG9iAAO8XKbXds
npZaszruAyVVB/7S2imamk888dVeJrtsn8NL/4TNtws7vHmeY9qeEj1sih4AheDxSkkRU+6sl8Dj
fAMNmUQ8cv7s0yYa+eKws9KWJDrlTDDMFh1jOyCaZJlnh5zmoPOEyVz9FcG15PQu7r+AaHupg3tw
YuDHeIfOcEyXwE66yLzWgSD/jyJNC30mH4TcDGwOGnJxjqTgQ2CdSTTGRMUpuDZbOl22KogWY+FS
lOHMyTTNOvE2WJiDIMsy8JCR8o64NXz0GxjJI4Q7kLcOC2D2aKUuCykKEcwZbR92gFsr2k9wgmHV
A/ZhAETub/dBQ8ABm+0aaS8sUdAKHB3jDRTR2D9bPrTE77y3Ydjn+AHKgAV8q5fVx1bRUSo0nar8
zCI8NaiDwz0XbLjcE4ZjRUZw5pH8oQb+Onpfc6z3JPzwewUO7ZHFViBmAeXAaVAmJm/+Crdd+4jq
cXTaMsKeNfriVedxnLKuIvImQ3FlLL6eDrm8vtuuf/Y/9fuCG+c0Go5vMyS2bh3lyseQsWDrDIb4
SVnl3bmDuneYtYqs2qNGpcu6Lkez1+HmMACK+BMw0ptn4AMjwceIeRqc7zZFzl1k1RFlcu+jpwdp
y9p9ejPQFW7PA/dChA+z614nWhjboQDD3GB+6bzYP2X4NZi+tkTdkuNA1Os771QNxSah8LpzUWWd
04oVe9TyUZYtSjxjDHOH7dMQDz8Nr1KGWrZW1SogkMn6irgSFOAySGuHDc8oHY8UJcIrBuf/RiM8
BhPDhx+LSKg6DwgDG3O99kzjPvCaef+ATyhS2pHYl0ZjVVjPQt5LWea1ezMyJDbtMKM/x2J7UOR+
GactJkwgaEKmf12YiFqOn0xdjtqkxRq2FtT/thLhA9R/sTuOloQwj/hECQQbXU9i2ti1P+DQ1Pez
lLXFnLUnlctkRI6lRRg4PymIV9BsyROV8m3PVm0eDWldIcor2O1OiZW8Xg3b4crumkq38Ijz7OcN
3dqnBf6p6grFm29NgzCwSw0nfmM2wKqIqhQRouk73+atMWv4Xu7eDsaSGlSiQFNZcwZ0Bcj7Z7bz
1oT0sQY36ftfrMmRs1Po0fJbWDfVmEoxDOzuAMvfmsRroGqvdGgkM6/7xtxlBf2ucQEH6ithTvJz
ttcWTcvQlwZJ308rhr9gMm1fmeSJ59yUK0jEz/+8KmA12uln/vQCZhPQRoQXyi5UbEoj3wPYRs9t
jTKC3JWB0DO+OhPoE1d7Nh+yd2OHzvo7cSDUhsClPVb4xO8mYzEuZbPLrnTUj5+uImkx7dHqARzf
qIt1fPLe/DqPT/P59EnkSJz9/D/oRZdeG26IawKIhpM5sjsURdW1uJlYxoAU13F+kmB1Ue9BQFLU
mODJOfnsFIuusqhynpl16F0bVFFnK3T4O4gHJIb92Dt32KKehJ6QA1LSGC+ootZpCCG8M+cyDDDy
ih2taUHGjykKDsoAxvFe0ESXkr/VjwdfDgE+/S5upF5y6b8MqerRDfVHS9E5siuI6rJ41uNpvZg9
i/YU3GB47WxmI4N0ojH2fMjbOI7EACWfRZpC9tI9JAGA9YxRDLTm2WOIPZSdAGoiHstTdW+W12dm
eUjQ5N9YUT4COsfsm62zMXRWfT/lcY0rrC41zFxMKQq+xGMDdHEWzM6WvHdm2kksmNttUfddxXVN
W1QkWuZd7kN44VQRX96QbKms8UuIX67DYn/WseACy71K2sDN/STY13POlTG3q+pzARKwyXK6tBVl
Itzj27E59qfVOtBCPRurRo2F7NzkRQnmL1uS3QqmfPZ6EycAIq7zR2WLRGY5xGmNfUvfGlCht3n8
XLArh/Dk9vXvcDMchRlAxSVG9DxkfWoqXfNVAle3waRjbdilkoE4wTe/GUKrwWxi+dIKA3YMitcY
Tvl/2bRwpAAG/JCePnbMVWnTu1jCiLDzgQ9yKiZEtcSltQ2byWOLt2PYHVYHN2p3NBjU9av5gjiA
aCLzIbQrlMtF0K1pogPK2rlC39wVpb39KhZSNhKYsk9zqALrhlrFWkxa9MGv4DvxWXB3AjGwHkll
COzrB+xDCLeAhXm+HwZv+u1dbnoKI7U2KWck/1Vo58xRaNXAJovQbu/RCF4YJ973zQZu9gze7/hQ
mHYtdVA4V+E4wS4k269MXUbFEjjCTyxWpiKPcZvIOzVnoPUjr9Y9mxf3nee5CL5/rxuDIlPwrfPv
CwScLHvzgm3wWVfY9uinI+3Ouem53UPCmxt8jvTatC03bnr+98Q5Q4vmBbhizNA0OdMuyKPCrM6i
qBrIrb5Xy2DW7W2OUeF6Wjd8zJtrE9NtIGx8xvAA6guYk2FQOErPO0ZeaMrkJJgKADpN+hQbaWJk
OUFxd+tGJsKXNgCAkaXDNeDMUIEI/JZ32QkNaC50iOr8Ix/fAznjgnMvJ2amC2gqq0GzxpS37BE3
+7u+xepi6gKFVL6Xr1zTkc0Z7KgNuQ0VTZHgA66uUssu4zBu3w60qSiqelAEfdi+jX005SVbq32X
XbqsmNyxIUh+V54CjXHErrbFQ54jttpi/OfKIBNDDQ4+LLjV34uTX7ynjgmw/Db4bZo+1wWRBS17
HvQ02Mxi28WOF3aEJmXKcW5ZOq2oPdvUZa5wu9WWo/Rj4tYtn0wpjeck/S6WA4xhQir3AuyFNoL5
v19wlngbTCGRC9o6hBNeEjyu3SDDX7eZz/1DwWJaoyynez0c0ZOux7K2hbOPbywjq3164JcdXrnY
dxdsGrA7a9dzNrDzk02RHL41CHmPwx5UY86K6ge9QTAPHx1EcvY/Bj3gZ7XQJhqH49mzxeTVBUEy
xNgXKB770XmV8Np828hDcJGV96mB0N9QfYoQS7whqaMBzcvykSfUDIUXL36aM6kBg/dzCTOi5IFF
zpwGz8cBcXLHpkyIUvHBm0VdyLk1dmiWZgpAzDVkNutIHM3CYXtKBPXmtIFXO/dAbd5dmTWLzkZm
CwoZKH0C+cxLNGwhHaxW4Sc8XSNcklL81EOPnzHvOs6PcPf+HZz+4K8rG+mFeotX1pfbp5T/v5PQ
gHu5zcv32KTDGNVhMxh7EmrQdSi4PqfFWjzqnNm8SBnEZVE3nZQOAnLHsAGjiZW13f4s8w/lChRR
/vJvSSfNVAME16NJwUQ+ti9maLrFEixONXm39I3xSYWnn/CpC0TUpBCOWDq982qrqbqAILOgjRJA
THy/k4mquYxUxLBQoAgNVyPDMFyZKFK1eDT5JwlWZ2NHFUaYEZh5zs3Tn7ZTQJFgj3YrTnD6VbAI
7iU8xvprUB52ZTbGhGprZoxGZl+O7fUC31Aa4buUhVIrlWanGjvtbGAXuViiw8Xth2/Eqyz07oFz
X5FPGKTTxm5ji2/Z88QuX/ZfXXJEFwK9omSKnROqvLyx97eYA3HFHMPTxZqN++ckkUT6v68NjNWW
EHfP3iSxKsOsBozZUc3pwLChPF65LvOSrGhjoIKRyrC1stYRhoMVc88zPQlrbqAYzLFTIXJKFKzd
OhudeGZypUQMVkY2snH+FwZqD4XKdmbI/ierXUm/Bc4UVasCA6jaZHKKSTusuwbtRqacMCJKzYud
7NmJ9ASx5Qol95eSyrqS/zOTguN+AoPI/PPOkYgrGEb3N3U3oMc08V9Pj5JB1sUiMmfcdCp9Yx8e
KIQ6FP4/bXNrAagHEFCEZXeDJoOcx4WqNzPnIVWb2ZWFIyXl9mvCbuqOFXUwmsbFWToJoOY2u+YP
vQV2WqvcQ8dyiwJ8mrgig0bseEERVkvkumnVKjfAZkCGAXxvzpkTVEX6zgiCgVaEMuSzW+cZfLdA
XXLNBbBMFaTjPTBPeENRuDTWKV5aKd+ovql5OMpMsXMSSsjCxO7k1ZYA+wH6R1rDeI35VJKbpWTp
hAqd/2gJvKliORBuq8noQ7J+YMH3m+BQikp9DRW4y0HBvVWm0zSKdsgqpfnq6pLtIPWuW7NKMwnM
bVOm5FO8xJwt3c7vdrl6rR6dR/pEFf6CeBZkV3KoTH2Nd1uiJWTPFwfRKRNVXojXvzDqd4wFJAeG
72DvEvK4g0SvUH4kA31pI7R2I1asbW0hOo6Z1RlkGsQ5jLvdQwX3SiZSe+AgbTvYIhynWZKb6rxC
WDIw9xPvN5ohNQ2rmYAj6SgOEdhwcbR/Qudzd5CYTO2zdx8oxNOX8RcjZSeShDbtqhB0wAICUz2S
78RJ7s257SsUegc/WGodbXThJGelmANYdc6TcyVLqL50KqdM0KuwAqAA6zk82iesPt4ShabqvNnn
jK3/+01UW0jBybtokmltLGKeSLGyYLZNCJl4a7ZKeeRwKT9u2254gg96B4HfNyOmjdF9aR5JngLv
Wyxqb+jYxAEll6xndKJU85ZaEnfya/rwBU0FTAzmLyAncALaCwCx4zQgXP3Z9qXeqBSRJZ8YCn9c
CXyn7fRJNxje0kCv5Z3sQWpDVOX+PNpfaPy1NOdJX69wWmOp0KZsh5UFvBHX/+JTzCZMgoZSd4uu
lQfJtaLGrQ7OiRV6n+/+ZI7+eMq7sPs1aqlrIbW23NeiYyzPyvYQiYBEhuXcXnfyDe1/yZV8R1xr
oN9rcMt1wjxyECn25ZMN+x5x7clGKDhc3W/V2OjuEq5pBQc1oGw+rtfSK6UnBoI5tvKTwx9D1oIu
/wRxPcWrBS9M0Pf/BUAepaEYZ3UXuhhi59HRhpW7wZS+2KEiRtCJOXRW9RM2QYj/x9UCpfZ+NEB1
dp5UjEn1WR6yg73VMAFw1AqJxPfd019uFRabDVTzjSmeO6tj+SERIVVmHoqM9AUSMEPT6PaUpglj
IVaTq8aVZaPoEIGbvzIbO+6Y0J2iUagRW6xiJKvXcIKaYOaR7jzeeW6Ap6CXvRTnlXVC6OONzMmT
gZB9vcsbcyqdkC+IrQ+qZAxPABKRanm4e3XUyr2pSVMH19bcA1dXLuis8jEe6Vk6M3H4+QukO6F6
kubsmjfc4Cg3R3haYZSOFtZjzh4VGc0XGcZewvwEM07aSPilnYTYLaqVsec7Ir35Mvt1for3K/f1
jUitHmr6t3rWo50vpBO2Pvb4LHmhosjwBRXaBfMv4/3l1uOZoBkkc1CHkaRprltV1fU8TOITfUj7
Su6YhjSL40VTE6cLfm3kYGxJQ1Kw3O/FDYF9qhJONu53NxjYFrn5pCUcz+dOO2lBB0Emy+5SjRc+
OaolZqsZkB6EoKsZVVIrvefhF8UOQEjftbN+TvOJy9FJkxd/YRDKVWA1rkbd/4law4RhwnTY/SvP
IFRtf1VvaZ5KcA+toRI6WEhQWVLwpbVtjDSRiyIEHixDMyu4cVrBfoID1I/CuMPtNtljwYeHVATv
W8kCWiMK/CBAQUlEpTmWQ5B4NzobS8tipgaIvsPDVYsC3vZNlZzYV+fCP1jN0VcWwjco1uISVKYE
vSgLRuaXgL2bSEU8Z67npqROJYaLidALiGC/kD0RRl5hhTfyg8wWna78Rmi96huYYzjjbmof7I8A
qt+xGpsKjVfxTEumrqoee0Kw0pKTCh3i+eQ4/m/ExZVjIsiJXPTIJw9mCXQ3X2nroj4iMiNpVIAN
k9whhI1aV7sbNTbgN4zWAWknwCJVDiPZ4vMNniY+aRgagcPxduPTSVguDTa+1smB6b2cb703udrW
skitXO3kSKL5bRqPpxs2Z1ubvFnwvDlu8NO8TneDlcXg2ETIY3YugIkg65ae6EbaBNkdN8lMr1QH
6XFlD50uBy0ozvrcAsiQ3fZqSYzW3exx/op3V94gYshUQZa3NZhl7+0IxXdJNNoVE7qJwFdyAQjD
W3uCFqQXWS5LcpC4R1YNlfgjW5NI3VwMHEapFHHlY7YbbOV2oEAwQGOGDNuTE63hMeUVcLAa/rQG
lnBDAOmJsLHd+sAGvo21vM7/kJ4U0goKv+AvFWJvXEjiL3V9fUd7u6AW3mb8UMjRj9gtpPGcYifY
MrOKLo7ThfG2UDEUo2uQ4VUDtkRwFXqCoeajwEkXLMZGW5C7GShnwoDnpGF+91Ja2fnp+2zyMYgn
lNXczlhNB1V3ne7UJWiAeVEWufrxT4sjdUB5sAGHdonTLCZzEmHYWm02ymW/ZHWj4CcZkttJqU1L
9s/xcDriJr3DdZWHOelUxl9lP9QUb6m6sXdV4AHrk3mjIDNC4/zFqso3TozmIM0U/UdC0T/DkAft
oueKgN27rnbZxTaRunUnJegWrQb5DNyz0dQcp642hr60FlxvZOUAAE6y+TBnCaTXBCwJ0YAXcJSw
3FhoCmJ6YF8l4ZYITimybitW/oNRsO96jHKKsCR1tua5jOre0Dx6ASHA90u6vGwFkca/sWNDBEjs
tbCq2cj0YzHeTjGIlbCLH+weLyRkusnoEC5cI+M0E7yljHP3i1/iqa0YocG6b+FrN4N/PLzXloXU
OTqjze1uanG4JY8u3ZB7Ud/O6JHaZfidGcBujNaIJP3WGdcueo2z0+AfUtRiY7BCmzNAE7CFLmwa
4qE+HGihSLxXYSEw63bsD5UMecvclSo7AKcts3zMHUv1eNKP/bTIu97o5viRfrvHNpV1JGMmOp0V
XN14rFxmHBiaHpF0xWSI1Bvdejg0Hj308OLrJ42aGR9F82jh3BvoyPX7l4KefxdUGGHVrthjJ44s
t2nLot9H3frDEb4ctZqIb/TBr2zOj3axy0aLInjh8kvsub77zrCCqOSr1mCx2lllXQWSqugoG1nP
rJIVexTF7L3XJ5DpzSHsLNUdxBXeNkfmdHsn2WGrto/qbgB32CYoeO8Ig9WRMW+I+Y3YaXK5UgZw
X8cZs7DYIKHo1dFMU9yNNQDND+XkHlh6645+QkxGdCjLogfZ6LHPkfA6QM/NB12ZQOq4GejXfchq
+XtYYFyFR1HqcW9Mice6RL2hElr608jlm8CfXSMYumzDZ+DA4su/1/MnX5IXJYUGbRe1nleKYa/s
PL1IsOl35mv7Lup57nvBgOU2o6P3iOJOz7+zD/Tv92yMOJTczwW82IVHfSt5q4sdm6LtYCSfYWsU
M75gMq2Lxve4U9uiv5s7ogZGKDJEt2nh7oa0UAsR7phdQmesBc/DoAVrP4dDXvBm1vU3XwY/y+lx
YcbpJEbXAi02wZ6kpyxtSsmjHl1EaNtKtr4TtA6HlyDARiyoNl2hgtPw0wKK5mNz2N/pTTDOAi3K
5Od1IoCkszS8WltuhBy1RJHOt3Wwpx3NRsb9WPUvW8+4lOCjH+dkl6Pm4G70PTWAfqi3tvxi7Mjw
VsNrrSE5J3aIhAJm7aTAX2KQb+YiRFd6y36HFXD765JN41xTSFbejRdP9L95krF1+/gbivveEI1c
TQ9Zrhx/X0KC0XdOgknVA2Bk6KhZHdO7yhiWavTGfYBjAiO1Xp1YKrMneps0UVUcRY32oQjrJ6PE
WrHdkxY4mOXR4Za4ULm0pXuUV22vvb38Gurg5YfLgNrT4Coow/+pZNkXyBQAl5hT5/7kuAFmmXjX
N5DM8R6TO8za1j3z5sIUvCcvu78ROfRhvDRCumcPfcswhQ3CIWTFk6NccOQbmqz2e4i7j0QL/tRL
gMtgTrbVK+SVu0wNW+Wteruln5StDzqINRmib6ynlZBZ7eev22MYq826+AuftyOldoII6EtEqlvk
tGAcN4+ZTunNcxWxgCzUe7q0YfKXLny65uG8lg0K9NP7ZFAk5xl3cDM6kMuUbiQIeRI8/NCtjnAg
2eeaKmqqph9a6MYOOYgBCSD0igjXpdHArRLFOHiC7DyS61IuAdAWTeGHjEEq+V4u+xFEJDVtv66H
PSmiSa7vRMF42UQzVQTwv3zvcgNvoKLP/H6gU08vDwzyJGfsw5xZdZEFSWoFm3OG3z1+pUR4vMSF
b5tsDz1AkZ/MKJx6EAUGaaYjNPy1rsO1kauFYqEGPxKY+FeGJi7WKoeJGAbMiUQ1yQTiIbVPjFZx
o7gFZR2onHjBoT2W8mocYGa+EaA8WXHhyERzhOu5n3vrdxNZaMSJrRsGWKL8PZG4XMieNiMwk5EG
nLsafNexHrTma5BH676ZVSYVO4dZrUhwdI8THIXWe/qWSKvGGfRE4Wz4OxDYZPaBEyoBhAtegyEq
vwKt1+FIROI5q0Z9EOiedq7X6O1LMTu82LuMzyOCytLerwLr5lAbB1CUa7KwbZJkFfn5L3fodsWY
wkJAXEanm9ilCho1Y+HXcDsUWB17q8N1JZoSprYKKwPCC0+e2y41rM/goEV+wzjvJxM9F6sbyGVv
Dyfd+AcV+ZrpX6k3b1LwvZRnVU7totaK+G6S2SsLwDob2DIOLL0XDvIjZVKUpg8WmGqzvBbNshjV
elcvHayFXsdRL5O/1ZeZlXnyAMKY1wp7G48esAyNtPHIIkektttCWPG6YyGNMMvHqVP9Rp7tM2V5
xJAJB7Ny9q4PRw2+V2uBgkju4GyaOiFwp32/3Hxzdk17JQdx9knPw2f0m53uiIUK+tTz82doAxAG
hp6c6394ZuZZdtr06EyHHtLN0ZtLAyq+nq7+r1/M97aqWAkcRZ00630OqEQJ0Dkm34gz3jtD4iJu
KsdrEnYFhDbfI0LP4YFFVrWeC2ldXNNSZmS4GYns40+XWdVjFPwvbXM3REkinudvOC9JR7wevS1q
0D00UrGdUdIc+F/g+nlC3uqBEOtOInVQRhuO0r+Op879UGqUqnmEPmMHe5aY4YH1F42O4lMtEW6T
5UhaH6TzLAUFSe9kAiCw4oecfThneannMulzkIC1rosPVqR2GzGl2m7cQUIVTTGqJK+sMwwi31kg
vcfsM0Ej84Dtl0qX1BZJ9OCoJO1ku+NesSGXe+FXO+csNBtKMo84QN0IRPT81v91YCXXc4Dhifh/
iFxxK9pe3a89psc7tiROBCWsN5kWeKytEII+ZtUnMs4B+9IfY663spvwJW4cbLikFr6cqpkHfAIC
wr5/a3RJZXqBpAu+LlzT5VNM2aArx5khH2fAkaJcjoQm6B4b49C2q6wtdvJS+ZJ2M88/5ICQquOg
yvmD2cB74Q3/Z2daHjk2kLXgLLrf7lLS/1c7PFZRBz2K/E2PeqhzmW4O6myZMDmqVbpYtDYrEMQh
L1Axjf9zaRU2dY+FPUbCRzdwEQdnQBrcKYk2Bd+VkNmtxROqVsa51sQu+8LwCoqmJfXuivHJTypR
1hdtHrHWbexc9hJjJOKJfwA4Wp1IFfW4giRm01Uz1Cwexky3r5O9SHH5+No+rJ/WqCehIErzjGoU
+fToyi/527plCJLpVASYX1t6lMOtnVl4TnmN3wcUvLvrFVrkYccBnZZPEnu7FW8BOc9X9WlE9Wpg
N5t0NgUuVwqr3YYTFD5u0eqMlUk+kb05e/mUi0jKy0CyILmLwgRvfjMdhXhrHPN+CYfoiKIKBa13
cVNLF8YVVK+bVghpql/BLEsNNwL6xukqSLPqIR3JnCtYbKKgHyORFju16q8nSSVzyfu2VCegBKOv
mbMDP0enHATCsJXrZROrPyRsBJhFJeECcEBwS1pbYFAyojiq/GthStlpdyAf/aNwM5dI8fywXvY0
b/mqXku9dpJnWNWSykjOvvBriKTStsGl+0vaYkM4EZhuqulJyktxMlHQmOr6gRojHwrawM9qzeg9
VQx5WIOAvRx/vfjyY5WMadQ9t09bVF1wgXl42cVAHs4r+pL7UmE02w0aDZa4xVc6HfE+6S8KKo0h
WHysBeQzOVkDXNOzjo5It11lE0eRa2IjEr5LDTeBduigCTcEqmobKKz52q7pdHtR2QHQavhu1J52
0u/zU2tOP3c5INHDK8q9sr+MFaxzcQ/n8Cz72m9wB/t5abEL0kqYgHELNTYUBesEYwbeJu/l9bh/
r+IgpgndVzTQa7yA7caU5quPiCZx8uqyJnrMp0mGZGCzchLYfrs/D9K+nOXKeLndYTOyOh4gxbAy
JKvB5DaRG3Wj5BTRrGdBr8l5FDnNN/3GS1yj8AIdhVNi9IVSrS9ZII2KsHwhAxRsSHyb/3mXfYMr
KLHUQdCq9/14owxS8I+2s++ZxBy9TPQKR4k1xBxAifOll3UntJytdUtXhdQPrRqCdiCoxVslBE0R
jg9JxnityA6To+g7t4JL6sTMqTq9jmZ5QjrLEwrbyi6z6EL++iY/eML/E4yRjjbay87BnW+HHO9v
zEi71patm/3dMOFfJNaTn1McOBWI/6oXBCK8QyinZSR4D7aceUqyLwqRuvBNSUUiqjLyr76MxSUU
5vAioLfnSlnhJhSU3QHYGV+7AVbduwNBgzBGyPrP5iBeEtzxJU7qJpnBlxaSobbeAYG6iLPCpps2
o9WxRhGPb7O9g4WfsrQkP8xhLcw7DGMpG4wncajuYf0IhA466YN55KSsq1RtECdDfWXhuAijp6RI
hmEs53YK4WbrMahyJTC0GGOx9YN3//VkDjPQn/zt7VqMVaq703gytXkCLjXh6wgAYdM34TmHYtwl
X1MeUwNJz9jNVGXQhyQIEPjHcvFKD/YCegJzZIOi+mW57LGUIX8nBeB7qd/0SOD1pQKMvxEU61V+
/8+Yz1WWO0zCSjg1AvAM+CmRoyBi6KUf42eMIL8uUvFcJHZH0Ctku0tPRNmlZgmOvMtILjdv0399
j5KfGfy9QDIJXvytKRo4RA6HtqPe42iaG1wWfe2ON1mRCFFTLL7eChRsAex9tdy2fRZHyurpWOn9
dvJKd0429sHrgFRQ0OBMabBlbHMPV/cEJiAGJtdr6szqju06cBNRYBNTNIyujTmQ+eQ7NPpRotpf
hewZKU7ThmPNpo3z3E3eHjGvKmUQfFKqC22ifmUHdeh2Vj+SVuKevXwNd8W5nAD6DnbJhSvtl5w+
35QUXVxcXlrL0M7NxghbaxUG/ft58y8DIaCaPyvtiSzCyOEj89IJ6a4xpvB6N+fd93lV9Mt59woO
QYOTBV8yNT7+t359NigxIGq5dfbuQ1Lid7FqZwx8OE3xSPc3rWPkRe0Zcju0KpnLeUHxBK428p3A
I7lhrLQ2+0Yqv/EHRduUZpzFpGjHV06KcN955WEzT2QMl6rePXbwa6ByXaYmnevGFcua1wiCyr+3
v3Mp2qt6zodgXB1YQskdkwjxeDwI+afzsF8qT5yKp7MkPJmBBXiugI5bgWzslTYHRKwFKcMv5rGE
JR33jy3KLcWbdxBklYAzzgvw8UhErlwddB56Wcenqp0V6armbeqk0OQAdDY24Z1x7THLM9dm2IZy
CF81svBohq8URkrGwxEQfFb8HAky7uJGYF2s+1iQ8M/+1rC695wIh4HyjImE8GbLCzJYxLV8KMzd
FRlqIR+nUXtKhLv4uqXr0uDKTC1iUpeD1BPfo9I7e7oLigcEvLUzUdArudA7x4SDNg8DOr9Vlz5d
qQrk1pOLvJyM7ct8vdHVR2twqYuNzAyA3RI4pEVUNVyHddNuFmj6PV4hEB2ZbFyMRjKwpYJ6SyKH
N8mSweY80NNofO4AwkIZSGoBQqybUDzjqFOavqCWWk70dF6+1Qkurh51oIoTJqwuJO/Nkanwr+QJ
yNbTZFc+QeGmFfMr4CH3Beo4iQdyo7l1O3WKv5FEQ6W6FKpeNfMPKniuZL4rIjDHqKRIoHjoYq1K
cchic3paDf4tQBZVboPJUUHXYo7OKl6sW6xWeMQXATWsEUG72yP84reYA+8dTXeRPBlxePxDRwVq
Np+I/HNWtoyvBgxShyyfNJMARYtfhLX2k08LT+cdmKnJl3j0b0G1vdVfVP5+saEUI52MTQp9l8Kh
BOjy4kBC3iV6+YXGJY1ICwA+3ZyqBAa5y/FtguyTH6nbNfoa5IhJc5l90rFcaHq5ugybVd812uYF
/I00lcu8XexIWUBozncG206gXal+cJjI6ejKxrlJja2WJxGIYQDcYkONbxpaj1m+kiMrzBlsee2C
3jiU94ftstk8nO1ESHHak1H2L4m0g3cxCR4IJM049WYjccCelYfwlWEo4hsN9yOUptSXu8g0UsKT
/GnJ696xf8Fxj8M4Gc8US1pHnqi0nxWDbsCF3iToF+Il6FKJEKoRmjNzlOlvOsffDoLrIBwnJvkU
xRDrQf7ePtFfN5D7Npk53OL5tOXW7KolQNUkAoG+kzVefGwRDGUntwNN2xUlCYgFXD+VfUQBb6MO
zgVdC6dtwb4MO5EzlY71vZntXgKzkjV/vN1JOw0P0m/40HBgflCIdKIsUYYMTW8gcaseshY2/Ghw
9gImOOi45Z152FUuP2jPgqPwSNMaVJm90hVKSCgJf5JOmiMlTLF4arTCPQV+oGcZ1UtkRBM1GBPi
1bSEy1jtEw0FeVHDcUkeQpbyO8173V7wmaalE/lny/gHtzZU+6Relu3vEBXQBJO2hsv/hYjuId8z
C4ZZcZRywmexckdVSNWRELGM2oLvJJHYiSOEOuh6Bei3TMeOuApRwgHrvat1xi+98q5eQnj94b4e
5uNUF9oJ4PbqKg2GUckOpGQmoGiF9HezpfZ3Lnn9YHFtHcTkR4u2iiTCh+6up0/owDv/SdPFP28q
1mEPEMTpg5unXPERqLLgNkmXcSls5TUvaVDDE4QzxJVo2W7r0/4r/vb0egtzdB9vWcfEQeP8+s6D
OzmZUbP2x36c2Z9BSDCGV47HFOC5mrqUr9+UcpnE3cDQnMKObs2Q+MecJZ9gZQR+ZoSxXWMYEXk0
nHemHPE4yupZRh3pdhCSPBkZL7rTcFrv5t0dXRHd64UMlOHNFKf5svoMl0HztmiUYjxnKW8T+xw/
uAFzbj8tQ4EEvQ1mabPBsK7Y5LIpJur1fHOlX4PETWfQizAPJ1WJrGNw3aMA/VtiIHTxTa5Jrxdf
LJ2tWWkrGMOpPaG+7pk18I6F9jtMLZrVlmbGtl7uacQgXfdxRO/r2LGRimZZvoQluWP1SelXWzEl
Ts3Me29SKSPc7KDpjtS0mo6hrxuPRLe6S55Pqn89WAflITL022A28FrMLdt8irDNv4Fg/4FNL8/9
MyvZ7muEYS1XOfi9Mz3qdQjrtIJmYeFGOisf+PbefBPJ4Deuk0N16BsCRJMUhb4L6sDTSC3mrpOS
XBYg+h33cfeU/Hx/TZeD8i6AwvZeTpaTkxrJpTR2hSYhJy+Q3ICyDt4LwIucGzJDTBKMHbAO0rbo
FkXg+NjRIauOnV4DaMfzNjzYsAlnsM/lMne6ufzRFnH4S93vjrQQtxk4YvBjJDDVoiVCq9kdHgnm
tDisXLqrI/65PpibJOVAqwH9UpfTBVS5xrB2GGC8PFqNsevZLC0EqfI0t+GXywiAhCpCVCfbSEhe
qbLJEyiV2ckcrwryZ9/1dCoWS//9ETzklVz1RIwSGH0WJOTpel4i/zxzWPtSHpRftweYAlutnP4l
Uu8quEhYSwSJXX7amtakXrgnzXuDLcglGOfXOSEz7JsFgRp9CMwsL5W1EDj2yZU2sH4DKRzwR7eV
0TskcBpfOnooirFoOX91Xrj3NjRASbrj/7GN9sm/KM8/XF5LFLGv1zqPSmURl0HwOF7YhUMMh33J
w6gEWO135f/TydrNeHpaIdycgZyX8Ns3qNUivz0TYZ+IuF08UyA/Ac1wAJHgOmLV2zNsQAos2uAh
fpluxUmz0tyP9zkI3/J0E1hKEx8bDS/V98rAQmYZKVlmyMlkM9Po/tY9Wd4ou3xhi8a37g+IT0IT
6cMISLNTGVNrfXiNidOzhZkQBmg4mcL+gV6yehJlXkVW1TiK0X6aAu681y0lule4w5aXO04bJZ1Q
ngQslFIDKt5atSSUdoNNCjoFCYNlaG/5chXBsshK2dUaDCOEfZZWUaPVt9fqK86zytMcZhnvDQKM
uc7jZs+wkqJ+os/iUuVjewH39zSd5xC7mgpkFqtu/+4Az8JFYmTRO6iZh6rbNwiwPEG2RkyqGmHi
kaQE/r4KN9mJuYibXsNYsqwu1cmq3+QUw/ODt1dd47ViweQmnD8dymj/feQ2xkQIGpxXosPbtYvI
eL4fSuPjz2Zbx0OpmUodMAHRDzoG61xIkIx3gkWj6qVp2biv5aMBuNa17/PHYfNQsgKkTMiMZ1kc
4QfzcgITzxuvKapvFGz4VErptUwhakOLF2rLpUMfO4qWSMMsdLZXTcRo6m4K0FDh85OiJxQN5Um8
85lz/wOmwisI1KGuqvnnS/KEDl4AY03irgr4zyduKUCIyHd6dDnUfg7tKe/1alCSN0IK/twhy+TS
BwbK9ayVyC9gKkwSfJKqnQWIJVejuQEPKVthxRetzv4q+3Ez/bgBPc3V8cs+S+cDLTWBgcOIzweY
g9tissVXAlV/Jj6Q9KRQR7bjehdzZ78m4McP+CHm1a9b//Oa3A7Layf2LA5W2OirgXmhXemjVcZ1
/zn49UCYutQPSdfuSWo3L4pQ0fctp5+99Zk2jeQ3YEw2iEA+bTqibw3LVbc7/RC9XaKxs75631t2
oTS1T7Hh4U86imG+SbBWeAPOv/ieh5B0Hg8BmaNDloB/u6DI8RB1R6PMOLFRtWsGBAhT8hAj5dAC
E+GjF8O1kGSkf2JdttmxvbWF705gmpk6x83B+POKuNqlrnHQaSc2O3QWa8phVBZotYPhqhEyM1u5
kPyxr1Gaw1pZrFjsD6hGGBVX1zoacEsfteOF2krC0jhPallddz+ui3zh77A7NRZxleyu1TQG7Bgi
JcbD6CbiDC0azyptz6oNywee0KOZJu4tYsmpbDpow1IfL5Ww1h6bbDTlMMwkby8dh4K7K8TPTpTE
Fl6PpTCn+TeoakIYWWoICFBBAneihi5Jk8vQn8Pa/uGd7PYPiQ+Dt28hUsF6gVgv1U15vDcEDRgM
dwwCopt/1ecKXv4I/aBaZCA1+xXQUZx0zCNcI7P0MLhCPVBPiqxM3KDfaQLGTM0vLiZOcFLYC/9t
lfZ1VKW7hurIx0Qz/TsDNdnPF72mggM+sMsd0hEO5DpX0AmqrLVtYvMLVsjnHf5zqBuP/puobb1F
0tUL16pfFFgsj0U2j56TL3tWHM7FUwI0k6eRU4BPJS2BvZpBNyDVboD6ts2TvI1kxy3DQmLLWjfg
Qx8icyCm9PQ/zeZa4Msdjt103eZlgCXa8gvxvlMp4UZJRAH1asq35PaKSdS1uic4CCDeFfjHDObz
XlCZFi6Pq7f6BmY1xp2/tfddMO3l45yFNK+OopBclkGyKCvQ/lHRi416NAbXRyjt1W7nTdlvlYym
Q3qrsvrVoOf6q+zFW0y9VdSTaQUcx49fq8Bxxbxp+l/igKMLoh+dU10NcqE6mh4CdqPB5wOMO27H
hfKDp24lbcR4s0nxCQvi4tMrHfpvqCNIXAHG71dIGYV1hvY/O2efxmfek32V6nxIwQAsmXO90dQJ
2J2MIIloEVaNqV8rnEhfkiZJK8tsy3tQP6j03tisXrKxMuijVCOpgpkY7LBgpl+AmFgmB1M6zibm
RriMWvSYxyLe8b46k51AeX6ZAFlupFIMrF3GkVBaElYH4TMS8X12G4GeMoEPRRGovjW4tOxPh8B4
rt4wgLjhkBUX6xBK/stL8nqw90FSOtS/fqYEdy2QXTPTaqVFERz/rAEdwcI/8i99DF0o/egrslWJ
VNlbQnkVn4t4YkJbIzMR4CjwG3GmFfF4ljpPcr95BSnLWH+a+o2F0lucF/a7F+sd97xUcI7TrBX8
L5INoDP+4TQZBACCu5D7k5GL/gXoX7HaDSKQqOz31gE81AJQDg2AMOx/I4pxkN/lFp4GfYJeWWqn
D2plrpuJ1lTdB27yiVEHsXu+EZiM7LsK4ETy7Ljbiy5bCG39FUHtwOEJw7ENS8CpTChMTLSy//kc
cp0zXMnVGOP1ueleUo7DqMvEnu38clOJhHUjU4EZwKOHTv0xtpGkQJSFa8b8+GK/5pfNXa+hE5LI
I6teQoVEe3vtJyLLjPqmE7vFN8GkpXodbQ3rjpA1oT/yigTGEkyNR+FGjS4B0qn7T8nHvBoRco5M
CugCyOvHIwAA4BUVKtfRwmbbcj9p0lFdK7PiXYXhCJR1Qw6d26k/EcIxqCo9Kge2KYKx6rPtEtOu
HMh3mLR76rPCxxt+ziw8sxK2P++Af78QeEM9nVDfcbeIkD+eOiXJq2XGdqgT2qvVgYBYaIfJyISC
KiaqWpFbaiTX7IdBbA30N6+kHM/ECrvZoVGwh3sO74hJp+F0/JvLfGVKPqshkCf8r5BCB7zv9rOC
GKbjsAiWUzDdV2zhs/teq/pin3wabGUAmuDuGJjXsVEHLzUln3WlsEeBTbRtqJK0dtgwvZcukGYg
GHeKYzYUrWYNzwBG6H8j2zsUgXgNkGo7Y4feyp35pCh9k43VoSK1K1j71CS8bDUh/e2cuBR/y2lK
zvcINjvJzEx74VMiZtFOzvW6hgCuG6Eu7g/aS4wMWjHIAkpuvekxRwZ9ZJDJaw/ljS6LAKqErnN7
5j/cGfR9kL8ixTHuzXpfE4d54eTn/SIYcR35Wx5VInTNDtvuYqsqB8ENeWiW8jgy6ryg8rZkPtIk
tXoww6JXPwbAkVVUqUhTO0cCRlmoK21PU+PXtQs03n9uX6+JjbPv1XP4UHuMJdD8fA/K/gGWTzTg
MznH/vEYUZ6gZxQyqr1jh6cjeGVJJRDVopK63qqxrP3uLLP2QkZkHGGhXEOwyvl4T3AlywpY7ShF
/HnxZyQQ5mH3rSYGCXtv+X4zi/nB8AC/admwmxfScAYetpjaAnPqijA8buJFbcs6PSuw/l22s7tS
48eZz/RcOvttjZqPduVftFP4F7NsIzFGzkkCf1kSNk4I2YyMKFz0QDKQW8AuJhj6DEKV3Xb9mFk9
WC+4fVxFHAlD/4jSqoxZs/t5CqdWf9LczIlhTTS1gWM16/xokRxApIwDlDOPf4hd63RqovALpubZ
X47nVZcapRo/iIC82g8XPSllFqwwRICNsQpcq/7dkO4wQ0n0Llae4+UpLfEOnUQve4vCez0V0wes
I6V7dWiiQGnP0fksN/U2/VygcFHkLPvTyOFuVpIelf1JpoPkBbttD5/9jvRmfWbCKJ0j6TQ5ZdOu
8WwHfF+j8Wx1hFuf9dakAvawhS6+qjWlMlCVmOKReShfklUdR2vD7oPXQ23rU6Di6jPYLEx3W42P
oNeHVfhvhvxmKpoPdA3SqB1OTNPnL6iQ7SwIdUa99q4AwW24z+6HopwNoX16ItKb6bpYBSHjj3bH
y4e0+9Q+tcbJgAjizysyydsojTWOt6y6sinYW3o6gpzk5AHHSI1M8DaO6Vn00FZZyG/aT6I7Bdhe
778apujk4cHxdIbCmQE9jbKfkBK9hHDg6Th+dSi8NS1wjR5IkLCKJgGtmh3ab9us+zUrnhs8u65R
M0z9V3mLFyM/waZw5ENHWgtm6gEniZCx7bc+zTXylGDDWmcDHQxKVuExVfjZNoQGnrlnjxIIN+h0
aDcXO2UOo9oMnhBM2NJuZrG8YDsE2kQ9rlYP+iI2TDxoUOEo4PfjYXzTVrKHUpuluVRyHPamJ3xr
LZT09tdv/zeIh+y0mIOaYkxKLH9Ge21t1N3o+90A0RzZmBJJF0TKPQIlZ/h2w0nmuInZVoqh33Eg
dA6kDGnPVtJRJABK6rcW2scqDDj5flrk8fHxLroqDbp/zJ58MwYysN0GV5SjZbLnwtr8uUI+tteN
CltBE55PJ9qAocSIwKdRGUb/ijzPUJmgqPYxRDv9QrN6bOaQOjkhm85JjzMieAzsujrkRorzG27x
kaj2E00e7892eVgtsZ/zio7Pacc4EdX4irBl4F16C+FL6nhi8Xe3Z54uw/4Pq+PmpEvL3S1xT4AG
EO7ATm1Er/6j/iAiSZr9ZOsPJOq6n2wRIuVceeHpkZVDlwfK/0G6i3GbaE/wdgABHDZiz+UtO6k9
R+WKeLNxXsolHqyxoK/g9HRWIKOImpVcgRVyz82ZihEyBAy81+KknMtBKunUokaBeM0bayxqc+Pk
WGf7NXkdU846at3nDU+WMra7i5PgjiMZOAahvdalqVIOS1I/KbPlvzm7a4/JXyHqAZaxRTCzrTNX
bFier1VOCsm0SAeZ7mhasmEHKQjFlf0GhcYyitRkTvFwwdr9nIMnZDhymKxb9zOGWjABh5904bWb
zQ921XFe6EvZDIMBkMbRMzyARPoFssZGBnbWPyEzENKBVFAQDgxuhFCx1LoJ63Frl76JY2+rY/yW
5u4HbtG3NHoOjjyTTvOlyE3t9iQ3loJWhJJJX2lOzCbRkTXfTCbkvC0lC3i5pq65OrE4ucTSiWP4
d26aaNm9xOKxpeAgdzZXwhl9nBIXCjec/D6V7iTfZMUGEf37p9NFK0yKfN2dqXuAES2rTkbkH6Yy
GONbM0tJD4qL+nkV1HNQ+aqkq9SZ+yGVojGcnr9d36hdClxYhX5IsMkiZzpVuD91XGRMh87nGmis
fuopBD4SB/Ee3qA2t4kR9hXpDKzq2sDuH2btGJZj6Wan2/jhyx/vGtCJk1yolWIHSkU6JOAqqMs6
+9+VGnyIPqKdL434TqqUfSlt3HHjQxUgA4r+22ztA1O/dEKdx6fo9PdVWCSo55B6AXD65pkdJFXt
hWzb/8GuO95jbtHXtreBdejj1GboGZHtxgsoJonR2a6F6yrai5849aw/wqhRokRKFZZUVa7dMpmn
pV6HVtn3Ft1qUBmlgSdsKOvzKUIRhYSBTBsMpRHM+bInRpe6lnSE1hSEOKGJzxbHsmKKZTtSyC8W
SqK1p23MPdOVtcnU8HaC0kwAf4e4mFEXyh4CVRPPQeEQmWVbWC4H7TIuXgHHC4E+9KK+fj4Xgytn
y8eWgmYi2ZSjUY4Fj6X3kAWkAFDSdb19GFELAHk11TmzHMx/etxTZvpsZMj09Vavnnom1Z+rSlgp
1RL1pVVTMIy/Wa4qcl1utI7SkwYlqOyqYq9N5QNUNNgGueoLwJIp1+2GssuV+ZmsaR+bNpo4Sxxo
iYDvq81C3kxd4j4VmGTspOPR/k4/7AKc0VidKDHc8jUdSOpbc1ArW1XvEZKBQ5ClVAC607kdHZy6
5AVSR7I+o5j5h9YBJc8WtijR0mKyIolU2m0qiM+HkAODfq5Uzs1BTRnYt/sBXAB/1pymZwdJh05F
pl2K27Obq6JZ/YSJ7h2OeB3H5T7VF8SdrQ1TCnNKwGhBMBig/i9jFLENhsxkiHOsVxTR0Nj5hXlh
lGhNsyXddCf8HTx3NvYd46aAsxj+LXjZSyjXHz6fCvAeDL0+qG9VK/m8JtWyc9p7iZ+yn/eSmVgt
k+O8e9tpAv57UbRLYzGK4nQi1fSVuVAiojpO5M8fH36VP0XHD3U0JGvWJw/ITOPVk9JgAvgfXFhE
2FVaYBHQmH8DLgials8yb5MSolrCSyrBUd6CsfVvZxAPndiu70TwpBbGp/41UgIkpNc4Lz1aajwJ
rumb35V+tUKJJwaUFFD/IsolRQ5zc6J8MQLqK135p/eMHI7ZSJbGOJ4r3R8wPl4Iarm0G2pbd6Mt
DqIQUZyuELNe0jXvNiExtf3RgFEpX+gTltr4gkEGgBpP5e683FiHd6FHxBCysClTz2sehXuVvUTI
4q4zTlGfHXCMssaOKQvln63riwNGR1LlMebaP2rR7+Mx9jQ0pE4UWDm+EzY8w+AsWQvkv5EURW0T
Td5psCQPNkdYY8CPa3K+ubeB4BeSi9Gby+LY9iHdCy9v8pf+Mu0YetmxNE8KV/+AmDdmQ1gRWB83
Yc7QoTYMlmMglUwu7dN8JkIx/PQEfwiGJaZojob/AQnVDP+8uGK8VveltiNuSDsxHAV2pK8QU2a8
ELazonE2BMWTa/+ei5FR716XoeUU/m7bikrv1g0Z8G1nVxhVflFwqwF9ncSsx5UMluqAK8ZwFOf4
Ve07fD4NcrAgIOn5ywC8JJDmHtE1GNBeaLrm4mWsm9rbtqLkGJSApFarCCEgTX6/upqTx8G45bhw
4ZruinOwWmHhx8UhHHDrG7yL1h8IQTaJqIHnn31R5VviPMmfLlsP4J91FNaKB8EIt8ZNnOGeEmdE
yFkyo0IZtDmJvK9e52ECl5OYZTijQY05oOECFD4oD0Zdjay3l3Z+lJdalzxcNpGpxYM0+tc2qliD
iNI/mahNf+aO5g3Zubb/8EvSCiwj5qmuvH7AMc8CGM49+pZNGyV33aoRUS1zjSc0YMmTRYan3KP9
+qJ68pnb5eE8sjH4scQ1BEHKzxNc123IkiK14uu2s87VvY26I2ozMGclOwsVr8TaQEFGVLC7FCKY
7CduCnYV84FVo8vkf0gaWCgt9b29C6XCvK12FotS2Cc2bj+F5HU0wu2fZNlRP8U4F34gvm5OMwxM
N/XwItBjDgK6666Kbdx1Hy329cy8X5OtH/TrPKBsHcRJnFYdBgYGa5rX9FHX3wtTgIoHqppK+fnk
QqrxD9h6TKBSLaIqets2aIfJ6mGZOqOU4iNg6qdnjPE2SiEdRPqb+42ie9l2fdjOnh2QdYG5bqhl
9pZKLqliIeTMujnrwN+lovlT33pIZVUkNYKNG8+FvcXAToCPyl2VgoBTubQa6D8GHa5OLddex7Ac
lV7LZ8EsfMsXeMAXytbGZiAnFHrzaVwCbpL2KgILxfFKSOQe8hE1+O9QcYE2IQlxYz2HdjzrKSyf
D6XjXjwsQDv+mwgEWCwgzWrf/v2TbFyYCQpnBEkmuBfIjRGLFoZOgL0lQrYb+HsARwy8ceg/iseM
+HHnP9Bn74wBz4XjVuAzemLFYfjou5oKjMJO+6FJgYYygjMlrViO+jq7VdEHPTl0ST2jADAhVAMS
MZ0bbd2Ez7ksWzDy4pJHp7u0DpiwRQS3GxIK3VEb51Yi3QlIvi+/ePMs4jqx4OyguCkBWFZd6E+b
RtHvBQCGXB7emYg6BsxjBEyAnszDOCfZ5CLkc8nLCn9lfVta6uCB0SM0KXXmgC+aGoi3sGPUolF4
7AA+xaA9+V6dPGii1uLuKq7sq+9ghxydtXhkRGoO6xSm/jaww7IKMQwvE9jO1A8mkaCOHvqDLxKT
0ZCqvRpHkuMhlVZV3VU9rPTKzdcxbl4rPynlKtQXy0zsot/isq3kV/rEJftOqLMZ7FA7ERF66qo4
LNMZsKyP52Oywhmn6GOqodebarxxYGsFop+rPK9nbWXSaKMm3HZ+pE0t19o0Iv1ZD3cOd73D5L7b
o/S5gWBQT2Kd0HwXOtrmbex7OTrzB3/ugjDKzoQDga3DmLGr6QZRABRSaJIoiKDL5U298MLSWYZW
oxtM3xBiXqZAPGijNqbVAgeLxezK1yfu6MgRicGbgCtupXpCy3DgIi/QYAggfGff7AfMlPTDgmKc
NCfUZoWr1jrX94fK6lVEq3Lr65s8ZIc9VIdKYFOw7SgEcz10xGd74hfik3N6P+x8SlZto9Cs151z
UKvg/NXbqQD32jBo/+32hj7UOLX0K5j8NDqK5jfnqEVEFKnuo0AY38tjO2GpY+2PggTre15DTZC0
fUz58xTb1J/9YnFMDllEnYpf7zGEey1Fe6pxiEfzDjrOMFCpRVUHp6/iGcQaOgSMbc1VtiVf2qqg
G5JlsQP8G/8GHHtkMU1R77jORjCTQavMRxgqigpyJ8ygulogf8sdlF0KlJ1JaFrjFN0BZBQjv+XW
hzNhj/WTUdKGp0t+czd1c5vUqoSjQGBjLq0HFOMPnb1Q1ekAhmKa6oljfZvTrXY3JXkyINAUNkuY
UkbxwDeDAqx6TQC1afdI6Wu3o/OEaZ0VC6+VVWJqhNbkve5cty1rTdNUMMdcicD/8WzsCsG0eNtq
KQ6KbYuI75eyMJFc+oX0i8A3FhRX/mX/EaMIrC8BDGKgB97jIDY1YG2GhDZMlnos3g1pMDeyf5DI
zREOshty9F+r4pp6ygZSGOsHBqOV47d4br2rHilCyqHoRi0qXu8Ej5xXQ4fUvyGooLmJuwzjxA/R
AAQwCciAwC4nnrRqoG9A65eERT2/vrnXb6s3MGT/1Hso5r/aQIsd7CZS0bq2R4LEvJrQB1wTRkq4
lKcVhunZHWCaQUvATOd+TE4dfhweK6+a+7zldJecegxHuagGtdYNDpcBARGrurSMwR6QVGYf+bgi
aeYvIoDjY2DIjxDchi6cpKp0Kbr85lO73EoA/wHxk3zN05vRinDLTLNunw9gM0r5CZQCS6t4JPtQ
MbZUU3VeHwKV4OMrzCwjOL8DumK1flFy6NqiRe++8HoqRjukLhNl7OGi1b+qsKwPtT8GmL4r3DES
I3fGx0cLISLFLNPNIUVfFNYgxtpzdwtk0xW5vpZPN0lfLKAkesLVDAN/OG6a8z/l4xz6HQ4eu5Qj
h3jKajw5i0R9wN3X2WFYNgKqMoimaX0+or0LULrXYwwzcdaD8JI2S04Qh8qsNKfF0MCCHJ5zNp0M
q273fFon69PJupYGYPvm75gJRfW3Vbbix30xsY+OJdxfN6Y+EDOswYFDN7vuYzXOKcKf9k9oU394
ttsbxu/4oyvymT+vKvrzyKs0KucRITcSc/C5O74DEHwQeFjZgT3tLkyKR9rQLVYOIAnpl2q+oewr
feSDwdo2wNDxj97hHNB9pX5ulQQ9RpNyhhdEPTYctWcdm72Aa8TcJjsgRzRA2raHid1C6WWIbTxJ
6N1Xy2Thc7iR/Zge6yhtD3Fq8scuLpFIWFLzr88+6VshPpmoteGmCbDS6DzpBC4Qf2TldX+32M1R
oCsJv5Pr5HNECn6F2qzoy5Recn48K5yvBs/ery22ecV5aWV+8a9j43dU62ky0HFcun5YfKwGVaYJ
0vuJvtdyC5eSyQbloIyfA9vED72JaeDEJJmwL0MmHt5GIdtcCJW8QTLVSYqkPWQE2vsh2bRtmFTS
YETvMT9Sl3tMDt++GyJ9KKNZI70C3vO1cWt89FA7kyxPzJ4NqjL5wHNGQ//KQO3ZYUJEZRCJOBeV
CZey7TAtwjIyq3sHH7tonZ08ilmz6LChYgK9r2cVoLlQX8g4RmjwQBKDRGV6148kaveOTVSrtmJO
9ZPZEQnq4OU6UvEwNqDUlmLucvNIS17Qxw0nJeBpjPG0Phkg783LDVI23M4Hb0xhMvO/Bvf3o9u6
eAPi7XidGSvWFaNGs+gfyd4yP1lLkbSTkthR8LKrN2qUJxAXEKi8PYtatz1TCgELE4D/88D8B9Wg
fwlAFB2bzXnOkokc7aU+QCs1qfFf8ff65qH1no+acE0V+3xOdvUPgwFDSa87oxGHfYna5b8FJ0LJ
/HKa8XQCFH9jSkRwXg3aSM1AbARbaKLNjNMwDsd7ErggTyTHn+gdAY3Xdg+UZNt73hFaqkeoi97J
IbqZuJ9uAaZvLB4lFzQW66f466g5Gafj9RrwTzDWt3TRxle6p7sM4NMNZM4BMIVXk6ajonV4/UAa
YsBkJWHWjuEb38Ci53MwMW4CcWKzy+QXfZjNz/wkIt7Y1AGyxUHVC+w9q+/aVPhwTg9SGa99kA5Z
IpDtBXeQjJSPFFOtqIDxt8e7jF3lCe+12BQkOLJnxs9vLxNEmaCUmsNbx8GhTcwKXC20tpd5CiIZ
l1+Y6h3tYGL5GaAkwRcEHgGCo9bQiFNly8mw08d2I/Rk7JNzrj1+HTTVlOwJPA9C/QL8mlgVAc/R
V3E+nDO8osmNndIhr1JuiG8CdPrXTZzt+94xowhWXjGqUi9vUQAsPQYgWBs8aaPQHG8DQQM0KB53
6fHxxtHQc8YumSUUez+yYxYEFan0SEjeYakaVLqigqbkAAyvFSa2zMOC85x+npU1ru2dqy5SCg+2
/yB570iPjWUsAALwrQYZb7pyReaKo98K9649vDgtV1yl7KBUtfULlJVs5+DIHSLuB16xN5WtSW1b
bCfRMczyiPtId6EgIMjuDjqmiycU3yTPdgp/bsrbVxYcroJBiJ47mk5F0GpT8M9NqoXD95m+uu0r
gNq4xQ0P/1GF8AMADtfjBmQAPUZpGwq/apmerRFblOmeloCJvEnaQnkUjRU9+tjOCNPSQDLHiNDZ
r/hlXA8Irp5VRaziyw12SPJij33+kL4zjqLmsXEDNTsM8aIReOI92t6x57XNoBhwiLNAhki6k8Af
XaPpo1ZYTUGY0QUhGCxvVYn/OxjfocnlvLosy+GHmcnNY+ryULHpD7a1K49E6FHwU0l+TkymZoeu
kDeqdzbvM0fwX76Zu+o0mFKFiTOotLnOt6hMe48AlJW2rUnUhLI2TEjGmnBJQpEkv5cHe9Q0acx+
noKaR5vgQLJMmxDD8wWaUngSTNkX8w3YH0aFD0UzbdZJ33YRsEvUdyx+qc96zn+ieRrYqK8b0vOY
RuWVo0VthQQG2W97c4xwLlaRyzdzfqGMOEaLSZIaJL0/7VbfmrlZDIoiKhuZIM5lleJlb0LxOdx3
/gSlQxKTC71UPNVJfBDdxlez2AIvhmsqeYxXRZQVcWnVUUexA3tU5n4J0zxZN+70slv4Q0FKtmdw
Mb1pxmlTuekiQD08XxS7Ktlf0/vKBgeKwqk8/m9PbIj5yk4T0N4N5hNUeTQ4z4eLeP+Di9hu5PSD
UwS8dV4e4dUb/YvRjxC7uhCo9x3w7QQ0Q/hSkAf7S8A8PV1aozYJCEExfHou50UWiD49N+qRYoRj
+OO+23XWb8I5SV9CgIHIML01vl4pCLz2LG4z5pG4kCOqkWjINb9eK04AbhCHzUAiNlTkTuMlRWLH
jD+HFJ0zKuULJLB4lzYx1O64vB5dCoUkmJieqdD5VVspz4Tja3FGL4NlFDE0gGk49D3FfNmJiiTK
2G81k7OcftKW3mPa2O64aEriWdSbXS10FgCOedHfEw34O5nVUExSxo9ec39m5tTNLWWHPl4erU77
1OfwzXF5EJcSHiw1QiIAnExTNOmlyX1JAJGETHz6/BF3FyMpdi+5ZIIyYXzEWV6MOtJrkIIr8VeF
i3NRDCb1P3KD544xZGsPzOd5rS5pxFrn54hhN/IFDyKCLTWI0dpTvJvMG6Bm4Trg+U4faW1yZj4D
3c8OePzZd2wimtRPjVZaGm+LzlJlLPIw2YRPgSFja4Tm+cPoNa4ND+H43JA9sEtL+/Q79L70Nm28
ZkgO3AzQwxDhEKxjYwcxLqsCnChlDo4GNikRt1pr+XD0AkVtQvfpidT/FRP1+4FfOrpvbTGr1Jgy
qh2UU+K+gYIRncrFM6EtLrZR0er7gHdNHPnhW6rCVlkgI4QVc/nO0KSU8U2rU2b1YWI2J3DvEFTe
gKtpC/4j77usTLTU1XIl1X5l7il/5n4w2ker4sRZv7WhUjnXMYcZLRmGPdavPNAw1mdePGbTtvV6
m3MyyBx9z1l6l/pMTq5oZo7o7tShpRUgVQCO62WX1wrWmT/V3Pxg0mrEsGWwJ616DQuf6v/QoTYe
zxIsAvq5q5ihW4hAQxfLkj1DoRAVkBG4txam9IzqzTYjOicRvycWbONsMTn4au0CmVG68INwmOqt
TvEOpKJj3Cv6VY8KMvkveN278bKm0EP+CR6rnYyMDjR7xLazMJQIh0N9dNTYFs+2jr5tCEBXBlnw
F9ZamKfQyK7FkSHWJGP2OuMMxajTGMgt9cyuZZkPCogDeir2B3/gQFgHVRLi3Q1NXRtyW7CKW7rT
XBYBf9Cvjwlsk46QAu7gOUiRu8JHoRVYwDPgRWHgngjxBei6clcha5gnj4OTxFLwxvwSEXYZjRl0
ts6I/3Xal2vKJSZvKWVe/Luio2lgHk9NygYSdYPXPL8vT5lThcZJ574zSHIFNt8NAVMUXvw9cwSD
ePnCg3juQIHTAwAEbZzl1LUGSRVZ0m5hqFBlB1vMZudCt/e7qh2MMOFeTOXprJJWZoO5YqoB+SZi
YUsg1Oy3YVwc4fUWJu5fI8LwP32lGhca1qYHs+t/GkcKBXQVgsV83WPH2DK1bFG3HI2xBUcVUlkq
jMAfSVWPAoK5cDz3ax37zlRWC+RFDzldFpePUDWO0bzQHUgkH470bYYld1S2fX3rPuq4lsGL7bfS
p/+SuucqgcJA1I5B09YRzsO5zTetGcy8ck20NqxV/AdeKMYOeRbt5l+Hppl8QTqiWG3kri30Dtke
BdsUxOtqXSu68Z7UdadJosUmXNiS46fdnAc6Z2Wvu0TVrZA6zLkfaJm1YCzNwjZqXNx6QQwVKo0E
wAsKl5P427wGUw6NQloyBc3kpQ2cLQk3fw9vbd43MO76Sce4vulxbUZQhs/MPBb99GYzF5aVyL/q
SOOZWsCsSb3LWyxd/fvvKOpj6Uh7uoZzeBNBmuQxYfyD4FZ+Z09wKQ4maHi61nB0Y4XPmpELi69c
PqGpSXpbFGIjRsPLbZdIPBaMAW0Z5nojP9+eZ0ya7SfdJwiUtzyVIi8xvG6HV/Twtpbh5f0nP2ZU
KokODtTTQAOolVR7mZbARLLTJU/nD4FE2TILEkc7NGiJrv9ZcLZoo7zf7mrIQm6Attl+Cz2PHtkP
3xTafn/bMdfnYCsbMSWA8KkXcWk5fuWnJcwSbVqQk0kLJzqMWef/jB/lRAO7AaiwxsM/uA7uZWH4
7W7ahNPO7Y/omHIlYhtOY0VETVmhhbS9WG/u/ViHYquTmdlugIdyVhV+iHPSFLLUZp9AOKP3c34K
Q8dV1Std9p/u3sL8q9QKOH27zeC9NkCQovqLUNh3cIul6YS57KAdJTa/DV9SlH1lEWyKkfvCQ4nA
lUbJ6bLOS+ehDfSgoyHlGtawvqXFgwADTPBpjjj5ec758x4rT4cl/eCFJ9byz+oi+BLPo3pHICxQ
MnAGv/DUDK/TPfxg25KY2yH1XM8pQtoJzTwo5klmlAuQx1Sm2QWkwJRRCw+U3WjP6v542D2eCFjH
U157e5K7StJDs3GERtmvAiy5vbOm/On41n0gdJMTyZEa4xbdqPboE1eYsJgvOnFT6W/mkBzIZnjd
49fSEAF5RLHxP0IX76i/w4pqME4IDBMEyFciKdmeahQ9rGLdHpUgFXuM3kuSJywEzmxniMvaC3lr
0LsWnRDepHAF3df7iiU+6BmE3wim5IrY9tLOJAn0R8ot+P5EmJUlCm8Qltz/hylR4bOruRbxybKd
qiYO/zcPlHq4eNzNgcQ/1tS9lL41BxG7oZG5O2NBZWvcWxSMwWaaYT8Ji2qqi0pEgZspXufc6zAI
XSBbe2V/suwLG2APCBibuG6sutV81xtHwuSqAlc3DsXhhaf0FBgTX81JDd8LRKF/JxV/G4Kx7ZJz
i4XYas15wV+nagNzW0DprBlRID1SsN8TChYWI0UiW6ymVH6ejhb8tiuwqSghwQtxhkiT3VRv3nkw
9RLMLtWUKXQX8IfnTzXUb87A6PGWTEQurOWvZgZzvSOZ0Fn1LzXe7xYL51wX0JHn6a9BHUCLFEII
yaqdh3PgLNlk9rl6z0CLOXs9fxRyKVUOKOIY/okGQDcYISUkgT7w1BVYdDM5ltgZwC7EQ1+wKgq/
axwlqBSxVL/x8GCibNCkjDykR6bj2VPvL+M9XJpL5dksNCe0yEWfjTLW2fH1zzjR83VMZcCBU9gC
7pqC4A3H1XyLyXr4qVgW1f2CHX1nd+nGswSfyCXWVCjbKV9zbVXPzHqL0U/b1kOFICM3D9pzWXsD
M/nEYbS/QzXyVxwP1mooJk6iAv37MXH15NnM7IBeHvnvB0IHw51ITnLqg432Qde3yGY1QrJ4d7++
iOLLHDvLH0SsutZdebTAt3QPcNCmgb45kQ72WXdtok6VmA0L71mX51CMwplFgb+pItszGofuyv47
LOErTakgvm0iFlbrBUVIUEcB/Iqg2XTrfkX7SaUSsMtPUmwmn3t8HRmocPC0jWTIw4RuRkkCCyXb
B1xRl22nsZYWrEUr6DCqeDw9xbnr6d28kEVfcIAAAti/zQS8yZDJM7h8iQnVg9a7C6aI+byWqqTj
6pTZOIf2OGj6zma4PnObyzgI92JE1fkpgD93wJvXrR7uB0elarcANUHmSDpoaU48UVGcNOYaoHGj
qSoAopI7hyNHSw4lsoA99J+6ixS8C0TGL8iRAwQytP4YbQ5hn6/fItrnQLw+YWtGTcLyb0d5w1lM
fAbANmLw8aK/ZQvmqQVEoAspr9QQ6jH4UUZvfeJi0x8nPzh//o2H/JMjvdVTP+OjlSD+l1UF2Ll0
apPTSvhqlv5XdITFG90UHG61JMKT+hyq7A+X4mDLzYnwp+lHpBJHcyxhogTKWdWgjh1VPEbNDgLK
ozyPjkJzdWPcXeyKbu1rMzS7Lo8CYJElEYsbmhOROfKoyaVOjNEB6KtG64yW+cqQwSZLX7TU0iwE
mrAkU7KpjfxJKbaGbREXsfan3Eq/JsQ7fMbYrsF4emzZacBcMzZlgBZw4RuLnCHl0A9N2lkQieku
0+JDwsT58SsfD0UEFxhyJTq51iI62b8L4mtNXiVyxJmhEszga3rqvN1vKqVbPUTzpZNzQ1GH/tuH
n/ltoIaXbdqjAJ0+1XBqnoU5l3DjabRVIZRFyBkJ8KX+3rlpdDWqYgP9gUQeDV4sW8c6is/wsMwM
qS6fEQsIXclvZWQtTSMLGhrDrrQWNcFEBaRak1bVV/wzgsajEwYkv+L8LcFSxJjRX5/RgFpjgzJ8
+4OD7e+1mCoIonLxTWr2VvDhb0NCfsI0g5h7mdWIyPOZZx02BW6/utEmOFNWw9/a2adOEy+tCDMT
b8kE6xeIaZi8aVWUxkg6qo9FMulC66U0LME5lvzA7ykCWxScPMga3ff/p7V+PMbJP4QJG2v3zxAT
DMt7fiQkv39vf4qJVNoUOJw2EaQmsJ5hwykT2tJOa1ljvna6MkExo+7IbR4ytafUC0KYPVp4Ko3h
nQIY/DG5WAoJuKtPrbh2pQDoRMJq5Jk/0Ag2S3o23jspf/5rGkc78lr7VF2vHgX7FgqS15SuE/+P
hog1YKIX8yC+0dLBQBz0oSoNYIofIiYC+eJM/ettptfPvtUngP7ViCVuukbG7umRbayTDRg7B/vL
4jgqicSr/Ig5SvjkHc3E0eaAOpM+40/wDViOu8Z8Q6ZkL3IYLukSNM5PVp5w+7f15pUpLrK1NuXb
0ysvs+YaUdXCCWIe/3Cio6jc92Eb2KhXvrPgA6Kjiba+S/D48ZHi8V8QMhR3G9Ym647HwJTSWbLq
xZUt4KzzjyFv4v8Gxc9rNvMH7IQfpD+gBNqJJcLVBBoj+6FeickAKhnH9J9hbhdaE2zIBeFhxker
ZgW4RB6Vp0jf188JFn0BRJu5D4iefkL2hqTOq1JALS4ujoZHfJjo/7275WlJCnBw7YCGNEX99rTl
V0fOZn8oxKCsPSHxdriJhdZccNom6EnAaKv1/+th9jpQxJNH0Y5VOY5mNLM1X5tA7qoMtTwkvU5Q
Rhq5xqU18tKuvq+jXLvYL7iSouT/V/EhSvESegUJExfHbyhdX1o+4svB0CYbjfnsX/spAwhzXICI
/VefmAW19+T4/PlYA4auN4Bbw9ebj2UewK3xRKmbBmQRNsexWjaeo7namd+/otdDQuJcHNqAhlgF
50y0UtufuXlvT8LlQfdceiEF9mzB9rK4CEFzZ1kGpOI/XMQQAZmsqu5CtRKLt/fXDBVq8YrSVhsr
DUXm/NsCb3Kxr1/B5dI9B+br9P1OA4yMD1OA+/+/voplg1ng7Bz5+fqLmTn8bJyDZ+/AgsDD06Rr
mqi2iw1z+/MNR1TTCZLeb3165Nrz9uSe9n29nLTdVSbdmGDLnr+Wbe20IioZzknoSPJagApv7MW5
Z6Bjvz0MwN/YdT8ClQN/wfTkoXUkaI+kH4HUIVYts320WJU8X+4StCHm5Ec3B+Z4iny63V654DVe
UYauFeCpPaGgBe0CM9ssK5zPYdGLTpr4chmYqRWDk9UmVdVEPBouzk75qeElT7cZoOSofF5t2Rbi
uZFK8/UIxsIJUHe9J9bRoWn2Q3GazlbiqIB9SlacDqpW/dS1ChnAdwI0CF/2Y2XKsoA9mRxb6MmI
be5MTzu0Wqb+AXXxHz/pCx70hRNd64UnbuIZzFPSgm6f55pRD/W+kdYoH7SNuHSshEERwFZ6f7B+
Nd1ARgUR+ILcj7+CsAlI1SA+MbhKJC1kLOXXO4atxcPXDaQOdrJSynCjz++JmHdFMXTomZYA8kVk
6kb1WMACUnNVDFVUccM/LXpCiGeweVrgfCBWJKj9iIcMmNAgJBEpGu5ahTKQpM4QEkzfNOtu/I5a
poh2QTx65F9Rs1tJO5noo3lIRCm7YX/MsjB7b36lL2PU6edP8C224g+pF2lNFlJqZhtir0CSguyW
E5IsMS4AOj2nY5YPHUPrdPPFyCLVClAylMm7RjWvUfgQliWjYNyocCBJlUEfN1zq6UPd3+Ps23tz
L58nmWaBcRINAgAB+2xz4YuDnmz4yIMdCnqM2YKTyzW7Wpl/dVflLUQt+5WjFqWtqgZSIoCZMrhh
yK1bY2DjCaBGmkGFpcorIR6zJZU0+kN8w/dblpd7YURvZGgz852pHR4Y+Ek3SqWeguHpX6I5vweq
tfdScG+Zjj2BFyRNU1WI3T6ay36WVWVjezxdhINeCcXZaxLN7VLt6MvI4H8E1HdNOilO6c6WJkWH
3ZmoxuGELhBb/qWj3+DQ1qiADpBho2iUUGahO8koMdLTdqDfrQtRK9TeEzKuZ1y5vOjVQgI3UJU4
0kO07LL5OsDfTMpUQL7iLbno3lKdrib00ffvs4DRzqO5OBwPaWVZlzCl7zZKC2OMJ/mD359pVfQq
pr2ubVDVLmsGR1kPfLvepqyRKt+ai7eUiCGAyy0oAcmqAMxxZXPHoJPCVLqIr6grEIMOsnHCmrGS
fOA1lNavjcbegbbsEoT6IJJT/U+yrfJJ9Qh3NY6JqRR39dja4WQDH52erKxYQjlGRRLo9O/3aalc
YbLW0qQeo+Mz8vY+eQd7oJiO+b9f9olr4f0AhcKAlWwXFLL6wGIomk49fsKhzW3EQ8/EG29PK6fA
747HM7VVSiX3Hg9TKaKk3W3M+4urKqIDKWzCU6XNGeiSFON5W7G/aifAfyowHoQXq/y9WapJBy1a
FbzuuBOCdEe/gHczOX/zUV2cgg4tCBJXDiFlsQK1GDzwFjkEp/N+OW6rZGtbECWUzMLJCrzshYBF
U1gxpNHrCQ2P7OGy49R1tRpAOY8nctWjF9FgDYV+Gsz+ycGYoZmpnwy/0e7/BWmFDx8RJs2JAYZ1
hCWfBRNRZx121sUcLNkPP37kL8KM46WB7DS51TBj3MmH9ZKFoMS3bczwen+kttBrweLgZTOIvQ/T
ohnrv0jIPqGc018UxLiDfLvoAjcPvkWgn3POEpNtTHT6Jw7NcgD7VhPqPdGgbLFS5IoNzojI7rpv
oWtWs6rUDaMKIPjDDkx7vcII/p23KxWLpQIMDRgNKdZ+isN+GMw3VcihfJkEM5SiP1qTlkZgckkR
3mQPl/WaCqarMJj/Dlgza2HceqilNxzqdyoBaeyI3HgvD0EKgq7QbQr8KDq1ShGAQOu8Kz2DZeLn
aL1sqGIAC3/dJmLWMVvhp6KCQ4MYX9xEjSOafOS11kzEx+8tt1WXciALI1/sUerzP+62XxbjCrGO
ext7Q6HKJPlnl9WhApsAYHTWktkVp6SVOa/RJZt3QWZg7bgAfKnUFj0NV6wKc0KyA9zMvm3OUY7J
NDPLwrQtRyfwY+dOMn4IftaDhKK8tIzMxnUJDUE7nu6/qppU1LMTNcb2hdmnQ+15zGfQBaZF4gTf
S3dkwvV6/GK4N3oPgM8HA2yJ9wADbnhHxJD/TWpwu2zO5rukGupJmXPFbeVMPMrNjRTZ2iZxjnoJ
ZeFwp5CfUkRn55To0Rs2iTrk/07sRmUfhJIhAH3OEJy5ko9EitF6IP/qI0xlfNV/Md+fet+rW31q
CFv58u/e37lp1RQ3UiAe9oNoPdX9BltO3mHY0k/f5foHPTbsxvvzPnO3yEaz2L+Sd1LswjDWaJZQ
FSS3ij8lIYCUUdymy14skschP3uOxlHJqXL9cjBsQijLdYxhVtMAxrI5aZISgxJZ721LMshViK5u
yl5MEjSwrcXwK214d/TMxNUakDnZD9DQycItWGGAl1/7Akf1bAzxxvkS4dDdMsLdxoSVVeR4gAuP
ZfxVFh/4UZQCOaJr26WN55TNTqk3JYcKdyrCkfgev0OfJby1oK3wQWNjBaoooFzkuA5/XRuuw6jd
Os1G0mynAa19h79q40fSWjr7ADH4mCUu2EW2yc4q4wrlL0XOP1vq15GlanyZcKvBvndljkJbEyd4
si0+dnyZcYeGrTZeTgEqnH8oLovnvld5NxHxNtolL/AzXG+nVrZFmJ/rOn4FTmLZDifMjONPnCFO
nBh7dEHeywWVL8eg3tThXMguYT1xxZ8nzdwc/qpI9m9WVop9TvJYFWG2oPhgIcjW+q1CsA3jRnsz
80b9R8jCNtJMED4j4j19x/BVWK9DeutF8vBe2fugBDKaMZhdOX2tpyKVmOVOsII1zN1DOHSk+GIN
b9pjgp7FCZ1J3Ru7VsoABoaigRGC7s7W0pTTczSOTnGqpkC4tCfNNhJieSOAZ5sigqOEQJDaAHeo
96UVArLrfTQmP7ta+0cXgJdlmWweB5+ojlwoZ9Hu9hI7b4v5GbNkNZ2EIVhPnTKJSVGldg5qbBFC
6mVZlhuz/ciIpjW1oB7rOpfZx6LXcV7x0xBjrNvD6yTv0pc2fEzLZqqoIi1+z+/zJzFe+7I3Wa1A
wGx0lz56+0bm53a18ID2n050VsPACjRm7ZvAetv5THLu7TrVEp6qIBOHhT3LQrjlbNroteKeTRoE
P3Zf6AvJtyhDIHHRkx8WqGw10die5fhRHcF6EnEz0CBYPTvuP+evpT1vgJlVH1qGTE+B3DlNvH9/
1bNoWpveh9QiVFT96F9Zw6/LISh/JW264wH7FarG3sK2RB/osbivjHTm+PK052l72xJ4mLc0HoLP
Dq8pkrdLIivIj2oBg4iKNIPRKyHbVdINwGR1/8o/4K0yufwzQM1LO79OSdIWMDBqzb7VhEY1OWZ4
GmAw7IUaGWyYIGL0vlwhDJpGpwWBnnKy8R6T/2w9HKmOm5qV38J+VrOQxcatbTEG/sNtcYGlcOG5
ixZxLqJyWsKXBbkxh2iCEz12nowjDwo3IcslpqQ3kuth7YagCgy7766hI4oxCINpgFVk0M7kKzZI
eSX+AKAJjN6EeQfHGgtJMRKxdzqsPsfpVEbE/z1IDYw3TE7jKeSg8oEAcDRIwVpPooiKW0FT/zpl
ArvA/bwVk5/74Ye7X22t3AP6f43QYjLPD5jSVAbtjAQCMiIq8pCUbXr8CCASldMiGEMHQLIVepZF
ztOf12T8WidoPW50e0NFegpflz7dXZa4Je0lDn/3Sb1pWo3eMIe19Z5AWEcxhBaDSraoT/rewiE9
aEWysK9BEXECQ9ligtBfpY0N7NaRU2hcVwHhqtcV4vqWqYecbPxI/uPtdfv5dHGsl7VF17LN58GO
kVvSqBcpExhs+8hj/AxyLN5jwHfAl81+OqPvOmNaFN6thFZH3CtPn0hb+RoEy0uFY9h7qgajQrBF
9j/kXPacuvoFGd6MmuufLfscUnXAbVjXYjZ+/XI+NMnwRcJvlWTviV32ADjFdBSqtNYnvezuyFCO
Hg9rr5wdl12W3B8k5BikcEEucR+aagQnymfdSruwNRLDVfJKipRBmDa0GxgRygw/Nz5FJXMyH7h7
ajwhKjK9JTS5JTWL0Ixa3jyFJiBqsgE2FYlu3H7kdZIc03pmjHPiKbQcXLBJCdPCseH5pnStVpF5
FLAB1O8GbxH0FcuQXDiHEbUuLlIHlemklbq7XDCj4VPVO9WccTGa8vM7Iufw3qBALahu7lwC8VTI
IJqxPFb/axA/g9pss24/I6eqx02ImazFW+XeKKYrAE9vF93VxgH4wonWawiEGARJUbL20+xvJzSK
Py6KXPT+b0Yv5GzPQA3k9Liw8C2/eQWzCZX/QXXNb0yfDyTDnsxHP8O0EhHdFcRaVN5OE4qgXC13
xVc1Tb6/zH+T3ttnZHs2lmPDw7A3BWNHOU27wLISc4AQ/32MjrN3QmVyaehZ8FZDSyKUYGhiicV0
zk+4nru909Gl43IUptHiyPqrEzMb18SnQDcOJbpKmXWPKPUCzYS6eqfSyZqyKJgqCvDAiBTMhIAC
jkKoszYKAPtkqGbOlwSmjRVGI4GjKAEMufBVRSTEySHY+3nrrPy5ln0zOAYdlhxFjHnaKBzkVjE3
pOn7FEgchnzW4ZNcq0iXpdIZaZG/fbeX8Dfkcv2kF/9ASdPdIv6IIG704Y2Joo77bFLpZAm+CrKF
WRLYbQqPHxSsLk9gwoG0b4xAkuUxJsi5TkN7SHmg0weyibQuHmhrWHVVm91pIqH8xfR5sI67SnPF
t9SlkoONJUgs0BwRiPwuakBepypPwHejmreihRtsaybuxRBNWeA4ow8MwhcLKmNgudCf8N9Eyhdj
gUwY4nbNPOAjRD73Y7NSQmMPAR+/mZGmvETpxMBhIsm99UVMnN8o8VhApx6vIFcme3l6iwohdc40
AXfFk6J5v3kS71DHI2bUp45reuLrC2UOhRXiRoRsYJ29FVuSu4TQrBbUAqlEC5GPSh+z+0M9Gw2/
u10PKE28O8Z8NShaWlCYGM4nskXfqfCPB8JiFCr169ajtJYyrMJtY+BL10rbEQG9iM1yYc0b4+uU
Mb2Py48TznvWsjpW5OhhsJ9rBOiM/QEkW5AIKOa+YzMbNEYvR9OQUJCljB2mc/SUGmHhYH0umGOv
6Tn+p6FjsbJz7SznE6lrVxYSeRVyHjlrE2tve8GGWDUalPVhT267uOio72Cud+bnEAcMq55chtfb
J5LILBtOlAp+HZ2BhnKLEEeNW9WBxy6MxS1RnwTtj2S2QpNvXEcG4uBeYkUyN6eJlgSisbf8l8jU
y8abh6HGFFDYsxzQ4XGe+tYYO66Y10CTqkOBv1hGqMDAFAaJDo3eXSsxphxc0IbjEGnxp8bukzrk
5p8YY9Jp4MygzwF4Xxwbu4A+5e6q6wyXl64MuR7mQOr22Q+WP84fRhqy0GAIETkSHKkGFsT/t4Av
Fg/oXHWBPGl5XTprdAdqkn+IGVDl2DkBr7cgV2sUo7BU9x4XJOqoqWcWNiRN+ppoiaRCXHmCQD0G
GxwGa4m7aSTgrzhioLxdBkmJwNPuJa4VMmc2m0W5iOopbpDH//pLvc52QQ64OmFGB28M9pA/OYZn
4Wi6PkILb3r7y+doHqG4Hw3/m3fVI/N8jF4aZXry9+9YPSyXNSepgjUxmS2wlq84pm3O9utD5K4s
LCJodFDBc/KWogcmG4X94CJkllF53Ao3q403+8rQyFJi3P31vo4RZ5AX7gYGhu45WVM6jjf8HfVt
xAeUSuUnlzviqPfdFpdSTqYKSZ40enFTC5YcS9ZPLLpIOykkt6mFPEHxYJ9l6FzYLkDLDIkDbxix
77qipuKmac2tNxvoGUjpbR55jHHkKlhMaHuxGjNS9MIIPdCdNOISDxBtt8IO8bsZ+elpvRChJ/nc
rhK1A1QMCT7AQ7U78hbx1eG6GYBr9NpzchtXMI5R9pvuA1UBMQh9mkizDyGst89gFf45xUsQVmAQ
I2AIYVCxh2linZp3T8q0yOvQiuiRaL5m9iKvgwB/VJCk0rbFdYFpuFZ/6JD2Kukga+2uEjKFGp9/
/jDGPFuU+zIXVEF/vMsFU3M4B0mJM4mbZnErLe6Kcq/kmVBV44ywD0GiERf61BouFsvWSBKFkvzV
mmYwTqNbWWRLU2X9v9RXyoCLe0Fu6+okgxojKPj6oH3HMZXOW+U+g2nqTZqhsREVxv3S5edly/kh
uiS+cP6NMd/Umky4/QahiCf45w6QDq+Il11cN78NdwbgqRxrEV5/EfLT7RFnRlZToEqKMfG0rD0a
oZfBDXaAE+L+OnswZhQ+8aZQweLL1ngyHRCx6ph2y1+EmAWG7awcw15O2rYwT/hDsHkz8k3fA5mr
OKHow/EegE2JQfnBF0LysENdWyBKno8Kis0UiWV5R3b/zevs2rHyA5GHzKjcX73J2GGcrAzhSEzS
xyuYuQkSp83MYaSsCjUP9yuRf/TLVTOwH24qir7APMNz5vtVchIwIodSz0SNLXU4B5rr9u6RcuGh
UtNC9tdh+hbOy18HMe/WNxgi+ZqO+A7OFPhQclSmyID5ZU9Yu8QHT+705Hdr/UyltYu5BGVTWtu9
f4QG4B0V4YuzzyFT5qy30olB3FvQQTdmrf8+YoDv+nDYx+R0MaX6oVZk36tnwqf6ZB5dLRJX6p1N
c/9Ifor9Swh5GgUlJ1D866k5T3XCBCIvCrP5ppPPEMYIezipZkbBT8lb/6tItaLughFQvzSTFE1b
KvdjUHerVLhp7di7vTXHzVSRPe961MC7GPieprQ6YIB8+fd9uEZrElk337g/HnobabKVS25dDxrj
3S+0ATq5G3f5Pzkzypq7dAGiTIe2GJdNirkKtW6D88E7pVdevE0Al/PlA160B6nq0Aso6urr8kUT
AOUTaMyZJRI59XRvgcz4SRzLY2NihIc0+EAGAKXRVT5U/AXDL06TkOyhMxbPU4ju1XPpMB0ASvgf
kp2jFfOCMz9t6w7MCIxCk86uEx4BiZhJa3IUgWF2ImuAzZ5sVJV9UCupwGNzwitL5UjOaT/O8gXz
2K7G3tdmU9aOZ0JK7oXmeJr6fawbgYP5jUDg5Q+HXixOTBeS8GUZoi7YK555mGhR8d0Fgv/2j8rp
w50SzFy0qWqelxYAvQgD9ZGgH8dxtkxE1yy2cxjoj4v60zbaqBjdLKDxzF6W6Jw/qokVU6DucO1+
I2Woutvn17+9FWGaWFrIGlUfyQDwXzrD7r53wckiAhR3eYNDVd7ecwmXBvXFJPtFt5gr3qhgbEAw
/OLQBUnSKlZPOWD3o3Lq2P8cdDj6x0lwX0FtuF+ewW3uQqhFYiFtyL9ZOB+HkpTWkthbgvAwzs2M
aYLGZvrGpwBz9XOZON1cEwLD4ZHZikWNRpxVEU6mlE82RrloHDPS2VSg4w+o+2GnYCfhlECo0fL+
G+fBw73yCN4tdhR6Wbc8upUzTr88Ff9HdUUhtEg84EfY0brABJ6Iwq32J4WjxDqOM8fWuDI2j/YM
leUOWzwWWMCumNvVb4+fYHpHPE59O1DfZNhyUt9Opz5fXO1x/Uc+P+WMgd7u2q6OjHXGvohIWVsf
GQivTmPxqIWAFVB/++UkX/uNNbxtF6olsxPxfy6Bf1StMPIm8rKh7qvQIfuwJ8+PY0kyVWHJ/E+3
lqp2KczKmqaaTsctPfwRm7cZUwjW0+OLQ4PTwnoebXM7zZTIk3/KtxYGDFyRND/tQxERAd5BlBUf
ToYdRuvjMUm4eJH8Enu4lA6c7887FhoCihtxSqZ6n0cdteqnuf/IMEFw/4cCtlLOkt154ac7np9f
OrtKxo397zbkTo2zKQMoab/4ZAT0CWBJcF8WuEU3vpSIWCCiM4SXyDLQRlvrguPqAuNpkzDVOWsS
QRcIzuiHXs80GbsNo48KhpIQPm0Z49kW/Zbjc7JaL8n8vCcjrk1u/Cj46ZB0y6nlx0KQAfjQuLWC
sOyPgOmTQSEItIPMQ+NfmhzVQWp085G34oGQHDrKuudp5ux7mhqEqda9yCWwbKdpttyn5KAA35oo
P4AbXP3gdbzZxqWm3TWlv0JlYBjniCgoW+RC3LhMMFIO3Sh8outTiwHvvt3LnrJbRqpnD08ic5RS
ok1rh5ozRgW+0x0U4Y+WeT/Y4mI/ZuTLr0Hy/vM55q8RuO4O49jlA/DJ9Hp1hflC0TaE2fJVPudZ
WtKrOTWCTrTkbQTTf7r8AXZwPaXp1KqjGdRj9rVLsLnk2gQ9rK7rhZDw9CCSJSfYQj+drvZVA2/L
QCufbSYwMciaTuzE4yeqeVbPse7jGKFW8z/Z0CjxBsjvkOie/S/GKOtHPfbXD3K66ux1dsKCZZIS
SPuz1xosfO7Ec45Q6sdqd9eyK8dDMbxg/Nxz2ignSSUR05HBDavDKHMstZ/LCqT9vMdUfF8OVySs
JMQx3+wbnf0ZsgTSajpmmu1Ok+CKqTLSSFgtIGxSylOaUxiMCUX/IqNAmKJoer0m8ZnN+Yho+c76
O4x0exNyu5LgpxZOAU57KibGYpqrmyldUrKBj87fBdWY9G6/f4zWgm78QqB0DuZBgr0N285o/kkd
4XjKVY++ST7P287v1GkgLKuFou36ppZgahJuBrTTMlj3AqsG5x3W0LW6bnQ38ECoX7i2/9uCQWYs
vjYu5ne8XVO+6ZILCs86hRlmIHB7QFvuckrNs77kQ5Np0d4/FPLCJ02W2UH2AdHR96T2SHGbAvva
FXGnLxx10JJqMJr6wHSigT4/IrhBnkC8XZ7CdEliuLt21knrZ5rqewg40mlH3EvZXZATUQVV4zVU
6rM63T9/JV2ZNbAJyBMb3X9EGLI05IEkcEqJ5XwrcOghw95PmBL1Mh97UV4TojZ4AZ3bS+8q4PeF
O1ifL74DqSDb9wfDjhL9xwfzxxDWN09beVdeZRwgZNIgNrFwxUzLDeRXf508O3BhMK6aZz7q1I4K
uNKIV55F8OfHhan13bnR23MIx+66AzL3bkul9ok8GtHPbbH3bJZ2Pv2nOQ+yRwr/kLrYvu8IJirR
GzjhYtj/7SV/2dVqL+sYbt2txss3Y95GET3LSBc3wK/JgwiJm0SuZNcKTt3lpQDEfQiOGZohYnQm
kCtq/GJyTxnnhKomkXtufacX6V7UBe5JFz/2zMbT3ehwxKDTwJvOVIpGk1PZ6b70nxuDy51Sws4j
pMcRpnY1asYkdXfntYzxKpuyCJ8lGFzfe9JduY3NjVdexv6YIGUGlqulUOjIZrXNE+lKwc72Hfcz
JrJ4swy2JdxpCOV1Lj3d6eL7Q204X77DB/7legnqhofMZACUbgv4T7rec6dnR6F7s9hLgxbr1qgt
hlcJ0msJ354XW8DJRFVjsWnZN/izFoLB1o2mhn6J6swSwcFcsfN1lORqLYVuTi8q9QaEhlbyhUCZ
j4aQLqoqrO0n6t5o/z3Xg0RDwYuowi0561zUpqKnCvWLaqcuomAUf2hvgQqQVFXi98JXwMbQ+jLm
s1B/Ljndqi7+hmmeu8Mk/2djN1G4/1T3SLGfi4U4v7AhvS01U0xjpwNedqxomUvka/aEUVCnK17I
3qEqwXUVGgGpxSh3IlTPX4gHKlsYyIni8dt4U7QEI9umohfAmV46E74446XEr5CJ3T2MTU7aP+kL
b1PyTbxuU0GQ5zXtTa0kSeLIVSkSUT1PjAG6sm7N8ftry2oR7iNQJ5qGtifQHyjWlacPvyxfztJC
+hGW9s2P0LZkDBHBRt7AxiB8wu+NfRmvmQybOhujFQw9yT5bTyR5d21YMothuHM7QvevX1isaVso
jMUzg5X/M/AGNtARYYLG/XvgD/vD3/D/Nxxn0uCfTc0uZdKw5EUw86r3VaDd+SkmAQp+tXAWZvu0
S/QLjz6m7EYOVG0RuLqwoF5ZQD7jeyBSniiPX46R+1Ywd3m6HxreOQ2OQHpLBNmEim4mI+CEDj1b
tUeCKGLV9UTZMMsgiikUCpQXy9r4o9HYeElG7Dv6aLpk09dCFIdH51ASQYkSp+i419tZkDOIpvh1
MA/TGmAc1jI3gzLiuDL/aRueh94V3XeMrS9YEFEcbIO70Tw+Bi/S6Aoyl/30VNC9sqZlJgmYkFI4
/C9lkSAlGNwvSCCE0hcN4pna6b5Y5k0usm+4jBSX23SoSAnSqA3uicfCtCV1HKtVPFhwq9sC1SaR
Ia+uAMivriFrQmEsaJNN1ztOyVfFEebEkd+2Jfj/dcnjkSL/V4n+zV2j6n66JirYkKKVPReEU3Md
LPfj+Jn+vCXEGWxGLG1OzCMPG9+dTML5TOE5qJr+2RMKLqpSpWSob2qPXIOpfmox41NIntSXBAvF
3AywYVvM9oNLxNDOnAJJ6gBswsjc7ihfUBU0tv6t6JGWPwEjiweA5xTsFrfbFb75BCmnThshbWom
rkDTBJpEo4pCq7WExp3hiInesdzmWP1FiD0W5+tjx3E1BSDpudpspW8fAmD7wErhzLjvfrllfaZk
EQNXmTFvFRJ1WnprS/ky8fiUWguZjL83Qm+blyA83WMjbwUvgiyqY/xL9Xjbv06vWnxYvWzGHpus
gtk059vZF3fYYVPKWL/gK0F/TgM7Db5G9w6Y07RjLBHSvfVJB2zHmvBwwvx9n8wI5aglDQWoQFrP
NuVA0TxBdD75GQTnLUteVDQKSjSuIOwNRTT9KGeEX04vqhFEjf+8/hVWKKPlNBj08Ggr/Iv1Ddpq
3kHhQGRJ42mNNKFZu3Fz0ZPegolpFygZrZDPyD3gQCl3noY7qpfrb/FTzNE5X2WcB31/8OwH6L/A
khTLVGQhcK+nJjPgpUKgNsFetCKPySuWnel0J8YcZxeq1y3SldflSEBoPQxD4PMTBSHl1g0t5umW
BX8IlG9SIBkZHi2S54cFdqrAwZPMAkYYw3/ZZtfiK6jiOCBv84AOLnWYkpOD4IadyxUDNVoV2IHb
kK/+TvKMGbMMCHxLv8Am4eRb5iJ7CgPZekK80byq/LocpOqLBzvF89q10hqn5Xd8Qy29+do6kypn
zcuPfyrZ0+2Cg+veZP/jNg1DYT6Yp+Lx4nMeiv1Nle2WaMghHdQXkKWsZy6dwIoDnOkhkwjrdMxN
mG1VhSNd4avaISHqp7WNN9ZfazEXdrIF14lQBlCzJhkdd3XSCAZAOLY33AmaNRH3LMPJngAogaUC
VtIMEIBSRdkGD4Lm5J+Q4KRRv21Zw0D67ucymdZmn9Dr/FLU+B+/70OkgqnxjnUjc+dYMJu5RGfi
6E9EUUZxYs3Fvo2TObOUWzIKA/uDHlkzh9jvzqpxDed0CTX7j7PW82g1dRvAKRwa65ukoaH7ZUBX
Mwy6NZZXGQZeoDrZa/SDGDlEGL8f6cKpzCxHj010ghaxLJWyi1612LVGZUFcQBalhE0/IXyEtWuM
Oez4URUxXCWWlHPUXQjOJesQVUr2r60eFtncCmhk20hsMCJmId8AErDaJBRN+RqqZ0ozEqHdvwWI
ynf454UPO0V0u/toHUCYjwEgJiaWarxdKzTGBiEMyacugQKTrOgXOmyJwX/fWXHSY1JXhb3Dr+L3
0mPcV3wefdSE/Mgm9Fi2i0i9WBz3HFhfwJQkNaHd4GkhR5z5wyhglzLRhf+hlN8ixDzFxj0ggBSL
z8CxB1YLxthAzUEA68510h4ndf3et3YwMUX0kZR1JBtIrPGXUIG2RcGGgk1Ffcx5EyQvLHFua46E
nMzn/rnDHqk4t4HA21tFF+P3IRAL14XsbG5hUUICB1M2uPyUR+GoqOiJWz+7Dk36YKm/DMZyycC/
S3rmnVF12QIHbKxxMPCbYmL/a3GuP97L6Kh9tRqPC61DtpZt9mEQsG97cvvVx5CpWE4f6U+0Ikjn
E6ORaj/2qLh5tXxGe4C2CY7unQiKO3lX1ZQuwNb3ZPsLvtlG123aPxtOC0bC2xXi6BHFePEZ6DYg
/U0D5aIoOgOE9m+u4LojCsun/xPNVTr/mseHQFUSJyNcAmjxqVRZzT0Sx4AV3FrPL9E2EEpV0ycb
hLEjH8l1QOKmkZetiq1v5k6TmfBelhXyqtD9xUyySp1mTgbi8snwmNfvZzVyEu3SqsDwIqDm0e5j
XC+vzhllI261FTLr3zPQYf2gym3YGXKQOMPVd/OQiJIAQZ/+0S0JQaWbebquTuF31iGg5g0TqtHg
gzeQOfMBIPn/Nrgt/1bbo0gOmSTst6bKpnikToPSV7bzKhZ/+UG/rBEW+7BMAs+jplkPj5cDKKdM
7cygp1JUoOvaMOQXhgy0172y9d0rPspcfPkHZdujIGaR6uwQZcGSiBoTAtTFUXcAYYyKJoptjwek
3VG5B23EkUfeHhB41unczIZ8z16nDU9OwIbuWE+Ano7OSO8UwW5h4+j+oj6tze0K/GmLDi1ExuQt
KR7PqYH1IVY+DgtBWBr5McbddTTf8z7iw3OfCK3IjGMx9yLCU/+6mfuQyVVf9HCyK4m5tHjT7aEc
dqBIO9VMgBzByiEMWDmSDIFe29Sx6uqSXvJbWHnquJfGMifaYHjs0rB2x1A1cWcg3LGzlNxkdeCE
LQYnL/48C9gYojCk81p+3+MQcRVZbyQN2JquQyz8chzrFH2cUkZsWGhuF5HpKXwdUGnvB3F7oBJ+
/qXjq0cX3dvlG9LWOXTLPVCpMMQLOTg9NnW6oxIHuGNsE8yFiQhdFkdK3TL//lD0NsKwpiALBdLs
GO7UsaQvgPeAc40yAaxrp2FHlo+s9hprVZtKcoW19E/8s/cZM8YZQZwkDnDpp9POdO1tski3TnvF
S+8LuYwo1S3wcj9H/ubxM8+KBq8PhTJlzKbNg/kByos98uqa3yO7UynJkFQgFI3f8WbdGRVcV6Fm
XtBnZjq4UdbWafeaF7eLEjQKTdjSrrTjjDsAPmNGFYwdQrysWgXzCOz7gJ5f0jwNvYaI04YxxUs6
HRZSrbBR0qtHLeFO8QeqbL00ZtivF1WRftYMCO6DNOKW3chJkt+tY7KDHhgjp3U/0CWnvCyFUovN
Lg1rmq0hscib0vChrunFDADboyocROyKJG0fuKKvz8aN94KrwU0fAOc6oUW9h9EVDn5S2Uce+GEH
k91yr3/qctpKi/FiZFzyq0C1vXzGbqSFWfj7lG+Ljd9nqVkQxUCQo428E1cBfzLZzjN6HeaDNxSS
aZfV8shp3W0xv8POHirkL+oEeSebOOvQZIqvR8x+7vbTbmg3WSH6l6nz1+/nODAzwyd28F40wKpa
1ekwgy7j89WMgsMnHkg7c5kLQkEuZziu62RDbMMfIRVzaPeg7oAZcMGfZXOnfVgTMHXZjUImJSBX
Dncl0XqzqJgQ+7On//FhiBJynOQKe1Vsd90UyVlrEkfhdoccmAfUIihjybY13syzS3HuTT+AnPAh
gtsVEHvQm7Yu7skp//F8Y+9VxJ4TdRNK+fyakIyjC/DbSe7bBVRTpz+kvkPOlLT5Sr4w9slAr8bV
kzF1p9iSV3k2ROkZ0o+/xvC57wlURfKmFsW/VoP2DL8uHjkL2HhfZLrZhiIaPlZxQIZHvJcZJbv0
FSp0sbhLJ2bK45Ng8yt378hhi1M0ARi39A1NmC1AuUb78xqIRSQkh2XkNPPbMXbk8282VCnUQAMy
+NKXdmbnkemA7i42YEDB/oKaFmnuqNdSGTI0mbhlMGrzGXJa0Yx+ESiTqNeKReGK/pDILgrEwF5E
323qwao2QNWaou/9wPta+yZ1uxPmr4bXSjIlXOtKWCeO1/s5hqTyFwZl/hpy53Lybk21YNPBzCOB
Kl5ZG8skzpxjF7JdR8e18MHYPXe0PzxxFPGPyw3iT9c0IQvddGFsNXAW2eH+9ObG6btEsysl+m3x
SRuiaabJFVWfFzcXGHNF7xzbeVDypuAk2zeZHtJ11XosrnYTr8/3GnTkAK68XkQWUTnlXcLTeTX0
bC2H5e3mGsPjB8WZYAeRX7l24Q4sV4MCyOKgEaunbvtDYP3H0PBX0nXcVuU0b/nyW6CrmdQFKKQg
FgmeWTD8vbSGLP0nLt3oIPcYaSZO+gFyWyfHTfd2Fd8TQ20eGaneU/28eNkueQIWkXf0w0SdVELs
3ruYVZe9LBA1g1LwLFgXC+uQYBVTvGtZh3rOZWbRn24dC5D1lfm/kekXPi1l1UVYzALDZ5qEm8HH
BLoVclxs1ri5l1yt5/9ICTvV9SjKpQEzfAfGTVMTx+WcBBjzToYlchwNZd5/T/Ob+SNk7cj0PYo6
Y/mLhQuP7ntt/b7IzzlueINsdjAN1jBra/wXyCGyBKrjNY5Baqyn/jgPvgG9BPv3r4NKJeThL/bx
xaLbxpryzmAXIB4Ta+o0IhoUOHrOVRPlWBR+xlmVd4OBrZracOPavDjx5R14ZTAlD8VZ5sPUaVj5
E2htn/+Ust32XHqLo0+nLipBaEsL/++q3TjRKb+9VM/u53pL/ISvNZkf84P7aUdv/VRolQhZLFqi
vnYkWTGwdB7DIJ19wy0lKEMoI59I9h14COZSWl8OfsGmbWVCkjivqANhqWEhyoEiUjRIV43K2cGQ
qYE/+EFweAdX5oFsTBNUZLl/Bhk3sXAy2VxH7WAqcf+kYJQMRSdfn6rxnGq7UgBX/Jaeluj/pfNS
unBdEZAt0cXXtAdsosMXv+knwso9cwpiEdj8R+edwBfHYDbbnZ48zTrLSyVzu9pFSN/XhORWgf/R
PHIjHKV6i2ZNxzznGG56oqNjh5pV2LidfWK5AOoJF22L7NpweHOfpqMiuGuyIHd2zzO6P3RSrKQA
ziBZzBHA7nYNEMq7yCm/rSk00GrahVhl6aKwovk9Mjt9KB4yt7GRCXyBDcebpxbR+lLz1ZFPEp8V
EcXcALwaGL0cWvUGnj94E6VCSLP3RcYiWZgoWVLHwipirJxu9bEtOVN5ZMOXtxaOiNzx7+KtvyMU
6sHgssva6ozAaNLj1UiugxixvBo9lNAT654GQpQ2dGfTYS9MezbYAOlHlLt/1fgbwUxsWg59UICn
NXz1MrPCKwsFLri+V9IVH4u+L6KZUXTXHZOvQfY/yEBAjbLPa7jkPPsORHCVyWVpfOAqMzorbZjR
cMOdE+4WAL9cCJig5FAH8wPDRYmfOCwgp5TwKqKFAqWnPldw9amSOBGvxTBgYZRc2N1cDIBraam2
GzT+7biLqoqqvwSXIYgKoYXQIRgGrOZXq6/TK0LRlkIK+ntokZBg5+zLrcdJZVNRM0UPubFY8Bvs
YvC1v5zLFOjvkN4eEbK+10l+sp35nWNrDIQPf+foFiEzeMvFa7TbI5QtuPx+HqauG1iRVVBclDxd
smdlqrpGCQuwSjxLYjwjc1cNTw3wBmM5XguJ0HwWpu/oxWf2QG2hUG2ecs13yaCC2OTeHlrHHZwr
iZ5QCeHeuWMPzA/6gMfeN3Ge+0csY6HevVy6QROa2Ku3pXNQHDqG1wXbpwQvtcdavb+zcjM0O7MU
si/Fo9kmcD1+aOvBOnXXGeK2aCew4e9t4hLkZQ/C6CmlHL7zVnVDRNk3eGMuAPRtLwMui3BcjIA2
ZEJHmtOyYzn5TXf/mzV9/PUHXuzWi4lFDC+QHi6yjDH+cFQzmN0cUTqwxU6GVrShG8NcuNbQIC3W
N44GOz5tM2fEAAGNlAowxD1ozIZwmGlwRpDp011zplxmNJs98+9RUdz6T8A45KLkItudrRNV673W
xK9l+5qBkNRYl7e4qdGG7PBphC4aG+s+SPXw/y2tJKTSO7FQck6uoz0V3Lla58O8QKTNnsgt2wLm
XyJSDDoaRw7r8LlzpChX8s1SRRFf6MU7mg0cw1Q7jdnHmrZniM/gjIVdqYRhXrOLS4Qe1oeQnV75
kZiZId+tSGLn09m/FdJbkFRIEB4/Nn/mQXfVGHvJ7dqwstU6hof1pLDLm0Qvw/myWv8R5+Y+9RbE
EG9iz9FDoP0v1KrZBimcLRhHIPK1/DGR1wty8NrAsgTC8IqsCIyba37T7TeA+yCT/rnHN78mcOJ9
+c/XbV12sKWrqQBuMp0nO6FoloiVi788SVfsFMA375floSM9zJ4zCKyuprrrZyPf8MskW44sLgjS
qLqPPwT0jYBv/QSZK3aNBFydAYNGXP1S4/A2vN2/M3/kj1k+oSBFn44bDgnt4VEXDOXGtlWmv0At
Mx8YccJ3V9d6U6QnY+vNm1tE8iHW4N00mZqO0aEi5PocJtwypwkNiiO21k43VkIp4Z/VcfF/Mxl8
3+zwM3qF1z68FdxsoNW/gWxP0xZHo2CyUr1Om8xGxYJRdVW/Eqa6t48UhhBl+h7910N2IzqSzt6h
ceLQG0DFEmIw8osOANSCawwbvhbDeEDUCvvE8qBYp/F7ig+XtbW7LB3xYu2yy3I5Uo+KWEvGKqR1
EV+mTEPLg5fZ04glLsErl4OCfpYaEyRVzplmWrxry14bKXb8ul6b+7c+R9hs8p4sTJJKSDdlihNx
3TG2EbFr2fC87fTQ2juokCWJzHEdWtdtepocpw1aWFvGhqVjuKKV78z6lYXfGlYl4Pbf7RbAHoMD
byPZuHellaaOHOFSBCOYTtDfPHGnjheRwCRwKl3GspXHRaw4XgKqj0kmoZ9N7UBbuuLOJbsT3R02
9S94qe+LX+WgGG7CKRZ6PxCloblZ+17CS37pukcLAHod0AosM1Vu3E+sX9120n5ynANZH/atk3uf
02d1OKvG3zs7m5JKq1JM2Ko/64xKR/JaiNhw3KwWtyj5QpKHKTxfvyVupFTvjdeqE32vauTx/56B
CPWitbMYM0YusbhMqLPue9o0HJlrBcm3enULT8fhqR8tlsGQQd9Gb84IQJVJWZpgAtyk7BBLJKQ6
zA8UvZc7uV5HUOGrom9cxwd5Y8JWiTBFD2cZIccopYIhm2bvqSlcvcq0AEojIZxoGKHuPI9Dzgy0
TVPlcOhYttqOGLf7FQGcdwvhJh9NSulcc/AroYU6f4/ZH3WpE8zXThgbZjIua6o540dLQmKfLSt4
iXk19hKdSUTpwOC8cRWJraJd0oGp5Nm2IxYfQPUr7Tm291dM6fIiRcgbMxFSjHEUSYxrEIaPJzB6
I1DV9cD1VNECmLJAp91yjvX2ZA+zGRHkryNV0zL5k8LmVU5oLCJc65Rh5aUljEJbOheQ3wUvtN6U
FyRs7QWE9JxBfWFD/2NCTdxdUZqORxq37lT7d879V1JVqFg6b05r3Q4gqZbABfs1Rt4Rkl4cbVe7
L+BSg4ZQdmmQY757XX3NQmBG+nNUjLkDmrIH9EHDY0WQtewUJzqK6m0Ge/cbCuyaXcJhmvZHtk9g
UoIjNjac7HLAxeqPky5c0QXY2i4mhXWEDmQDO/J3dLQX1PWFIQaFQIuGIu4REqR5MB+4+yJj364x
IKmwFUfK4WbTrhDgxOr4F9e2VlDzvntDlz3QhZqlO8fivthKphs2a0T9DMIYWG9xpG5JmN6Xm/HZ
MQVkSYGwhCE+M7pHhnrI0c1qB3TnSfolnytCcYtpptpD25SM4m6yyS8NCHFTwi6lZZ4aKg5ZMNSP
0MO6lDYJYczgYIhLr05Edsq6W203oYhEtt5VDf71cM2K12lyi8onLifq3a1s0RGSCFssTq+PvZ1W
hoNSFbigk8cdXD3aWNaWPd5M306Q4hPqq8ng5n8uv1jT36UoEAPb/nN1zsr5l4DOksvwRwVS/qEI
XQUxSNibiM6XgfIT0KI5HVNqnrUqfVH5/zdBGKcSabzpWCtmqEylYAvtyDKYoymHZh1jFy2KJEVR
Hw1X4vNp9Wzrarf9j0PQbvWwfcQ/dcmSyfn+WiP0o4JVgsz5OpfxDmfcF6SJ75YIXpQVCe92jNtv
hkzIFJ7y6Z4su1RsNFBFsr2FN0h2JFHesBr87CTL+6snou7jl7k0rv4w0DQZ8ogs8R4FCMQp+3f9
X+j5WKkxid+FuI+3f+TWbCT2pQCt+WHTxu7rEPWA7zhs+SSOK+V2bynC3vhWrpuJ4tN5pAOdRXPi
UovUlsYK2hoEp5pxnZaxyBOZBPiPWLMOP3Ir9QDmjwh7cqRWLSRJ08t0ftXKcNg2K2Ar6CivK7F3
2C3W0l7MgCYQjAtMQwEODb8l3+t1U2zP8A/mKnSb56QDc6JNwZuEHy5Zq5phr0UencgtiLucTFSt
0XBvjT+Dj+MC0S9AtPZQM/qBjTH4P7wcas7MNuDrG43CvbIOjcU7/j4vVbJTZo4sgelMsnf4Olkg
xckOWd7NPGIpRZ8F71fF3vxJFzpSMnKdeiCZNYOnHcgE9MB+9qb9UO3nsNqYl4qyMOW7mttRsy5q
VzknA3O3efQPceHKDWmoh7MTuw4VB0yWN6NjmZwBpqPus6WiT7j40wEcBEiy/k7nomgAVxDVt7pE
d1i9JuAh86hb/Uqf1Q1hYJMYvMq7KTiKW28/tQdUOVvv4Jb07VJG7mK2xNXoP06LFVQ6G7K7eW41
6+3gH/UJwaWHJPMSoP3cMkZ0rIP//b0/1X7yrDWqK9kJs4+rlqVDD7kO6/UU8olgXmUM3aY0TysK
inStTFeXjoAAVk+w7le/oNuV00OzCywvRCyWOJ8jKsOuPxv9LUDLgDEDhF1ZKY3DpEVzgpa9dsKa
AaXfaQDg9MaF+FEJSxWHDJqCoiG3huupTQNNPBwpOf95hG2PPJk2eW1bSqFn/13GOlvmcVgckpQ+
1IOYw/llb6ngxl4Useo1BecG5ZV73KrdgfQFp5jif7JW4iao7zL3/8denC8vEDALq/sLEDISIRpm
Ib6JVsMcpDFIMtYQWCQj3UB/PClPDtCe8VjlHQp0o4Ie7v9briYowH5V+6gNWTp3oC522DA+eXpk
o3ewBqUmrbDhMEEcmLgec4TgancdLerpMmwVvRoHEdsDz6et4xSWI24N7PMgcolB2708Q9l9VnZy
ay/cNPEPQj3HLQEUU3YQ4+t+LgZya2TykRcHv0hEnESc+U1kaL9H4mtz3uerfzwGr4Qe0NdBJzGC
5ocjI3Ht0nx5K1E+spbOSYuFXSL0qsxMDheMzUJ24i5WtCeZ7aZetYioA9VSuTS7FM1tt/fbolBS
lu5D73q9Z/6xjXXJuND3pKvku+Y/EsvuvJGW1J9nf8lLNfp3by7n4NKCQhMG3gK0li37globZoD6
qmW/vjVNXnvg03+5SMp+ldl39pHT/U9ThVpv6S533PdgrKPh4NnuEA3zodoTCaAPdUb3OJHI4TOq
75OSIWg/EDlKH8JZ7CHaRuz6z9IzG7OWpOYbjhiSFCmoTvdckaBTdNaPg5aHxGGeYt3NfstO8ogC
/nV82ane9GYNwYEwFq5/0CCno3jixS83Y97FebUOHO1oSgSGtj2S0nm/mUwkdtsaYxfw5VklVqPQ
NoO+Vyc5t6PyltqJYJjLaGtokGW2dVfOd7OhvdMRMKxj6tcUPqDdD6BetffW6cMSt58jU8cNYAgR
elpEZmMQtYkZcT1pDYxEuvvFY+pojZeXdaB/C3xf14TwttDdfATOXqFYZ/KqKtGR3stNfYCtjwYP
R9s8jd8iZQGVGkSOthzYFnH1OfKXez1ev/gDXkRY5oQgpg5KHrGBSI1IqR7DeV4VNfuMi65Lsbkh
zDnGkSy9HPDdkUGCw98tEi9hdW95mVOo/opeh0j25UD8m8bfBjR3BtbmpJ3FH7upzKJK8APZ2wOR
pFw9BVC18QMPZ4HgHjB2mQMhT+HdN2lwnBaqdr7vxFNIOfHl3AByTtrBOwx7o1NfjwAkA1/U8fX9
47AKecZmzOzYTQvICw7sHyeK8Ubr4wtj/V9UW8Wn3SoR6WlXa9Bf5FtOuQKJzuSVf58/YNERjWuX
j3UC80A41tnXNbOV5LCrYAyxydECVvbVTIegxLHUs/E4kCx6i7jHP+CBl5yYEmep32tn1FIjtNEE
tZvAcxndFagB0hfjVBjIuQkAMKkDAlG9wPbZADseoyz0WDgYmwmunARMHah4Ie7uxfekaNWhQ7D9
1wuB8HJX2BGVnJ/g7cfScU94ILJKO5Ky368uEwB34+BMbGZJtaWVwqK5cfHmk6nbxz5+OElvlckv
OiQ6OyDZctSgCqDW+ADETFkbABJ/RVnw35JoRgdbL70wFT9bVZ4n1OC02Nqsu+Pu3PBk3K1GTgOz
Vr8J55QDbTh7GQDrn6OwTCef2MTB2Cfj9l1ElLR6se3IwEZFh8GCFVOfWr6aWVtNwWvGa7doWk6h
ommIoNyKtxl01ombTMFPhedEFGjQhpaWg35vZjn8Obcj/JoEGfE4+0sKOKT5qo94M9bg36bLmiAq
mBUOGiQKP/h3UVgF4wy5+k7U5vP/h96QhkQK7b5Qk6ioA0qMN/K4Mi5QGZH/noIEe++G0+H7JSWo
a/RGyA+3JFCm5CKz8/lrALMMAbSne1jl0B8Ayip80MY5hcy9rBbYrc13stEVsVcq0UBVrZwRciL2
btpjHbnklEeujEnsyl4piRL96xWLrA6NrErshbZBSQxd5QqXVdcI6Iht8wx6UHVtxW0LGbj1joma
6M042iRPB9iLm/PhF//N4m6qYX5jF3FbhjKp/k15eYZJSPfWAsf8FGcHsgcPZiEvggZ6dmYZ7/6x
s3R7RDM9WckSaeIUj9Rph+2q66PCzoh0qSY3jbAL83ZxMFSOamIdSg/eZ4xWBT5e1TgMk2arINFr
H/p6GhlZv4JzEhpfWCstk7bMkSE6g0LP0TavrLH6mmyEOqdPoHHnz4aZbtLDx7oB4aIB6q3YjIaz
pVi5jNb12TxPuiktJ+6y+myP2WfbzF8bUuwjryDosoDOmTtCBj6Uyi2kuBR9mFR5XTn8Ws+yRuac
VkFNgoTZnSxbhAhAkgHcpu9wyIA/2FmnmQrxYglF3960n39MKIfCVwysG7Rc2T/oqupYiXAd1Z8v
fc6ZRyRVRjV3R8eV1P6VBajhTylDuxPwM6mnDkQGTDUrDpAJUd9kxOr3n1sbHl1sP8s03xIH9nNR
OMiwXFZwM6iQ8k5sVe4tZO7ab4nIPMzVfk8Ci63srUaXfcz1fUMveVi0Wy081YE7Z6sae0PJN8N4
TtCNRU4klkKfSG6lutt6BeFekONyAT9szKnTVQwbbRYFdOUQw25dK2dz3uqv9JGl8cZ3zVKTRU5d
L9ekZ5dnhetJjRJqmjnw7ylD+zuo8b65SUILD7f8yACvjqtGKMuydHGkjGAcra2z1QjF/gC8PMNo
hawPlB4dKHj7P2BFw81zMAbLpmebc2B95IlZfFnvm4xtFKyZcPsRbvP/dqFbVc3uuLHZEeKsrtBQ
DCBfhysUwEdNgilhNxcEyX4iFH749/OwtBYTuv4aG5tlmBEAzUTsz7zaCUfi/5f0fJb7vx51bPpq
c9JJ3DE9W/tZrfNPNxPcqk+HH1Y0jYYg3Ct/aOZmMmHJwMCXuZUGlIF9+Ef3zC3HOHRDReONQtUA
idWIUBLnrnORKBfSHbiOGigjprzEeaEPkiHKYbTEMslDTi/E92t3v83hBomiymU57SlEB97qt+d+
D7juEWdy8d0Y4AeJlwxsiKl6PYroE026+dBo4tI8U2Uy5LBlH56Z84ZQDODu4joSjmUhonjWA7E8
m+oPoZ728DUZJeA8S0FNyZOgYLSkCdObuXWhnYa5JwbwX4OinMrhY6lFDvsitAvl+cSqojcuGsT4
zOHgtGPqZ/aEXSYzAWnXtxoDvnkuklBGm9YxCCsrXfKnnWl1CPV+kRczYa9vVMTPE8eBCvUmctMG
mGVcOeIoQoPWgnkdHwD+e96NxHZMSU26w6SNr/+RzT6qk46uglSXY+w/cc4fY9RgNNiRhJCrdvzD
bqACkAKWbdwm88ExpAJnC115wgdpl9xpB4GrfsFf7hgpYTmpLJgcDNSNhleXBxFYRh5PxTiNKRsr
06TK7Hr0jKc9yZHNi0lcz2U5byF8QIkNzXt8hk1DIKLOIKxFI6sjTZunPK251pXDXv6P4ZkFBVz1
YhQ52dPdk4EAisbvA/3muj5nSalf5O1k65DUBv9+jk1YlJ57AyuyKdivUekWrhDP1KLTw2MVBaxQ
9I1Hkp6ai2QP8EbWKRZSMTX8z1epgxqJz66TTqqC+bAJgFY8HVJcZzLObkPRBf2gXFEvUGo5AwZX
2f8YxNBnQsP+qq0FYuX2b7HvWugaWO1o73HDBDuB2IwpJrec+NjjGVtXXFV5MEWMiMqxmhxb379/
5LSJUYHkXjTOdmi95Kwbd76LkueVjjw5NzwyhZR5BzSxMKwgmBxcaHIWduiUvQ+NeLvWerPQ/KmW
XxDvs47Fkn1HNDeNxWBoCUbadAzDqsmA2rB76Q/4WXCVrgUxo2CFza95zNJDeuL8tyF81DBsG6n+
1VI+oUoRT3QbRwHr5Nru1WmmGWxK+W1Wz9+TSMMdl+nkPPO9rLoFDqKQm2Ns+cE2PoE3uFLLbepf
4ig4Tbd0bOLDwIDcxMtIBk0QgR8djiVD1H+ExjfuC1xJEY8dqNRTy3omJU7qJPbllQVWWCXuC4SX
IVdjrRJmixu+Xg41D1ZmP9y2itva/iBtPq/u+SIlZmL3KCCj/geSvulpb5DuqrvkY8uXOFXoCZIy
3aIHsMc1w2VoBpH8aYHO4IRAzZxRYRrp2KTOOIMAEEVUo2s97m1r4v56OAagUN7BEAyFRpy57tQb
yXQFV9bkGtbOfuvGFrbnNNaWTyQOkUO73NDWb9vvzngEKaqOZ2GNYV3wPBkhwVVjrKdd+bW3z210
eOkikoaVK8BJJc3FAOHtOaHzL0P5tvU6o1hsnIw+m8PBErmZ9ih7tqv4c8g845kX7oBWut0s6bUk
5NSsxCuKyWU82QLiYLsDsQ85LwZf59CUx0cdCXVWv0gh6fW9Zyd/LZHR/2oVYUqjyl9kbuTEAwEv
io9us4aTN/UF5s8wblIECm0JJ0GmQk+XmFE1JX+yzdV92MGn3gG9fwhWXWY2jOHgbpTBeKOaf28R
S3HG9HNJVNnnbwuaP7BS4+nVYi6CDBv/Kqwz44RzHTMo/FlHrlm/u0XQBIbNKHy4Ri+GiVoFTLWP
QpgBs8vEFdK/2NeltfXggsSA2mcFsTl55uD1ERAAC7aQnbqTmCm5yXhKunxnFN8WVQoEPhBlSt13
mVH1/W1m0t58pog0rSDw2+a5OImCDDUAbrr70AbxXrehwm3QXTumyCH9EpYbnAo3SXPd5BdXuDoP
HKY4nFftYESmqZjdsQgMhjAEA7p/Ta/QYFde+4jIRbQmRgVyAnudVJ5g1VI7bXWSlz0mUkDXbIMO
nQOAkgSUqysR+kCLRSpQvGXH3vH9CH+aFa5S6jdN0idWh3wcnzzhsBQft1f5y9/DC6AA3tj7zgs9
wDaDWpJlBvgpqRlqktAsntEb12s1yNTPHjlX2IilezKfhXVqnxLEtoR0nP9cYDLHMDKf7R88/kzK
Qkbe8zFvZ0jxOqHAI+4bZqmEd+dGAg5PZeKxBNI1Z6V1BsFoy9GvCTmdnu0XsepHSKkzSAC7Mw7/
ejnWf2yuijobglHRKu7GMZ36WldFEXVQ/flowY20aK0yBzY58UUtGV0EOmPXixZCGbCxs2E8D7Mw
jsFUWOztEQLm02rWnWxtVLbLi+P49OA+VHTBLn5R5UGZFLCG8DhiF6CVocYSnnAZEHrLMIcAx31P
cZMs7/cP9Vc2fHp4xR+vEPPGenPTHeT/GTvq+LPNsUxQJ96suqqX5kxXYdX97cLFjAQU4eH4pPlP
A9yMpwtd7MPEJ7O70tEV0+Ak0lepXKijlpBJORm5+U0Nl12CArepY3lf/7UqgyxcAyOPLwXncf6d
LBuA/FP2Fi2WluQvxFdOrib9K1jle5UIj7s8lz2su9O87BVwGdzDhfjCYmMVCt9p9BHh7C4doXiM
krKoXzZMxeQ/bNM3c7W1lHGwLFhFLuNU3WQRJNiLQiaSqLbsO2n3e56qxj77W4X4sYVZLqskdwWf
6a6Tn37/OhEvgDV43h/FljUkwJgnGXkebjo30ODKQQAHzVJnJAI/TOiucbXzUPfwkVIWE6Zfqf+K
0KFR7mfzeyebWymIQxYrtg2gyyKDzHXR3Z3WhylP/Vz6o04bwwMcU1lVgSe3uKAjVm0VYw9nA2lr
ajrAPNQtUXTXmnHcbGAGzqd8epnhQ9f8dAvdNeAeOBaiclUvzh366HVe04//DSumO2+sP1GOKKiy
1Wrqxn9eb84EZGbiNz3SOVLaCkgfwKeYmKRjzb8uerp3vhm96WG8zOFIH2E1C/erusJi/e6yMeD0
BTf+uxA1GYf7nSseseK7A8vDp4r9D45QtQBkTyUhBUrTx+JQPX3h/4L3Cuy60wMahlESF81Ltid3
Dk4LdKYAd8IQLWWQOSXyV/tujgNs6qaUI2/3J6vj/hwVLOV/siefoESE4JB1rjp7ceGl5opIIIsS
HFHsKwc+qPAmbtLhm4O0IolQHvnXipPDcRFQ/WIIhVbg+s9LpxUVGnBEOpslzDo7NOWENmMiTCOb
h8ZzLB9J3hD2htUugplDi+udXISOYh1/UpYvZxDZBQ4h5AwlHphXjcUJqs5cSQE0ymiH1CfrPtGU
uEFVLWgKSgf1pKIZTw9dl6bwCLwW0XEOsVwDW+9rSYyBA4w6WW8P9RkzPQjVhsmU7eTV9lQNnrta
UwgFzrKwTE6PncX+SB9Pyj+uE8EAhY9HSALgsPs9425AYy+uXRnPG7Ci4DNDORdHWg3c/fL6LdYH
1VFhU5n2CPXD3eLfyabZDTQd0pYBb6fuhvJyWeRFEZU32AMXFi4s9Xa6dGKH6edOIq8dnwsaahjL
8RTv3G1fKxD9zqpu08oIzpXUEnze5/X6J0W+UXM6vjLwUtASSM0gMt57LuwuMSkSMN854na/tAAg
fJ3OYcZOlQEIrXltUiIDtTUeWd86oe6lTBahsoLUUkmUPdmGp0oaWB8mIH9Ul+Mu8aFHHeRN8wsa
BK01Vs/ODOfkI7qUCvblXA5Ws3QwKJ8P7VQhgIAOx8EQm7VTvqFOqoW7gOUt1e8+L/bcMd4px9sO
BBa2C4KKa3eZCDDTCUloWgulT03Twl4P9WrelyN2z6uBxvCzPuV0rWmWPIij1Jr+0taAd7BRtR6r
BywZzaHxClGTCo5Ft1fpMPutntcqywwFqSv8Lxf+ZcGxR59pAkhdwYQkTDkhLsCwBnL7oDX4t0hu
TtyFOEMq4goUAhRoW82nP6gNdxviX8jyi8/A32slg8By0zk2AsLa/GyHbWOdcPkLz5EpzvS4rodY
AmLdNRhj7u64B1YWM9f31TwCH0lof8nCxW5DPFOVeJSB5CfpIB51EhSfQd17Y+MB4jwwORsV5V2i
rQoHNiC7DzQFc3v6QRvDy1o5LG05Tz8LdAGFM5w2kKZr1+pDuq1ihFTqtJ1gKd54fiq1NjgNeiP4
2GavAV9pWxBajeMoS45n68KPurhOACsrTOBMKJYST6XuftFwKypLCX77rrutybK0t6tFc1WwaGEQ
0s5U6TemUTZplR1uqMoeyObfNDvuYHwIWEcj2J+dJ5sQ0zFciO7hEq7XAZ1JhVEBF/mtgXH1jbny
t0oWoB2uaLAljVsuhpY/ogckHZYWu2zhuw4zndvEHQKx6kp0uIipYTnAsns5av10nl3oF87hUl/S
ZCvbpyLvYbj3xzrxJwobW9R/hbEAKKkplte7dwqfr1YMgt8/lxOGBOlTGLKxz0O6z7/o64098KlQ
1tna4ucxjZP85q6FOFi2WuKsx1irw5ekswFDITvcW/RzKzOYmrb+HFZjWF7LzMIij48HsipiwLDQ
i9+EYkVxYmsz9cMJkp79AQlE6W91Me8VeRlc2ixsn8dPoxn8miyiFSt3qXhktdmN5KUMamvoCS20
/fXAWUc7zJSzDDv/jRi8wtqTwMNmTO3tkyxEILD5CtUv59tXVenjj+/3pTCcCyyNZbzZIA7rAagu
GNikktNifUJutMjxhe23LARHl3+tl+zUqHQqVYpHG710fhOtu4/VZYHSSHh9zviEpL6ITzFlRzE1
dZYD1gegiuhiqmBLpxWUeea6T4Jxg5CuROJvCbmiAgXW01Hv15iTTt9p+fC3zBKC/nHRwgeMcFBy
eFTOwiYUQAQ4x8xT22RH6fxE0vG0HQpjMi4O9dgc3u+9jdi7T345EO/nmXtPglWL7htQk+V8CjBo
3f6FA3TbfuRst99FbChFNSnSpanzRQVMhNC5BhQilQVVaVyBH9DRuEtPaUlHnh/KDVgXY+MHhp27
QXiAAR2NO2+8X/kw7TEuY5HIj6Gp6dHRXOzb2gMCfYx0wrPm1j9H/VI8JUQexqmIO9t5WJHZizKx
nW/3yYj9En9I+hp7oRH2PLqbYKEKxthjLYDz4vw/mWqMdx8ArBqsLSpYzeXA53fSVl4rjqP+V3Zd
gOSJBEXH7bHghjQs0IOvrAtgrs7v0V5AKlC7Bv7HcMf/04uroeTH3mRDcBz+71zdBR/EgNBiJPgN
Al2jwvdqvVp2Fw441bK6983inTwe85kovjtTkAze5NlIIWcHtxJWd9meRrnNfi3/Gmp4VSptS+v7
rXliaujrf8M6xmJyAHNBQqOegVwhDAQs4S+z5tGbS5B1uKlEBMPghcWQrjcpG4kFdnS2RpFrQjQI
xYqndam/y1mj5hxLi1zeDoCOkpdmPMKBPDtLGTIUO2LEGnqr25l8ChK2wnGJamoRDm19FzozMq9L
ZcY49+pdOIAXF6onKGHnoRVbPC8MTVb4vQG1MeDUHboxAgQ8bCXu/mIIvZATxf6JdTX0oVDU795k
e34wUaLwE4+7e1mhTqZwsyXacoLQEl7y+U/fkZcWgvQ14WryHcG5IiF1eiyP8Rn778HDHgNHAQl+
NwYVz6ECKa0ATc95P/gdVonbt4SiAiy0Yo12HxqS9F6AiO9OEzacGex54siFpq8UPxOVdsUSfK5G
JONGjSc7ymju3QEZvQcNocu2E0AWUeS2ofnmCSroCX2fCqwnJifttVpREeDhbqPjceoSNSr4ph1c
ezEaxSwtXzaEGIFqUA6XSg61uQzQ0QfsW+24sDJItvCjuTzJQXjzEIy+l8bYGFlieAqDi6OLFLiE
Fn/pPvCGSNkbFHUTcvfCbN6c6mPIZuKFuPcXQ6opWmdVkSRmViywXdG/LDrmnDmMvXpbbgEGBc0h
IW0GW/PuvwX51abTVl2YsYKgkkecFXapzwqA04WWGFXJWkf39QARa3mLG3A4JB8UAwYRkrK0n0ZI
bxVOVrN9+jWBjOQlDW7PA05RlLfxFfoDVXOPsBLR088SXd0bFAw5YQiLtVE612qVAfZoMSBrHYID
PTYz3iJGXcSeV8cCBzA8V7KAd2i/obMaFcS7PAlT85nA6lR6ZvTtXBXg2hqAl7YQ9z4fXQBqM0K+
K68FM3O5LCCvNbsoFbyT+6gotbAsA9TKrSCV/8C2h1lHqXwppFwEYBSk3+5dgNEb65X8X+rYi7A2
Pa1Xq8kiRq7fp1+p7hwio3bbiqpSQOq8YLt6/lqiu/0sunKvZeB7GpX9plqg4tNogGG0tq2enXwv
WGwlPWqT0nPXzUAY7HZ5nEZ3yNvOaj0GGBiq+AgdLtA36rQzGc3GUJXF3mhMOwkRODBua5No4Sgn
2prW5XKLjxhmq+plwUHzpfdPnGgrJWahaMKA4ozSLL1odOL+NgxMXVFGOEYvhX6648b6uhsTOQ4X
VpwTdLpgkho6b0h4ekIPEbUMRZYcXDiy7uio1O+IFDYSkBj5+BB5f6xtUuTWewdKjna1N2eUUP3D
NsJRW1xPqQvVfJrCu1PgSfZf2YBBaB+1v7q3Kjwe+xPuhF9BnEgDq9IqH7TGwekCyixy6YrorI8W
bHHs2Z6/ZWIQSaa4u3a0bh7CqVxxaveQdnjDuW9xycovoGv1jG1ctNpCFgYi6SPvBaKqjHPIs9MO
uZ7yhzdGGKdfLSSpCSC0k7uhQ1KkdqLBGVp+Yz90W74gOYpIn3a22FRLHZLBOyBTsMMkWfXIsrbh
z+WX9dPKW0rHn8IDN+A5VStBuzPpGLRpooPEHdMm4LT/lCiA2L8QkYRagvYWnUQtPZpi/qpNhEx3
f9v5izTunkZszz3OSO7p/bNgdpl+TsT3MzOlx0xNJyE7Sao2XMCroqQT1wPSOx2PaI24x1s5d5AF
uDaPl78h0qoKHQwAYe+CpqDvnQZi4SXOAEHDOMU50GT216JymMImvmZ9K/BPX4n7nAuTbNqn5lU9
bBhhcCgzw62DehGE7qeb5SyeDW/WYjyzQAUxvPMprow7LZ9hLjMbQvxJggZDfm4mh692QyaFKNk0
I+3D+Ow4z5sd9g+PXLsv4wN0/eVWsE8lsTKarBpM2RQGxTqH0xh979DDzG+C99+oIBr30VJ6hALp
Azo1zGUaSmHUaVVZHyX4ePcE5vo1nS8memqfB4azfdQBlQjRz/qhcQ/Nx2UuHrvhw9jMcaVyNEWS
dVZ2a3yZDSMKg/kPO+T7hjgLgYRQYWtWTcYjWStbylaQEX3CU82+Og+lnfH5epLVhYGqpv4+x34N
yABczDramL6M6OP0xvCACVQ1l9AYIt1iLOd5af61utgaHZiqWI/TKkNEwFpIjD2FfCYTypDi9ZFZ
1IYXLZB4kcDDWIMJK/oEjuh9aNOz08z9me2YhQTDiN9mAIcOWQkFuyzxU2vbjVJezm8u3Yfnq9Jy
SnoI/Q6q0GC/rUxBNQ2UkLGrFkrXbeA0MgVCIN/PxFy0ja910pEgnU0qokMWpzZ5R7QAb4L5VZhV
eyL1hJvoLe+9OHV3LD9O9haSg3/h9kmWzpznXkrLzzDUN0YoiLG0cSv5vPnu2WYt7CAtUEwX1wB0
u/kO5mxgzVs7uR/7npKgilmL6Km/nd2wzcjJ9V4CNsHo3NiaAQwHK8XQV2RoOnC3y9vH5qTZsu0A
cGDDJB2w4r1Ohxx0mk50cEBxOYr9tuyho7eL6BiK7UNG6kdBiSVvNP7CmQWl7rhi/S0v/uvYl8q9
LKCzGeL3lku44NBM2Plt7iPAhITeu6Vd10RyRjRj5TtkBghea4lh5IaczZYk+Eb6XADP0Hh2elvE
+rBHCl5tybPsX8YEzXIxtyiXTERVaf3A7GwnwEr2NELtZfn2WMTvv13johKuHnTMw/12RYKEdU0s
YK2SWUIcqOP5tT9z2qedIdVGO3KcA6moy4CzOZEkTC4DEXdYeSv+apGSEBtj2ke/M1tjsfCdUJgi
redQhF+mgeG9vk/cmT2hEAzIWLrsOpm5p9IBJrBiNPIaCwXAPiNta4prRBeYoO4YbvvsqtU3hGgf
i+rPSLitiVhhGMbDms0jNapozaOeUyFeNBJnbbQoq9ohpVRvABq1PtEe6yRjS+j62L21Ay3gja9r
1c8phczCc7oQkCk36NaM+atkil4Zsxxrh8GllKwg5hqNgoQthClqEqETUItRmmadSCxMulMQgqQ5
MpM4sCpAJd/ppTCV6x7sj0Xe5SB6BF1Kh9ucaf1cNwpBxbPFuLur32VeBjtV3vI5Zkb0BE1B/TjE
kKvzPhTPKiHeRtamswVYefOyhTIWqb3YMS/ugCJCbG3OKu+iNev5sOHF42/3fsIl65KO6xCD5bYv
segFXGAfb5h7Fblnk4Tph8Fsdc0n4SEEICSXziaIpMcxIeRSjqA2NR9fdXQ1Dxp9rpyYilVR7qkL
Cv1VnB2tu2E5iIR2xqB9ZIl6clJ9duDsSZX66ufBkQTCm1OKI8p6iBD13BxQbmfnckMIfOnB+7hb
oVsJguMy1cqwIwiCnAqZTe9gsxGTlXd1/IaOnCaswz84EBLrR9wMLzLGhcW6Itdir3qFu6nSLWJE
Jvza1LMdteZj9UAAgsGngTEiUD+ZPuAk2652bNwR4KuFnfbwQz4JxQ7OVVCLAYlyKzU+UYICVWTh
xL1NV01uTVSsp9rrDZPGBA/nhyg5fW0uorFx2rW6YYHsV4F41EzxVtW3FgLY2J4l1AS0bQV7F5Xl
u1pt8dzHNK0uUOrsE4a1GLF1ksOw2xU2u0Yc+1NxKiTiFmqL2WMak3pbMTIMYBsLsDepAvzHJRAI
f5e95Iep2JUcvr1tvk099y0g9gmtcOJeFM6TB9BB+TwwHY44Igl7/kuAMpp5hpV2381gw1s9c9pc
h/TuETJEjc4Oq46IXorvaqrkC9kFfieMNmcOkxBjtHt9wR7I3uF7d2QEo/UkSrJVXMgdYQxAgDaM
Dnl7Bdoxiqhy0SzIG5DL3vcXdoWz+87xH00cFGcntsCAjdoFwouLHrlwQOs1AlylV7lQcuAQBk/C
m9yjWZyZD8h7Zpvsey/1sVybMcr5U/GwWwhVOTvZe+CCc5SjEh60ObEkNwAoVkj5XGaKK5VqUr30
OLT7VVL7yIdTaUHDYqm+JfR3AZtk8ZfSR4DgX/VSJ0AxYAUQFXOjLFD/WWYUPhs+sgkltJyQxydq
TQBrX4CPBmX5Dg4GUAgtUHGTyuBLqUI8q6Rzs086FSzGDzq+/7djAu89GcIvtJbPl0nxUTBPg9Se
MHWoQBnWpgFa+OR2Cx33PQCBLjETnsnD7jvrwbhIrrLY2mlb1LB1VT9My6qxcCmRkKV1Ft5U1mLH
MlCzjIpRIiDt7NrsTA4SHtVkQ3i3H9ekLWpE3MqzYbivkmz1xAAAeUfMekGAK5rwF0FXXz1kdQYO
4mAAoKT0uhCE/PZVvspPJxgppppgoRHYwJ0gFoLDN1qM7m/i5Pn24bOhHupjm9kL1K006DUKzu4A
FmEsJGTvDKDbIJmV/T4x0RYpMW1MKNnKTdLbHWMnjGCpX28NiqdJylSltclanFg8E0DsBWHkNe1r
JQGXSVTsrbLQvo54/NnpBI/g0sCPJSMt9yNP+hH0zkCtwbMEcDXalqBbt1mVu581YXPVTn4u85N6
Wl9F31fQB32wXO6oW96NKjFP+acaUUDk/lpX1a5JnEqU6E3dX5aMjGMUt3//tqdY5nLlJwIoG5qm
1THCt4sV3zR4Es9XReXvF5elAvPewEEI1PQQj6E2+9c3QICP7YFVS4vTl7j9BYTFbD1611RvgBLB
vhZo/EK6SnETaj/jA05BgC3+dRIfJcSrz1sBV6InPXEtB3xoYxNh4HLpXCQ3TvVyI8YhOqzXcWCJ
oTion5hB3UKo3n9WNirnsLUFwWmVINve5r0FPKCgAV/VwW4hmhaVpj3mwxYV8jR5Xa6CfqMr4Yr1
PZuZHzG+fYzRj49saOeZj65miac7fxY7KZIrsCfNfd2oYH48lsu8S4FM1Qt2sI2hdrnnWqfsUHmk
z0iTKGYrVjwpqpZ7XkOliemCsG61ye5S78kv6fGNwxF1nwv+s4aY9I5G+gdv3uyj7G5L1TC1+6as
u3SUkxjXl/8PVgbNcAI9v1zsf0UOFLyts8N/hHfq7dwJq3W4bhfeMWYnpps67eGL3DKc0V3H9soq
o5wSB4RC1bGToeEUtlsBLL5LuFkzSClZV+Ttvzy2j5YSKwp78KCPTI7wZQYG1R9BV8+9UOPUtTtB
4xLJMttS4iPAcf0Fnh5FZm2/9RZ9MYe6n69SyUnYBRFjrA0Qt4MaF2fVWt7/qT5EaAppWuMNu7uT
0qZfybvsCHsNJQjoYGGcD1SIw47O6whXnlanQ20QrOCi/d7szlAFg9l2T0WoDjNdq0F6f8xrskvF
8uPdeqNwq0Q437Qbc9hT7d25aN9UDZCYNVAxto7+U9jTcpPIjDTw3d1CVE99xYw+h7MuXfYUAPS8
eZX6SLzdADQmWCqob1h2N1YqODgAA2Go83T9e8ivxqPBSvDNN6kPCEYwpNAGlK+e+MzvVTwS+Zut
hs3N3AnCv6ZmFM973bixL7PzI+20LEcicju6VvAHF/X5+SU3jspxw3kfKy750lczBMfm1gtIFnEz
qenCUF6THSYwJ9tZNdLQQ19lQpV3J66ersUWocZcEIt9Y418bIbIZp/NpkaZRKZM4hxeBmOPP7hT
jEJHbRvDDfe2m/hEFzes0DM76DNFsYIZC5VDsexC1tDPRW/9/rOgYBcBbdDCLxLmcCFjK3p7HR+l
3L6xiBJBkOV258mhGMNnNRyeQzJde9dsvn4viQpNxCxo/vc+CO0sd9kaUVsgFrCMyGYHPk9cXXg6
oaYGKJZsFWFK5oZv7+Z6j/TvbbLaeqVs7yj0TrbaCYB9Z1nOliYhr09yl74jxcex4TrMHqTgVXEJ
E371XmI/8+jz7K9s5cq12slnraxc5bTmldlt+BBH0AYOtkazvOoO5HwJYdx30hVaCoJ3mIR45CKS
enTou/HRFPfD3EFZdHt3sIn1qnSM0874m9oYPUxGMPFFdPhPcnTAnqBDsJRG98FXpcpnnDdLzvyx
dMVfFVaExkj2brc/bzloEMAEAOHazV6I+i7igIeT3bJQRev3tH2EcXw71WuRPul6gOjwlDafl007
rFF4eB2D95ksmDqna7UfBNnWWTWDMj5Qf5pAeWrmOFUMbvM7kq9Kh/mWPDiZt0LMQx6zBdXjPF3d
idCUEU/TAUBcsgVKiOYa1x7pQfPFWeAd30bhG6owhAvzCRdS8Y2iMVgor9uqaJrYwofOFCx1DxUr
xT15eKFhoGlWWKandZo88vmWinHqfp78pn4mMtIMSgwWaxqllt3fcB2u2jdpgrw2k8RJL3iu8dJY
m75QlH94IFZMrMv1e4RpQJVgfUcnpEr4qkv6Sx+eD4nfWnOcXlcsSPNw2nSarInGPwwFbV9TrnRR
JQMik0fCtqtrlqV6yzRkEQRBPaSL/Gn+qSjjNyeTrpDm5CxZt71ZAATrnUvupBEIhmT9Xy4TmKdA
eKEVGQRvRvqXOSJBQvDrIwaquQDtTCIk+Rm6KObGBpkUoaMq0VhzlvZp7HKIB+pwHQyYmp5So7yz
jlg6vbEY5qztyv4Cig4XjGrb2mI8StjXrXw1f++VgMo7e+zGXvPNgTBFlh59kMttT/yRPLy65gL4
rp6V14x1xUaXp4cVV42I3+ese+HgmlmW3TlVcPdGmsSAKJIb2RNeUnQUzDKsqeImQrkQpYBvjE2X
Z/OvWmcdk1pudxM1MTaNDUL13FfTS4M6iYV3VI21baQ8CMRYemFdyoemGgK82AtzDHBsvE1oo+B/
wW4440r0+LDAB74HFmVa6Cd9vnN3RyibUVfVzBvOo+3zhm28VK8T6eG1ICmZanwgAUEGxNFyEGwK
2vGRwP7ihBPVwZuR5Q8h6z+l3frakUSVYTwZqcfV1yBPW9rtbvKXEEspbWCOC1JvpUhktfbON+CP
WPLHREBSjLIGPhXNnrxynWyWPnsJwWH3vSMhPBsRYoMYRswdRBa4N1cfoIcKOeFDxCWitDBSc/Ks
Bhcx54gSLn/8GiAz/nzbaFjNGDyldHgj6MRoXXe1C13JCjmv9XTD6jYOvICJ8jA7+iElGFWds6zH
KbWznFc9UXmT3nnB9B4O9x2PwORZqKJ6S5nWbti3e0CGuygtBsBBoKv37zdFCZAUCDPvUhv8W0WN
kvWDd80eczTFaA+cDpDfvai0iREvnmNKGYEKCYkr7UguvDuVk7REHPiPPZf+4RJmCjx+xG2s7bmP
N2aK/nUauo4GpdlU7lQfy6SwpmfQ8VQe5Bk6m68o2h5l8DAG6bOz9jClOyrZXioHgLbaKGjxWPw+
ddKxxoN9Y0HnzsJJZbfE44VQ1YMuRPeAK5XhjO9lyYktSLG/00gyohYhTZkdAQj6UVWpBSrXeiMG
mAGlVUeKM7htZofL9/En3wgylyu8BY0YlXI6mEpIc6cMQUIUvbw8OjvA2wrJ9M+4qILy/Lz/xzFm
K7nzn/+k7/eBG0/a45rBtYjGQLayMih9Gjo+5f606vsCTNHmATOe4JPq92bHB/8E2jjY0KAoAbcq
ST/Uhq0xKlOjkMx0z3fd+fJZyDCkFFMfeuqx6WMxmTrWBOJPtvUDaZ7+9FNiwrgj0M4d2U3LqYFO
WLd0+qIdk6GlccDDDL8amQTsNJ+CIGR5fFU8sQ5mH2zLZLdbyhZjrs0pdsy1UfpYOGuMk/5xoXbk
sBmIy7jx4plX4ghokfDIL64QcoBV5a6SW62LywOOT1KGWNrJ3UMwak1/dYkaOKwKc0QdXCDrHjlh
QJtXTqef9wPUWB7sJ92m3e7lNbPOiUCev7XvUgmpRroMHN6FoVQlTM1F0nhYm8fddQDNrGFrOc9v
NemjtVmaDaLCaJwpe6eL5aIgxSoD8DdJh8+lwW9zZ8K+YQUBZWGs+YJCtTHqL5Mp43c7atZJwXPJ
pfMxoaSs4Er48+hSchCsOvyo9ZxXYTbZh18zxbOw2n63x4cww0oc/1M+FBj7mHs8OFpa1cSkIgtC
JX7jswauXZtotmjkJ0gzE/KmHgTdP6TYyh6qRv4zl9P6bekniJBT5WEuT07jJM3SN0Y0fVqS7Rw+
NT/0nmWLpxl27ALSh9OEg+qzWDZUZO1/4yONiZ3XwjVcAD/tPNiQ+npDwleJY1vX+swid7+Zz3DO
2IzHrA9ByhFP/e277wikllmG7TQ6CK7uMFmg7+JD5fJsi1s1oJOzAQG5Antkqg0flsu3RH+TORT4
4k949svyTF7qZmxKx/bSjRCwevprhWIfmQJt3BCV2g10CxxwamaRvynsHSPPBbKrnowkQjPmMhcq
oqgZ7abEkBN1j1ryA4cHjqZWaVWhhT3VfXw8J6sRvd6bTO9rzYlwFxx8ZW4ELGPt+RCnHbfmUcwo
PwB4y1B4WYHVdOAxv9Wiss6gPXNWZ3Mu78gHFsb+M2DNam0AKQl5jpbfl3iddkyIgcwEPp4WQJ0k
88ZvuP0Hs2XQQgAAvohPQK6JlYTsaUANuusey6ZjBd6tBMsKDJBmHN6W2sjrQMMUB63s6294yTpn
eVm2V2VKnNBm7RsWaRaddwU9nYmye/Zn66xq33rlBC8y03XmSf+Hbni1irWEAU/KnLAq3cTUM4GT
nbAnIbvpz2269OBNWFKoPXVI/Azhnts5DmJ5Ozv/To2SH2rBPzSbiI3R6Ge82BX8S7fCscyw0LJR
yVndVxejKmiktWDErylKUZ2aAI3nLDf9VVnlM3Bo5pYQnuDlwew0sUskl+t5hh5G7ofvwEG2UemG
0MplUkaYyrOxksNsPhmAQq5pRjYjIY7wKxRU2qImjaDmD+vCfVQJFtmrt0SMa0UmdvyEFSr0KaIt
cxyHX9bLy2REAnODMyHK4DTm9HMpjsXZSClKV8F/gjohRp6JM1QGCIBK5+/j1BnMW+Nut1ESHHw+
Vm04P/n3yoOZLyvri97QvPyKPuYG3ZBo+u9g6/k38/XuG9Af6KqjJDn1Z6PreyGceG/mV2vKasvX
3O1FCuzkJbqkxl0j/WHo21D6Nm1S5llmD1PkOoU29MOEvwo71t/A9x2y2iidL4eQubYOm5yHWJQQ
UM0+tbt3Kf5KXX1D2vF7C7zMGm4SSlQ6GHCT2BFr6V3FInWKMZeJiluzZSrLdI7fmIfG4u86DaEW
k5tvxuVucKaLJFg3f5gD7VTG+kqr+YfXiCoAoPnSQ66AAZg1v0S9FSE2UpkrvlgJMcTS/RGyUITI
tlR16HkdS+wpDjwe6uZaMcx2ehKYI4oExaWOHzQlYgWJ57P41GHRbP5sK1M0NNTolR6FHA6eEhke
JXDbFm9k4DDA3bc4ikuZmN7+diduf1/CqDh2FVc5QP1zKmG0CsWjN7M6MaIMHl5wp+a8qtAVD1tl
bdCaxtsPpRnzM9ieNLIGS4C+Jl4WLvkLZXh/4HgbJ8k/UdJ20abICeWuxRIDsnoZjoH2XZhakaWB
wmfNoUQZwU6dauDqdNVumDhWGuGfzuudjhckfujCD5l2S3o382MQV2UDYChW6U4XiJk1DjVo0rmA
jAEOjRxfW2Y984ba1oZAvccxq3RUhAVkwmSRgUdUiLsk3zwjz/wWf5wn0XCXuXftDFhuF6fFA0U/
8Q943QXMc21Ahy/ibbQtj+GqMBb+CLJaRbi/hngiQYgj+qqALVqBkIwxBpxGIszL8L+jcV9wrupY
SExEpzPMJEaBAtsvvt/86zR+Q/ojUNp7dlD1YrtUjqmGZdg4mMbTjL6zZ9DKthVKKb6kZZW1ZHvY
NuB59MCMyK0EKnXqtsilISTXhBIgctj2kcnor3Hh2KzqvVNhDfGnuVYqyblayRiu+0EwI5uBZO95
HImELZhEWL9l+o002OZtyoEjhRUkO4fgCkXYTaaVNi+nzRGq849S7MXHJ/fdJ4DHvs/JKgPB5ABc
YRrLhkMDPdvk/BERS/0TimqnAyrB+qbq3wc3RMzFXNCnB+K58+fGdnkhYXEoW4oBkbHxpyHmawKD
wgmptDpv/cAWk2l7khLprFEa/Kbw+AjL7w/xrxeN7mVB5+wTNFM5cAsQY08xB/Q563w/Dbl1FCR3
QD5m3dcVJbi6RCX5SSnvDfw6/q5IsFhYbSaU2k3YiPUCDOoMwq8y1afXgyWFfeEI5NXJgTGI0f8J
eoCrwBlpd9kk2iayvXOTmhb22kAchasHDym0jri6xTivy7G3Kx6EZPDKoR5swNp63p2Ii3k+1kqb
hjf7t/fmlUSg92iC44xdaLrfbvd8JJRKEo0i1wHuTwLC01neMQdcRSbx5CjlcFp5EX4A+2gcv5vu
xGm8155qNvUv8RIUr+xQLPfMCyXLE60rcCfYMQLYYCIo2Zfk0DoxvfKo8QVZmAaLgZvsyTcHLaLp
gy9YF6jRlXX0RoCg5NCVjYmH8S9BBXw/JDvZvzOLeJXkMC21DTkkZnIadSsXuR25PgRvo0QCpj4l
4zdR6c7LpgOgZhFtpl1/y2UN4dlhctHgcR21FvgqXCl47jfLzMy/jiWxO4f5TyPqjTbAEF6ELjNE
6R7pkfKrLngig07nvEhjd5jZaroMOhZaAkZUcLc5yEjhps3Ilas3uVhnxJevJ9RDknMyVeYhZTWq
G7AKv2uJfQnTK0zIFnOXbf7N0gnJRPAKAcpPw+xKHKo3lIxF7X4oAAvjkc79GrldvmpDdLsRubeZ
KvEPyqrlCYRrsDutPtj2eUqpvGNq4R1FixAPn78iho9rTKzL5oItwvCQ15mGhUVbhmp05FFMOT3p
UD3mvOtnvUzwi2NLwO7BTHf2OHfmixw3flaV1Esf1Syv84RnrzZGkVTuxrLhNbRnqapZpbzReAud
hzghhDOpgAdzTyCEkc071hAr0hpu5eu+wbiLEdt4THDqLupMc3CvMnYknaJb6xf6eR2mtES7xYJj
+sdKv5iDGxqCJBRgxVuCXxM4jOEhBs08aMgjCtHHQuJJl/cZRKk/xMMo6Seo1swsucUtDtP/ItMX
w+mzwc8wYUYfNSNA1318Izm/NvNZclrrWFnitOCubxWKMKo9rdJ6rZtrkvel+b3KzUEyVe2G1DFV
EHaKBq8lNDcQwZAO5gqC8PbnKjCgF0hS0iLe228kvYZL3br48l1rNfqfSMaZ66vsdaTRJJgTnOD5
3stn9HzjZ6kL4AmdLenA4ApHu6NqxUfgxy4MWFjG73QK56zDuD7ithqOP0Zor0qhiEkNIF56Sjpq
tyc3UbJhdFNDfm+xZ5awNBRplynpM/B0Y8e1xhQJf43UVKE1ZxSQGTI8eSXgBxFHoF7DN8bxucWA
ArIiEhIdb+DdWQwmd4K3UchyVGqHdMVg75yQYmxd78WTbSBt0S6tYm3gGJQB7BdEOkiavLK1bk/z
o3LAG5gn5dNJkRnrf5P6SjPcnTk7ezWNUwy0U18ko2ZYVsq/2B2mX63NA/zJC5+zy/lGojJPEpKZ
jJjEQ+GqQdHqXfN54HTcRm5T7k1D1ig4EvedBYYYrJDo2GTskByl+e24e/SfTULlVohX86Woc1+W
xRWwBDK8T1Apaz+P8jKcUkZ2Z94kUIOIs+xq4XlADR32L+jXTf6tc50q7FcOJn0E5BJpFrGFt5G8
p8le9Jg/Tx+qY8LMBoX3C/aCydsYkHHLO+2ldi3eYoyxL4A0hYWwuCbNzMz4wfaJjDY+gK2u+bSn
Jn+uYTqwOeiPvNjARgYK1NvZoE+3StZjfY+2INJF6tWlcP2xqlPRuH7liw8kP9VwNK3jwgzT2nzx
7Dy5WBEfiMbj35rTy7ILbVb8uWYRsD3xDMjNYe6PD+udJKFxE6PucXeAcWgOt5hLkudvbBb1uwC2
pirNEAUDu4sanmaWaupu0L8GPXArm/2u/Qo35YOpZ/n/Hq9Z+Q0vPuIjgtEbFl4s5KEvVcYxhvPH
x1r7PDOVBAZlnh7bxd+0vvMQhOqj84LaiyjnnqrNBIvnv4ZMNVHu3LVhzSKwK8zcnHDc2hI9+5Q9
3UZLMzAXPr16CQQInTDiWRUQObPm6Sq2zVW+d8MLfVLxVK7bQIGsO2bDrSi1xCb+6oC1ZgbmchLI
H+8G99MOUMEThA/ApjT5h90CS06fWSwOrxK+hu4I7glJWOepsuHKb51NMBHyS39enFF8wJ5ukY6n
wo5f56l4I/lHMUBb6Dz9yhER4rVOb0UcdXbJnASAE1ewIgyNnqonHbObWDimxqwHdD3UW+db1NLs
ezmbLDJ8nWYSPoDaDSfxIFF5WSDBTBtjhib0dhwVV+HRWpndUhpiTPZuKe0mbkIPrXU1fn5Y6UAP
sR2uzVKPMpohd1JNOtNcZZly9GdlFAAQ5fyKAQIniz7ZqWr/E1wwYRipYiePSc4V+Ce2wW/04V28
w00vT8lxx8V0lZOo4bIrZNY5bvHyOR1gs7vCQS2YFHyKibDhLWkw/czpOefrmDkt6DNSJm75qaI6
HOnI0yMps9C30zh8jIEQ3zOFuFHO7LjZ1yz6pnm5LZCZNz5RffTH1iQP1DMVNQcttTDHnngolcg0
F9gJ6ETa9FbVu3nwEhUtrqMcSYH1CtP6Xfq7Ef+zh5sprJcO6Avk12hnXeiYf5rScJp5nUhXBbas
DT1Bh9+m0fBiSKzaNVY3Iwk+BR4T0dnVLw+PeNg4QYb1BtNUBSuZzCP3gTGYBttYvglafb/L3oVV
eIwoSkzyx4qwo/KloUndpEiHZTQ5TImEjZwYrQlzsz4lXfZTduBE54cXTVUTCm7VG3Zinzx/3w1D
0C2SGv9Ml29AKsvsUNb+C4no+muqeBarL/218JFDRtrSJYJLR5psHioCw3zeLYnqjD+05cXWxSCU
olQotM1bxXDkCHw2PJnSTTMlpqHsZ15+E9hdsGGfCfo7BKlf5aDknh5Wybw7k4mGJ79IoqJ/Kmc3
bxf7oh7YRhA2cuenma6XXP90JQRWcFtHU+i2TgHVsNcXrJ/EtsB7E4W7SiHFz1tr5MpqSeVRhhkA
uu1IWXKj23L4BzlHcIacPI1L2wPKCnhFV6DmLPJRBZ/MnpJdikJq0RKqHgSUsWsYPa3eL+hbGnnU
hjwyf0IerrkcDZ+jvTZQeYgiC9FqWYBxEVYng3l0GjP4s1sGp+89TaEdoBv4NWeFUqSAupTGPNJK
a4EFFBMpSQNJhVNQX05PVJKxQx9NjJ/vQSsfBJGwX7OjZGddK99pcDURJD/EeXdW/E5sm4o/Ye6u
d8l1BXxOIO+ywfPiVwZ6R7CKZgN60QZQAVDeU+8FZzWsSHo6Vb1CWPMO/RsEq0azmsA1rfe8ssSI
0t4mbnMVD7F2ecbKpMp9j7lVq5vxpNgrluG4Qq9zKAkmJN1iowUc2WHEI2IB/bOep0+EFM1Eebld
YI2yRcU61thCSJVGwQd380rSugTE2X7CxlOJAEKaIvP8DXZ7h7XXyuw77dKul82r+WG0p0HEZQeO
JPfpe9fvagCXS2Z/ade86O7h7OzDdragB8RY/K1Ex9l//g/TokqR9hcRrnHtuTOpcZRbVNL+U44h
tPfUFy4KogdpP+Hv0ERE6PPRwVqzaftLzt1Mpznssox8EHQuyaix03uK1hwnrlg1C1QbfxME6oCo
2vo+DH6XMCD8za/rB0o7icHRTvfHlBW33SrpSN+Tnn/tbjVE53G9cmY19Piezp2njOoqXbg83BMv
YNQ5EcZBBp9c7bA0omtA8hDB9zkUEBerYYu/4bpxmx6ZmhpZMi5c0YcgUGfVPyMVb3ea2MoMt515
mTD7KwCRNrtRnMMf3GBcQOr85MDn+kJE4qJ1mNVpImNwZTu/+El7ikw1sxQWkUoK/9vyedSBz4fx
TpG1fxEHuk+JU7S4ttl87y3cfpGhu5mxTxydPhaYCRXLkldrobYm6J5EpYOzjMlm5RkwtquUa5No
vsxpU8JCXbgfMBAigzjunimSI+eGXk8WL6a6RHK6vqCs3QKs3PJijPadMr7V2h/4vPj6LmQtNY/q
IjJpRtY+kcof3h4Kpd55Q54kXQ7l0/tVn4Tq1JGUYjzHPEpiE+4AIhD/fQUr+020gFgtB0nNtc+v
poncvJoTowkgmSdO8yiamFHeWT5jkPMGoE9FBDcg7AJUJ+JyFzBg6T9shL7J4Itzzvf9FxrqaxPY
mlNMeQsWTxvtxbKrZxi8Mjwtx3zbhvv9Pk0f+aaOjskmp4dng8f8DqWJDHUue65gGHG9UkVbMGQT
M3pG7LWajje8P0LfGpeLRMKXi02a6/tGM0Se8HBZFJAnW2oxCx3iYWKu6NzZJyPKlglSRYeOXPNK
Y5ls5dp6ILixPrLCKqrykB//Eq4fnwV66q79bl3SY1hcN/heHDUIbV4wFg6apYhKi0XK6OAssk6A
nCYbgdY/ZJuHs+FLGsif6g8dkKX1+6/Ck2qFhbq8P+mnxdO5OFYjUASXIFtOhQf4KmsRAuh2bLvX
nBPqUfNZAQiRB3Jx0je9lINBGxTmII32YVIl2fEhn3OH8G3gLcAjlNaPQ0IvCcWKraqfjNYrr3ja
UHQZhnzEf+Rn16hno2lEopbUhVWlsPsHDQa8/SIF+4Rv+jXEQymUlKaR8Qp2ZfmZdRSWddtVEfwV
2K2WPwAVrpAbfTJCYuNNqeV94Ski83ZuDUGWGFY4xYeAJLbCS75RKykQVmj1MYdWFc4nq1syFqF7
v25veMu1Mol51zWU6Ho9EIFh8NJRTeJO8MpMA81NhgwqzNG5cPCPKHOue2qyvvcBAfJfved/aogE
KHVqH7TiMam2XqGfvBe5yDFp8i+TSX47oDU28NHaeQ3VYQPckEAkO9wd9kDTzy5STQIytdRXf5iJ
rAbjIn3amGQ3yNlsk3TZq1QRTPHwf6vPdQt6vG0NPB19wZxQXnautUh07de13JfrrhM98BNl7jv5
spNC28XrNJ3M/5ZQm+Cq791ZqBiNlF8ccTRjROGHVvb2RMnBG3FiNV5sOrjPAi5l4FsPiaq9YvBV
r6IH7cO6rblTRyw/hM7lDfaihlMgaPfIGS+bAkCoBij2MLXG1CBa5M5lBgGhwzNQwO6KAxFR7eDY
sUuiK8+GqV5u5AEqsjs+IyCUN19SbiaDzjLK8m7EZ8sNixbW6MoPXhTZxcIyvfZzeiCTu5m0K4RK
aDKhPBR3hxDdX7Uauo/swZ5HVidgQ0FdTsh169uLBD1ThZ0bCTQdtpBMcdh3IM8s3ohGdb1aVBco
dsiKJBwn2NDr9+S2kdAKk6wQbH/SXcx4L8WyvOsBVDf+266JcaSCC0bsuS4bmUUDPIrWaIoz6Oyk
ccxXUOp7AHvx7qewlFBswlD/hOE9GogWk9TVMN1DY9AaZf3Qx688AD1vodNLMn/DheBnzGdGQL/Y
CTG6VEkIoL8EyVB6srrXWmE3lM5ROwputP7Kawp+wWOL5SykLj3+wKX8KzHr1RKPEA9l34TSJVZC
TnRF4cChxVrBuNIRD9sQT7v2P8kVBAJs++BI5dwKA9z8vG78lcjx0o6N9bPvRv7moWkDUzmgXtp1
WTMmm/JnLi0IJ8D48DCLPc1anTTYNZsxmkK+qWNN/yBunReI3Qd29awqGxZ/OpJ7XlgdSN8wUawV
vSavo2WoCOK3EpcCIAuuWIoV9SsYXiOruCFUkJjdSXoXkkiJCI7JiHmfHvmGDQKvbEmfp1yeBOJr
mnPmzLsODfvXz+d4hq+SkGcB2SUgnFvXBHfLP4krInMqWDy84AvFRMcym6wO945WEMOlSLU0TY5y
phswpyb+L5DNd7vcOx4lPimTHD64FtxuX8xXLGPHG4xVfY8DMwp0EtwZ9EzXNEKWp+Kt8bEmAZqC
4kX9mh3sZNic6PPzLwLNAncixbDAHMDvDtq1HUY98B7YMZ163PcpxMLbWpgziB93qtIlWOtChFyZ
KJaeR7E0JbU7qQk31Yj2jhHgTQmSfvYVN+NqzNFIf63+vh8APzeLz6jSC+2CK7HqN/HS0S7zvMZr
857+P3NeqZGSHLKmrs2u9IMCubkZy2liw9bDppXbAEkBdHcCeQkX+gohuR7gW2nOJBRJ+yTIccz3
C2xNm8i8vJ3EYQHOMuJvF6UNJP4IW3rmqsbSuCeRj/WEALWNB+UdeCdNT77Hbia33l5JVcXmNT5/
rby/H250c6qD3xZhIY81mUznZc7zNzKCTODK1QETn9ttBG/RuSKiEQ4/JBpHWiSVgEkQ+ADcTpsJ
QmrQR7GoYpFi6ruJO6s2aYkFUEzHOYTggmJ0jE3UvOCIgLAMQlylDW0VvgcOAkQ7TvQC4uJlD5+e
LhQ0fdCtOVvMqaPEqViDpRVL5nihm35V1OLeU3cMBCEd7NZvMq8t5xwZ6yVDkB9MIATSpyn1lK18
Gype2JVV+YEKFzU8MESn+q5v/c2LYvyoGgEt7FUJKWU4ivYwm95iRVkQzmz/4Aj3uocBQKB3ELky
WBW5s/FwCLEfOVO4zqpC+/j0Qju8wg+Xbk+a24SKO0yRci/adwuKkYEdazP5V5+ypEf3FexkR3he
BoNhwnffCtwtDgF0uvpa+h+L0y+IJuPMtvizp15YGw81ONyg278gwXlzjYjWQ6Jlk+vGydzbEVbt
6PJdMcd+BA+SAL2OuL2Ki4jaaMdN+3iW1mkL84Vs0uF2jTsnxZolHgGWFAEKgHSFjEadYxaOzdXj
jcY9WWm5rUzNka2HjPX4hRHU3Xjk3nFNFpzyhzGqdfY0Gv7qX2utfe7IFrW2wmlcFIHlxP+so37K
LTjO7fYlbPnBv+RZjYcvOj2NlzAvjZhm+pCLbWpG6Hy0QWE/EbqW5sRlt5gZE2LAWRrsAm33fTeK
mbhhnEDSxGtJBR46N3op8oclmHce8Nl7kmH/hRQku8xpPU0jm/33Ds8iVYAabEgDLclgsY+HZyba
RQG+qO870/q7hjbq/KqMQPfK4fGXHjWdzloX/KrkOF6egnghYHLreUZmMK6wmU2ncV51M7V4d/tW
bNPWDm0TK7adDtsvykZ6yRp1akUiwgfLwZan3Z2ebMCZhN43dUyA8t7ZY1Bm1BsE5vI9sEVrTXns
gDsA7Kf7dBZ/19NXbNyAzNbxrct76o54eIvSAx4YkUnEekj+2Jizgvf4Hw2Bkopsk0MXMiHOr/qo
Zm3+TVJ9aQHdGpyRImiM0wjMChtZXfKSgkE+VmdrFLC0dXde5M1oZ5+jyw7YYY8zUiFmxi4bWafi
hr4ySXBoqZpYPlC9+DLi7DJgYnSMkEqESHcv3CgBxQP7LrmLe0YpvkZHvvCUe/LeyjY1atXUAxPp
hYCY0oQbV6nmlq8L5z7R645yFU36ixdoz+AMypbUF1uBCqLKEw6Ten8+p1PacpritMtzgOiSvBhq
JvX2mr36HLG7zCdlzpV8g9NTVYmnuUg23qbdMPfsurhgceBes5A79tBYGH6ncsZAgnWvkuQvpPKH
CrHRY2t0xqPd5BEa2yEhmIBXdV0aiIJmmIzEaMnGLejTOFXpIn4jsHs8h1ty7CR9/+anvJypXUHK
6XOQ1IFuOLXq2XX9QuCrG6kjRIuQoMTLo2/Lir0QorrLqIzIKr9Mh/IqUb9pMH0A9jmi1mMP+37+
LQD+A3V6MSkxXZAUlArunVLtQXtT3cGeoHCit6yHr8ctQB/D0sS9LJaiEB67HeGUByBr1hAlbLM/
CLbztVJzQNW0TRdSw14m0Ckuq7DPo7vpls8pqUBSE3Jwd76ZbMlAaB/LSPxBvTVE5wauQXjuIqfJ
zy/jikDL7HVy7m8u9idOtvZpo0mB+YPyZCoM2NXivyy+3j56jMyJr+EjQY4duuESM3wDKtPnfYJp
shnErW8Ms4R7o+/48s16O+m5TQbFOzulKegeWgz3PYsps9uAccJbvz1iGycOy8iW2++zmc/66Plu
dojKssxaPtzvi00J7CSMmCYBlxnLMuxtwBpuqFQv4psaR2W9BmKaoJ//FaJGnEvmuaqVQKj6OwIC
T9u+eU/3ZdWJLKv23LMN36LTAlpzP+m/iXxivZWdNqx/i4/R6Vpnmy92YmyHBjSSHE4/5le+7sWo
x3fT9T7WEaSQX1yQtcAYAbH2Pe3dpmHvNkHza72pyGwxk6r/6qi91UKKju2Kujb9RX4Oz+C5OXgY
I9PMMEpAG/ZKUjkrYDnGU14AQsVjbANibBXJGemM242yeO8/NCW5Y7Bux/diRSaXjpsQm0llZdT1
sUUCZ6tQMIE+OHvcjyygw1TZwEmxcckygXGC/AmjVb2CmCZj//C/l/fTPlVIdzlNURO0xRY2O6OT
QJ3CfDgi61guaFLklYjMrKduSeNnG2m5gELMVqUVQh9b/sh1T8Eyqa+NxH4KL7lEb8oKj0nmqiX5
zWWESlNmrhk9ilrmjDtZmkYeE+bhlI6VVKSon8TvRwOLSnu6snqp50bV0ThOHcvrxXO/2QpYE1Sa
HclW8G+wbePMCgDqg9hZ+I5NdmXVgYDY/c5XC/QcFJRJAOy1J5850/1T7bIZXhLpmtrkU8Y8jeqS
KV9C+FvRoyQzQqT3nn1rjwQGSeiITFg/Y+YVgfXIQ6HYv9MmyitEeYm+EOaFQsH6zhViROdkQ5fO
6/WEbONoSrtRRnCuvZQ82JlQVerB71Ox2GPiFnl10pCIfLxMiiWNo/IR9L4V0pZpIQNN4Qauf+Rm
8AdkbEk3zdieTrm7r6aBuuVx8tRR+lOHQJuWloFCzYIs2v468CeWpDKROSmfskNXq3uSOSPLWauY
XFcWSlcWQUH+iVo82PZddH9H+8Hb0GNUFNKCIeDE84yRcUPmgIbKGPjMXklOEpCCNsbXdg8CV6sj
P/Da1lqdnGLpDUzkk1zirYvBBVAsWpMurX6ScnTomPndaDljjJ/ZJKfSKSYYC6OptVz4KLUR3h+1
N8hpHXRgeWZFR49FdH/ktDKEdx0rXYXNImyZmENbCEf+To+ECHYrsipFLeJJtLNpbH8HFK7in9ar
uHwhicKA8gKlmljQQqPwkVsf4+Qh2IUyBhxDAU+MF0Q/qIbmMZ9JMn+DcImwp2jjjiE+oAqYheDm
5j9sDXrqln0WfxekwZSQVwjgJpQMnANI3oU+lg2dh+Pz8v4OqCOS4k7LPrmEBjyeJFI7DDX1Mitd
W8eHtP/P9VJgYBqsqRWAEFJO3LHfgQc/zA4antje44ycQdDZBt0arqrVOpAh1TlNqHcn0om0C4kk
OcKvhjRHE6cPEZlo1DZOHMgtOzbcmpw4tOsAhJeQZRHG4IT+rEE3eP3wkY88sXmYHtEis0mlMv2y
fEpmuv27h6s1BBYAGV6DTMTw4vj6v/u1Umw2NSkCfSCRNtwEOK48BDYysXBtZhZE3gLoBt/UHnTo
XXvuDGYxd7H4Gw5GijZAF9JGKXvsm17OZD2ugwQGofB7DxwJTN4/DtmL2RMlGTM4w8eLEfvZc7Ir
NW3cDTwhglt3sqedechtxy+YY8O5ibj6kwzV34NDSHw0Fb4FQH+7PpIBpuC58AfeMspOJI9hUlY5
T1d/FCj5rv3+/cuZGn6sM7wyA8yyBUP4Gqp0Lzs20cFMCf6gN9/Bg9cvElM6STSTR3Z8EzTSo2E/
rpPERDq6b2x1QnYYdOihRx7vZdVOF8EqaizqnVbQDfWmwuYwDKsXoeXhSNdHViBm6Zw/+tdyH/BS
oPx19ZuXVJJMVc4f8PDTLvMPdYy7Vm4Gtv00F5d/3aXx83yypTpeRvmHylpUBrzzx9X1xALWnpLB
saj4hFJXbf9At6kIQU/XOPBzUlGIRLFA+upX+/MdGODiREGOoHF719Opj3c5jpWHVNV6jVYjXa21
b0FkOPNwXfR2MphQlZhxPIhLb9sPk6Na4/6+OPJI228TH8nzWUzHBx3bGLja5e2zPqpMVPPO7uSk
lplUa2rnY6GKw5Ix0mBgLlH9fxibT8iNzF3Q+mvDSqCQEx9rplrDgHaZ/evAuQY0TBRx1psuE/rf
6o+t7tCrNVIuKliORZRuduCbnTcdVvihar4FP584Jhm/HpbT9I++9VcTt1DEZt1Ce9YYhCpZuK0t
K9zCNzmU4HgMKNlBspbw5IIzoE0L2ZbMs3XoyBY3gT1RHm91c7umZXik/A8NxSLPQRDAofwHMZsC
1/UzUUtENaXvQ29Fu/UEQk+F3FpiOeMeRMD50w0LyKN+AposJW2/m8jPslw3DKS9HHmMerFWPgsf
UZIm6j2O4qVvrISnfmEUSHqGE2mUYPc/ugHTJZyNQQx1zGakljBiV4Z6YUbQUVIQExE/OWeN/9VF
znwPFhM8iJnP26JSAy7r4EIAls3GVQwZb/9CHb+ToTAF6fLykBgw14mpVOy7KUFulxl2TYtLA5YQ
S54b5RTo1WfxQpceTwjkeDznAuQ41YcgxV8nUe/QYK0Qz9KGJeH53YXmJ/mE9pr+CjW9fnhrOW+r
xFYK5sz+DZjUOtCgByRKI7i9DaA6LRw69PVOyhayM8WNDmYcwdMCmdULF0BxPt7OwdG1uWTiGj9S
eiyNuAO3AptPPKfRwzX6UTlOX0scRy9HyL7AJnnSHj8UM03tJuo167idCHt6ptZEydWEAr0MXtIg
yuiJgrCTO4D8aozAKLiIREDg6i8Bqp/Ho0GPlg1afXUyqnIxO6Tu3GUB5WMkPwONBfk3iEFVddAk
j2J8sqxrhG1uX95rT5KIgqaA1OMNFKT+FjGjI2t7Fq56N6pe8SVszrKHVBCmFTjbNT3Q0boy/5G6
f+LGQxiOe9M19a2TycE/2UnheUtnSbEzyl8V16jV4TgoadD8WtMwrFta2yg8mMccZyQQi6FxGoXA
SDWvMzdyzo6zng47enR+4yH3rUXtHZklJmTXKRqdPS5/wNd77tqVDh6Ab2Vr0QJSjUtASjTDdciv
tB+S6Za2A1OHwlhZYzjEtP8EB82s0WO0ImaKzPNYMMc5sAmwk83K5+Spnvum6JU8Pn2co5y/W3og
u57JA0ye90CgUtve80r6IqO9eRwKOOUXCZMfRFMmPmXSLvS6OC6qxUt0G4LSIranRrLfJJXVM6Af
kClFsbSJoxIztj1moUfZOwLttVblcv92vq0JxviqwlomkTKoMHaWpoHgrfIJU9FXK+qAWsleSd25
NofxctbF+yiGjawoGqaY3r0sA4ph3TJBq1dXSOl2dnJxObCFAfPGLuORXJX58YJps8UXtafAkFqp
KvocpcjsS+MaLL3g7MpvrqoNQSFwNBFM9ZMK+lP50G2HCaBSJ3FO8YSoFXl9BiCLjm3SfB6CCVvS
RZcsMFiLFJaE+3kdpz8mfWGdUJ+uH4VGk/SM8zpVLe+zBf79bTF3jsWJuFQU2IShwfRM+cguS082
j5HlimtrqKo6X6VqLZQZyrWX9Rqnlv8THUvOs395Iv3tG5BVrluWA5KKwHHMTmY1MKeoiCQ18PCT
6B8PSvtm/eKbtYZwFgKETakf9Yn3bSqbAKwKJvSJEo6utUmpXEdc4xA7QQIrlh5D8sGIaKpNH6so
fSSFBDCUfCRTVzIW2gbF5esOSMp+O+MM4Ht5sceixk49Lv74shdBxWHBiqPj1QrsL9T2BT+tSsPk
Ok0+yGc3bHfC4OmY1aWlHNj4plI0v3beZbPh0vv6uv0avYEO26oIgktDSlfvcE227JYsbqOslEeS
EBB1YWfq4SY1oXtFLHFFNW5Ajt95yT0x1gCwWlHqSY0Pxvz/4X2lGJ+gjBYVGNSJdxBWU+e4rq9b
aLUeiy1pT4F10xBY31lqhcBVnWe1nsN5B39xWIvbrcSlJ+Jd/BTPHJUAks2Kj+GKaCtJCoP8e+Yk
T/stHupIpCxWl+mN4+z7qfF5vjowh3+2AARZ7JJ0rWpBR27ETQ/nEZa9Xwx+yhdkkMjGs7nBY6nE
OFx9kh7Ss4iqk1NoGNXx1HDbR2ALkEX9eFyQv9dNx5XBw6kFQtnV4YAv0Trx75dpZmp1+JeBL5cS
WAw5Nd1u0HrIFz/1l1kJUdxdEPZjcPcFM2xafzIfZ3V+tgz1ytzSQ9/gjOxS9KY7+IGpJsKHAklK
ez8LMXVq2dzKmDHqKchUCkurdglAJEt5BdocXthojrGLn8N47409FNcGFigw+tKZzoFpiTm8uXCG
dq+6eKD0G3IKYIlfsmMCmQ1KrT4KTC734HEXuaMIb5fLABn0P5LCbSUpZeZm5/xRxUN64+47IBZP
7n6gzUjRy2uNZpk7r/nz3J1weDIGAwTKmvccz8tLxijPu6IQ72as+OLnHFoQMT1Xd/3w9Kd71GZy
Cc40DkoD41/DDmDllt/QtImQ5o/xK5SAJqbjAby4D2vQQ9henIfI5wh7iTDD//m3V1r5shE4cZNc
sQP++Pnad+qOe4MOFceIatQDNX0Mv9maRnaABApij4R5WisGXt1KYE0M1v0EQjWiM6hxjag4P8i2
stNRbNpSLA2TAwWEjrMpupP44X6MuNnlMXXbIQkqwI8xx3yDfSm+CLHjehxafMOzEdLjA5xhYikI
wgKqdxO7ObObLpaVDDGlOYGn4sHb+4LS5VTa8OyiJxNkb70j+EqVJsOq7HkybqSpqXSmjRQpv43Q
w9fMMsqpH0B1cIdgEPAxA3ZW6FOAOMfg41e2+PJ0TU9sTFNyLd2XeN+z8PODA2z0MHfdjFm6fb1/
0i8nf76rAZjk6fy5yksdFytRmUPs8OMIDk0QZ3RN7URpuvNGk4M91yGWjdU9lby8FzWJ2Oa+b+Rw
2L1IzniLq4r2rzmAAdWXFYFzmU7K9reQccAeXN3Yam/7Bffmr9j86LE5YwXToTSBNxW9WI9OqrxC
AgU72TAMLwkLj2ajo6202MAfqyWDgn4pxQKQlmj5KUO1qwsSMZv2+9RFFR1Qko/EEz/JITWH9fQn
ItEHr2qMr6laxElEP4lh5dNs7vm16r2RGGMqcKLr7QZg3fmVWskhpKwjowVqSzEPIM3DmnYlda98
K7ZflXWdQzLfNOP38IhOUJMXELnWpDvvfCElJXYQUYLzy7YwiYbnSM643j030mMAD0zcI3opCKFs
ubc9zmRVNiZKivtRCplV3ukn+f1t2WT2g9jsxtS1fnwnWYhlL7zst22+ale38sQuFNpNV40wr1tv
lymaKSIkqb1sf3CcTIeoJdV8kD/dyZYYcf5O65IXUO05pmKec1TWyIAet9PQjxWc3ciuTIi0Z2LR
nvUD6dRNtT9eiWlI7KxD/acsuXA1cM8+/32c6puMsRI1JOMQNAb//aDtokR7+skIJguSeDiSMu9Y
JuBw2JzgtSC9q4fiBdHOat9dTVX/qElznqccvxykilscNOPGQVFKzsMKJefQ+I+FPi7x4nPOwRLo
Ydh7NCHpF3ackgFfzbKFaAi3vgtPdrYMT3bDfviQU4869XEonPQjNee82EqCFcqDdx5ZMPaEuTSM
4TKz7HoD7Ci64zLMD6nbkgII0OntoxC4W2DhWRxolJKZ3vLzVonZJFDuEltVj5gKQcJzipr4cYL7
Wln0/HplMwcoeRhNPU/5KlV0ibjk7z/kWtAFQyYw85psYIN+TcS/OOoKE/rapTttshrWHLhRDMrX
VVNKSWs/At80E994f/Mi9JtDg7xjPWZmH3NfyQIy0Wvqq4l5XrTKzYCFQERKyaJtOic8n0bLDe9j
k2en6NN2wTOrBxFZRCXAFaRqc+bkmNflH+2wq1DwV6Ccp5Hjj9naDNuEPkgzpaNRFqttt7oeFmmY
lxGKEdm69SUFaCHFvMLUEMQRFY8fbbKCjZVIvuMU6TXlhbbjP8QfdcHrF4HUh38iY+yZcgiXjsG+
CLoGKTRMZH8MSEvoepgouBLVRAWKekQUOsJ26Ci2XsUxHT3A6njGPeTGvQ6JiZ9cQRH0BQByZ0++
Tr0tTyQmiVJ1Kf+UcLVJEfUt+mZmN3VIJD01rAzVpASm904Z+5EEAl3701kUX2SJwHG8RRvvT2Sa
pDYdipmG0LaxX5InCFb6V+JljPP2DlyayrswwkGnE4zory0QutcSLN4q82Ao4H7/jGnfuw2h1kSR
E6WL05VK8JeB1PsYAfNOaXJW3YldNZ8AGIBYcw470i72cex2u6inIPGNcByR4a+U4zrf6oHu8yb6
2aYl/wmvcAZf3yU4ZzrmnWleGSPBBdU25h4YdlFBfn3rX/RTQ/9cJUEnB+86YPeKcdECInNC4RZ2
35/5h/N50Yw9QultX/JzPsUFx1Rjl20Jqq0K3rzWcH80B6r85sirUSIYMDUxr3Hal7OOyEyfw2so
wqBE/suOvEyCuuQm6iyCcKmETQ7ncO/g8NdRZcgE/goULTGZiEVYujU0wgzdmmff7AupXTL34QDy
a0jyy89yieEu10K63pypoelMxHWIslLDml887Kqte+HXqo6A3okM+QUb5A+OFvwP0DVS1ZX3RG67
mgWDEkJ27Db5fBlkKZ7BuMS17rtKiVrx7YxYrpicmNe9bZ9vQe4zEPHr9B2R5dvhfZ/0CrPNLFVK
S03c/T9jK9G45zJPPF1XRjgIp/mAbzsUuxT2x7GQarf89en+rSqfm/E7lH4WtZ2jBbmrALTm4wjR
Y3s7JBMKLVwEhIwoRLLbxywLF03xwAdhykotowxPVnPYAccw3Fp5T77J8PCuaPcQ4GfsG6pFVnXc
/UFDFoJ70OpAPm+3fREQeZnz9iaEDyjVfpTJ+q2o1kCLNvv5nD7wwX1dK3jL17am5gB78fBsZ4Cs
024PFSl9MLy1fVNFG38MGKncTgiykQGb1vJNGm+UviuTZKaVCArrh79z/BgoX7jcllAthgrf7tpt
H1wasPzyM5eH5dKVqxOKj9yFE0NZiPy2NvsZykl/g866n0GQBcpJKvCqJUC3oLCHD4KD9vNvzYiI
pVW2Dah3Rdm/+ay3YrKPMkPmR0nWICYYDPGfijpXJmEjWbSJexTmuMDQt11Uhc/4chIQFl/QIOUI
AWv574LwHt8FePx71Xy+Z97L9u1Q+8Fv4TfsNFyfwzdh0630TprgrrIyVLeFVnBhwlF1UA9D4pm6
cSO5B3QXBpwGrp+NKIl5kKFw8zk49SnW/Z2U3VqLHiA+Xnl8i7V14WWY0We77MPOug/+a2EAgqba
+sO3QczZueMe1NfJUkDV884FmV76VfGtbg+t3sMUClaRlXeVgOVodtr/qtAGK9HytHLwrhYGyFmC
mQ75+7E6xVuBHqXa6Hjb0vy+gctbf8ltBUO6wv8oNlbHD4/gdwCtxPrvNowMMCukvxxwDG8ksWZv
8reVEAUDRbarbgDRKnHqEG0BENIHI0imIzx5o8BJLqbg2CH+j8BlwKGELo7yzsdgYvYB4VHAf/F3
QHaS/YRrMh+arwTWzcDS9ufN4tWkMk2MOKB2qUHHdWh5I6Nc40B/Ih1g1TKYWjuzbEXtE7XapJ8v
sRIV2d7joIhcLkpO5MhqUd0wUC/lexf4Ix765W616cJF15Odywyx7LDC658Q38MG+UMiztZfOGwx
xjkCSjYlvGBPUxE890Y+g2j/uSa6Le0YHDDXAehEIklqxbpVxYWpH6fFannY1b49swVbgc8UpoeS
r3oIynzwNirenKLYOi95LwsSDzC8Bfe6WBcZ5GSU5EkBu0g4yl/P2WAolxl4XB7rdL85wKNI7yCo
EJU5Y5uInraW2UURTfrsywvCrlOJpix+ewNrpV16HdYmyFcKubhsoszjmD6gz+AsYIZupMxXp586
P7cvvgY3EQaDaXWRCyz2dKvfpuypkZ2a5bDBzADphk2pheHJIHLfdDMU8RVkqc1aOF8TerEuqKbl
sBZ8ohUOqxlHlx7Ii4JvbUi+iBuMEKQu35FNTNIl/LT0J4nMlVimp5FAYWBcBb88ZXBcblyFRMyy
1qMusKu81qpAxYrgA2RfS6zkHzstyZR76xzS/FR8ZcnXQKJv8GyCoK5GmVxlbfakmHBTXnA8gaZ9
pM0ItEoiVm/0ob+pyWBKfD5HOnOqnNHghxc6RdPMjR6e6hXaimCFqIhhudLKQnL2SFqHUvKmbOYi
6/D80y9pG4gCVrhaPSE6omm9L17Dzv7jUi5EhVJKiBr/aj8xob8/YeirixEHrx/ceuolKOGQ/Uof
Yvy2h3zH8LyhgTKgPKPVSjJFz+fSO8DCYD9xyvrHx3h4Wt4lQmkBe88igoJFmZLhyOa5ZuGGCrCp
x1sZG7XP7WINem8QcI3F7fIUQbqVMHY4l0/NNzf29GH9gcyUhXXcbl22gpqbm8vxYzNYqoXjrxNU
oO2PXO5/I/n7y2T9v57mTSQ7rFOGhSdGz/PHWhFx6LYhWMvCgnIbgn2c+hIWXU8tOzqsm4cFssbh
p4YXLXJf+h03StNVroZmktY1XQ82TkqfS6KhCtb6sDN6ioH90AGpE/5Qki6PxZSH5zdspRd12EHu
MoNs42DY7jjt10GmTJL0amh5l5+/N/FxkvMD9mIXCDv2Jaj/+lfjgTNzzZ6ukic73c8Ur+Auuxz/
yCEMJIBLFj5Sy0WK81V3VMHihHWnZJL0V+v9riONVrdxlOtfiXEwyAmwDt0hKxl+93rxMR8WQlBu
XaHNV8/lfIS0JDEgEzigzcx5temd3KbmhyvbovSFdAffBUdU1Z+A17i1WKmNyuDU3NAyFF65pX67
iSJwZOzLJTfXenzhRgjQRpTObn9TfXqHJHkrHRjHhRBFw+kM50J8Y4Zl3lGrRTOb4RPSfL6QGTbM
nsnNMAQAI9HFANMmRt6ON5zjK15+Qc8w23grhHMPLjKQnemHY1S/FbPyk73QJmK/5EGyWoH5SMXA
rVkiIhpHqdjyPdSFd3EnlOCFIKVwwWxCGCXlPKzzpEuqXJ1QJS0DJJRPuj72vpAJuZ0NN4KRmPfX
HC1ckLFkOJQbXhFPwJE/abKsfBGfHQoA0pzuhjnbinpB6llTl/ptqFfIrceqCA8yGRo16cMArP3W
GaNBB/1SmaiAPS9n0ZUq8gm8kyJxW9tVgiS12WZlhRWeV1prIimVAJcSonaz2Zs85APTtW/BdW6k
IL5LIIWhs/vIz18VyvVkU88vlSMUr1Zgz4kCtL59xdkpmh3YApyM7RyemHUDBZX63S+vzFjVjeZ5
7+4TeHF8RvMW0hdynuvS560/uP6LJfDuU9Kp1ey6uoSVF4heIScB7xRMA+w3EaHyzhOZ9bcwSdKW
zMeBjEJpxJuOpfxWDiFGoUEM2LvikSDFcpJjaNFhEH/qsootNak/h9suqN+T2OaVMZpV7V0Ky6iR
hUCAEwk6BM2F4oWvkjoTUkRgl/TDl/2TsArK/Q+vavGx2xBCXwJ4KKm795xB6wvtMRBI9fWhBZuJ
ubc/UwPp4wzIdGb/1Bfysnkx+/PPprg8DBrca6R9aUCFUVef+enP2zwrI5EFaDdm9+pQMbYk8KmZ
zhIncimOtThd6qhWjRTwCzC7Obp2OToiFp7Y8vCM4XB/zWqweluSCnnbNF2GKnmqawrPyUnJR3oP
9+SKvLv0ISlp5o+AMYN5jENFsgZWVpNTMfFL8KLvMzGLyqAHJ6XXU28lWSP0FD81GuPB63cBKN5m
t1avF5FbL+33kLRTNmAu0nGhpIN2KWpaWGm8RcXCXnVn5Fv64aOXFik1FYdc9FW416Gytb74+DoB
AtjfsSrHp5cDYlf6HFF3lm3oJltLH6hlLf21CkUetecRR0je80NscZXIO62OxQdtywRMSTKGko07
fhGhn9hC+4snkiPZ9Xh/ZVxS7d/PsbQQ8O6mcHEt1hAZhi5uWPjF5BUWOk2NrWShqwahzulPOpC5
rpIEWPCrmA36aCvnZ2QONwB/iqzFWPbeVuQmq2yEVy9LuAiQkCF5ID5f4g75rthRD3aVDnb9BGcY
IxyBNbHgO9e+iNqjvh3zRj0W4mC+MZpxovfXTv4SLbrCduY7BVJOoAPGayBLzVQzIZu8XBpP/B9i
ZSQcOiRZQxbADYbyL8nXmxZ6KwY8n4HpbeFODT+tdjsPNJZUfYsSQ+I/OW/24X1SKpzdv8cFSjFi
2AQoEBrOLi28/7vyNqf9j448vnIdN6jd9JDnV6/QTc/5REgJlpK4w2jt7jw+ML7Ueb5IuihacAYR
9QsFWGkqSPlLIBJyBcBontWSU5kHTgjWUOWToEACyK343+Ci9RNej9VgemQYwTh7QDgwKkP8iQMV
sNQz+oF7O8lSJQ0wlyQ0ti8/QTKTSPK8y9TNrt0cvZ+32q1ShPL2oH71ixequutGN6/MPTk2Q7Zr
VgOufmFbtkUvCcM5oemX4kY1Nixd+IT7kmNXr5k2DDnvdNgfi5O0KL8gIsLM+rsSpDncumIOFT+h
r47pZRKy4QXOEWH6Y6QflCQhvYBpiRsaHt1HUAd1SO1YMmwgTgLK/fdgYn7rfynaPWRtZwJuIG6D
4cpB1I2YpJ8jiQSSHo9wH0TKRtru1aIDP+P/VDLlUcHfFkxXLmdSu5jDeS+NWaFLuuClrn1ZD10k
EZLhHbm8JimMMcn6ICpbOGRjmadblPJstKphbynoZ+p7aGxZen9+VZm89qxUIgL9spLAPbRutvcV
6zvLJ0h9SOVWGKbjcdbMhO/Ie+g9rPDKZRG1HjTX0bf9esrLxdximZX37hsa+o6zI1/YFxNmNq02
izhwujfXetNLbMGeSqASO6d+OYFdQ/UxaqmlO2541H+9pcYqqKuEU53bUh20iQmTC5G6HPk34EdU
ZwH9gBcRzcMlH33B3JHs4RdZpPm6TlbRe54nZdIm1EkDh0QEU2sDJY263tdEsHNsNv9lhuYcpjJp
8U6JOBwvDNVp+rwZ2yEpRA77ULVZoLhGGKHejNWPWgpxrV7CIY9huBZzRKT8WwyaNx4gsmFU19rC
UWI9JlyLoftX1wROu5UTz9J1+m6GPSKw9ANBd4XXAYD3JoWR/fr0HD/m31GhpgerihA0pupYe8aC
xDam50kij1sv7ZrYN1FcBliysDSVFsWLSd4We6yKBv4M5oM4tdsrR/7a4KwWVe/UaGQWKNDRS7Mw
0MKkSKEAN7DvgmvaYnZiN6goXNbDHTgHaUV3Ova1lyvKf+4K7AdB1+7ERyr3wol06ZsuCYfBxfxr
GkouQfokTMbGEAfnfAhXajjNZP9TPtvT1hpHwpmup+LhBmdt3qwKydAAIvLGnwJ5c4TQ5RYxzjj8
nCsbw78ayiK/Mz7vc1GVSOc24z04iGeqZGXVjhP76UZtq1FHqRpkyvbmy2DMvK1N7u/S89ulD/K8
uXKGdG5mqIGjfNhYvfqjwkBMmBxbjrMKdZ3WGOhjlRZaZ0BEyt2Zhm6UUpaK+aMqYuLff0x5aMPk
lUU7aJpZXtmWG2CKmbL6czZIcL8q4s3cWpSP776uCwdJG2G9dAe4sYctCIym09XP3Ac60rgCCmqi
XmbfHlwGdoRcXs7Et62J7zxGx0j6Luq/byHheYvZIn2z1j6d/awxSwpPsdn+lvbKbq3xog2OQ5Mm
ieSSEjFt9M8DczSx9aWKXQPdkM5/ACqvxkNAvACaw8ePc6/8G14KEPaDIxVb9SxaS21lS92XfK19
W78mCEUME7MuGBp9b/KFUb0Z8Vx+SoBtxaXM4sdKIGWRwl0qfR49EQrNvUm2fFZsouFhx8PdnwtG
L4KKxk160iv0/ZAh8i2JWAAatHCetJLwo86POMBdEp8Ny48fMpnF1NiHVmLY11TCONAEFnbO6cMi
rfJnT038u5QLJLWXOOzeCwvFOp23B6ABqcNmECZiiduktMX07fRW9RFpI2pp6/V9XR4K8fp04R1Q
vJ5NdGgENr+DGxpU+dA06La/IjpE2wpHquqbDqMPFsDI12qqxMl4HQjWoGXh9lFoyCvMFY/OcDyE
KU11QKeg4Okfgaed02cQXDLqmAqhMXVHH6yODS9N8dodmVSUdgS6pqz311pKpED6guwZxiimq8d1
Fj9ZwHP+5v5i7EucWVqUKPXr86fHPCNbJl/nosV6N8dbSPCdSmUWny99/XGG84qO199iMV9QmZt/
QBENBGjAUQjdvBakyukTQ0hxSDDRI0KGXhfsaxLgDT14n9wyq82ogsYn2BNCJ2LWGFUfLAnRfy0a
kwDFdxAboj0Lx5/YT6O+2VeezPieQBUvQPOucWk5iJ9CSPbPI/o/I6vGcNveFqMZeS6S8sJ6BDLB
fo1zwxDtbOcJFGRWr5tcCaYNRn9YDIIFBvt9bRhYRCif+wB1ZbarPNBQGEArIHsZzNIT2Pxd+Qg1
0iw9YoZUGHu9Mdinr4EdwnfmddIOBkp3t8y2Gyej+txHuPeU4PL7BVQ3p1g1Iknwd8IFHftWES2q
aW1rSuDKYaGQJJ6CNaFgDAWezcgeZU0QlCqfrmlIuzbsO2HeRZLDDOoeYCrp4ca84B1SKcO4ETam
CHOK/3bX9sTNH60XBCJMG8VnHV3aQoYsWCQYaHB9BpswavmtjBBgEiasDfzwUi8vw44ZzaLgR7lh
GJopTlBlCP/RevZt245SQtHMrl39JozJQF0jaREkwlS8D3GKJ0LngG8FGiH8IldGjxOJ3Hlo61Ip
uM4SPfpIo05eZ6ImF3YXbfSbVKwtB+TgKRERSSSgIfamW2xtB2Nln8PM0z+C9G33Y0n1v10IFEhI
Vcl7rZCS+uQotSVE82Y/33svex4ZqqhQNghamiE1phWKqD4B4rpIHKt3O1O41fDlaxL8PWNi0BZ6
TsKRKIg7nRr5IMJlDf8ZxLu4o833q9cNOW1eKVEbr8XuTcXpRz7f7s9Xv33uZGLuspDj4U7M4J6r
1mxMwkD2s2hugsQfP9Hhzf7aNWoQlU4vJe2MILtGLM4ZQQWRsD9NGSr/4gMAChflkr8ZXQJTjrXW
E8OH8qsaZRskTz1kQejIXDPUMgkCEjr8IPS1M42ewfZkFJEMIQNs5gRfs6bUzcxli5B6EK1z+wGO
dlb5MaVljD0w7gcKc0iUls8mBTnU9nyGBcnHLCrxIsUTkobZ2SRVZBNFAY3zNRx+nPNXrZnPZo9c
hJo1BlOHFy1tMbFRD3ZOFBsH5O7HCv86BfMpztFC0GaDQ1KCjbnsLncaI9UabC+myPhWUOBPSiYe
ZUrIGxA1dJY55xiP7JDZ5/QP+6PPRSSDEkIx6yt2sre0RB1EnChIWyeaVYaXoMwEd4ShRhaS7FdW
C6GQlIwXarhSXohoIbBpmUL6GK/9Hf9G3M3Aqdz6Umz1vZcPYrH0lT4t8LS+vqJ+IRHnjwe7Sn7y
T0nis41oaWGCFBG3pqe8cKIQfa46KrUrEcHhKTzhBk3P9IY9U/HXQ6xHGoKi4M/LB23YyONH3B8e
0udvdXhw5zChlktCVt29KJoetd9X8lvTrVYpacS/EJCQe73Q1TolVWmK4GDdq57ccMC+JyJhW16C
TJdgpyrwf0YoBHkgtE23tvSQHt9NBGRqlPWRBb1D7ByN7P/j3ccymdGb3cldLpmza4O5DCmt7PHf
GiuuWHmQwZmGKju6BLHs2Ur4QTXGmyRid0XdCNn9k05lbJKdkG3bJnG2txfpJFzMjcfhX4jfHcmR
og1fIiyu5usiElRSeThYEOOdh4v7foDDehKSvfKv6r/FUliYJzWchBM4ya+tqo3GmKTdP+VB9syp
8pEAhU2HVWnijdB5pmLSy4DJKD07/orxv6Oi0xIMg2J96ohNLrposAr/myLwYVoUebMLlU+FXuX4
lQpld2cgCAurghoZbZSkvTun5NYrcFNkFlmmhpYEls9Co2aIr5mf840EzuIc0e0GQ7I+Jw9sK3Uf
uJbGKiph10Df3fXzSD2sf1LGUpJnQJeGeq9bXeq9K/VFNB3ChQmqg8laCjfKa8KgQg6zMd6v7zOD
WTDJMLjQ1lt28/FxzJgwdknrJBpdxc10m8y/OunLgGPDx4GV4IUd8e3o7TVMpK8yfXwBJkIqXq9+
qBJGyUDIJ867iTuNKgQZ/bbPLmRZK/IzCL5xB9h+VpCHqbAA+MTmKpgWt2Wn5DQEhOoTer9DEr2D
w3dGtcBQKD8MAsgG8JLf+NVVR/cpGHpGC1YAId7FbAkFgNGtmZkTJ8vZLcM2BEz4tOOOFlCaWmC2
3iMemK/0Iu10FOnh8WKSIHf9R5XJtuNq/QGOlmoVtBcVHxv5qvrsmFc7H8PhKc7X81Yf7M6wAD63
+C1NUI5U6htkw0ZAdtsBZtXIJ2YwQ7rwneIKOJrKlRH4Y8AGMukVJX19GP92wPwsuMTDjqmnhAot
QYF9nd7vkFEM5DT/x3lhS4PKkZleNP07e89w4Q1x6Q2LouEWFf5oiR1+VF2Fl/rjQrKNzUrBSsyh
bjIm3U0dv5ox/vlOPu1JBzY0VUO5GBhtIgBxWHwkAFDMyM1Hn8KDuiA3sLumPRdqkF2oFVj6YBog
SRZsAIz79UbUypYLf9cB736HcYuvPHg9P3srwn26R8ouuz3C/lyJoOXQgNSPks4zMPUKVEhv1rfi
XopYSpvs+mgkPbDOen4j1t0SY39EHVpx0gOPGghZwOHMlB/aITB66TfHFHSAUi9t8hB9QE2We3ju
MvxihkCGtnfN+I+JRmg12etPYD+YUHOIfOx2jSk6YNwi5gk1gA/55OmtOW+Ke+KGwsAlbJDU/zQW
yzCvE/l7MMhLYDRPBv/vVCHiB9dFk6OG1I6O91NDpFiHBKVTUct8jJakMtuy03oB65+gWL4d5z1D
TeR3eDH6Xg8PHdOoLYKVCtREEmn0Hn8R1nI+p0131qIXrYW5d8aGkNzVrzjlIYu3MQAUDLswifU6
JcRQ+JggHl3Uv17YNBwztpxK+UuNZAwlFpZ6OzB9/AyEytZAFzr7GECZqRSy+3puK+0jUxVX9Wzr
2S5frMwr0vTwtvD4T/hRiYef8gXeS2ny6QIrA55up2HpG3ELjzXChi+uXOGR9UrrGhenPCNu3i4n
dgxGM3ANFin69qmLtG3ifHOTKxSEFtf8UW7TWQW+JFws2SCFuJSBOlmXtrHcvYI9PYzGd0APwNB5
/C5mSkKH+sf1B4fckhEISwyz9fVy/b9LC6pmlkVBVYZVOi89mFfg2zhdlT5iNBNOgApc2IXoqH9I
E8S2Cz4l2L41zl+1ywb/ATwRmsVo0Gd2szbPTMW9r+BuOwZMZahr/KHuM2QyhNLA5S2sa4B1kr/E
qJnSr9BALZHTCZLv2BQEiA8sfufJvWq3qsFow0qByu5W4Emu8bHc6wYngn3woGs9WQbKxi4OE0IT
35yw3R9mVFCaO9/i/KCZ1sTQOy85hniVKTOc9Q/Eu8/vKsqfdgMrk0ht47v8ktUUUNGg/do0pY+U
ORTJxrqIyqcg8rsNZUoW9JSKdYfeNJwuzL8MkKlPScCHnZGV6xBEIM2Z31GaiYEdYodwI1g0G29P
Wpp0PQ0t5btWOWIela8yNXGBmfc/neiTH0mDQFAgnmfJS0puVaZGdoOa3LB8mprUzq12kqMqUtON
ZEKN63SvTW244KRdMzSLQt+BV/PFtbejGRFfX+bJDf4mK+29B41kbmuPghOBmfpGp8FC/M+cU6Dn
+wew5LEDqVN/sCQ9AFuD3Z7b8zbaqXHRMgf2DoRu8FxaMRzOIlHnQR1DLARFteuv0edxmYGyZt2F
CNIexOtEJEfyw+uaJSJLKjZGJlCQ24y0+TY1/pybA/F3RuSQGS5QMD8nGSOXkmxcvPZJIWuEPdZB
H0Td9/+VERZgORWQ5zTTMtazpm1UVnse7gQ9GVf0I3E3LB+amAlAiZq3RY2ImYuDWNv1YLJLN3rg
FgRMJuybrl2cNB5CB/wykwo+/9F7cWZAeXolQnGhi2tdccXQu42R2O1kRcTkALK8zbqVnm3qMP7+
7rpZdPZmb+woPLzU+L/obRBOlvQB8R1SoYj5Hot2HNvqmOq87kVXiKQdcWeGWjJbZEfZyxgBtJKe
sISr/BDmM+g5Xwj8+HEyTMMGoWU97gN7AXYqnEoDdpfiw+clWgZDw/Etlh1RDEjoQcOgn7oxjNdI
Fy+3kZXku98nZm+RTRGqkKOfXHjIiFZ1fIXI2yhyrF3T0azUwQWtz3XHxs1676eSv7g8FYVICBbu
1kD+rk85LMglIPjE/m0jr7ncbOj793kCRXxEDLlyR84eBeUYqQ6eWGmRyHsY55sVLoPPTjM+cBGz
dzgt+YDknjNO4VMD8C5cGvjCnLU7JyxWIkcis91yNQl4aBdvtvct9QdswNBW2rdBj9PuPHGqQGof
nHdNy/gf+s6SrgFH6VsTv344F7Xu/yOzBkRiEZD8nNvCmAhKlA4UjNUoPPRzxaZVIqCdnhM0TrCu
M48Ob5eN6lyonXxyEFVlVUgA/h4Djh3TZ9XTC7RWVsKez1f554qh20ZGbseSaluSIFHlZsDutmfl
4Lqr+fSzF9QLJ4JRX50AWKvgfV9f8oOHIXdN4uXf0TklitcMx/BjYw6q7kpxzwF2TUP/JF3cYi2a
4bigsjyW/LoQ1Xb9nF0LeReqasXwIp/xcRGzjmo0p8gOBFFQA9B78FpyMIeyr3h6QQNASxsMevIU
hjqOsnqB/kQBRMTVGSSSDkNc6q7yoPZqAvpLM7uuWu4N/KVKnVls6CquAlpkCsKmrkdonVuILOpc
xEW3I0QTjG9zVxv/5T4gLS5URz9QNYK6U87euKENbg2k65+hX/3osN+tWJvcFk8mmQtuovreiyeN
m2PQeQv05n2937ftiZ9nifWBqjUkmRe7ibkvEO8FToQBYcsPaSp8AxUJwM9wbOKkt33i706YVA0Z
8B7kz39KE/zxqJG1NlgGukD8ySEzZR/1cJXaRLXk7NT8gmxU2T204ARxf9NQuHfNNV6+hQyINQTu
UJHh+o0ZNdLiIY0IYrMBu1lpZR52kHBUWSyLrrDsXWLA3Nhlp2dkLJJ47HolThsaIb79RJp2sGKu
F3gPy8H68xbTLvJMOpAbxHSiHwPoBxT5AMdBYhiKGBhIhixp/Tmh+qH1PKAZYmStrmY8jGmKgGOo
2wefwu5eGcH22C6uERFXcXcnrHzBWQ6/9o9UUzMzENhWLO3AqH8396iVknzmN315BUOdW8EV6lZt
K2qeTr+k902NkZFLJuYolZ1tAR2xb9P5EoRRB2fEvYUATrvPlQCmDjmpzdw2FTSfX+lZNZtF+eSy
sNvnvLPX0a0YXwcz/1cdnFM1XmeN+n3r5zCopws9gjabFwGUp1zqdlDm+cOCM36NfYVmBBsX+KNT
F+oxtXjQCGEsIko0zW+BYmn2wZB1dvdRCQpRWWWsEiro9sBrz5lM+Dsr6HGUMjtyJ+hIrQJ6pkic
BQzRsjM5xhK5bGRfgdy6Wn6CHdyZxSEJA5FEdHK43TyLi9fOoMnvzEUF/QTQz94dvv28MxZL73xd
gHiwTLw1jlYkfRSXekZL+ks/r2vAjMys9WfxHm7yg6Hem+oG8ONuLqqYmv4wH3t9s6JxiCRY15e6
VbZY6ZFjsPDUpl3xuOSxln1cwcHcpD2jNIPS9WddRzo9jiEo+qx66n12qr1DbVsPsNPZ8saktryJ
ufNlJmpMcfi92UpivMso0F90XTrgqequ73Uj4/w3j6MNeKA/kWxKt8spDRgQqrJErAC1f3KBthQT
GbsloVyKdkA0bVEICvx6sdU0QbbL23Zq15q5fyLfYgLxA449w8M5/Yr9aFK4+R71GMk1Y0e6XmY+
NnD+xK71whD0LU0TSvc8pt3aOHJmSE3JuMrJydGyY4JrX/mALERka6OvNgTdDH6aRM8W0fLPLVlv
tRxU+3yHB/qLKuHa5xoUctO5DpdkBSJHpqBbQe6M8HsYmDS/xkQBAio3PkG5ZRTIeJ13v/Ky3KFn
wo7ww9wcNphrQcnW7+5ZvG4TzAJFVGBtHn9DRSlbTgzTf/xx600SmkHS8xmZ69s5Q0xHKzOnQA2C
8HOH6qpg9jnvKvQ4XUg+Z4k1CZe0a4anCCDrnH8KF7cn4YYq7c0ercUGHgJLddg57M5IboJF6oFX
TpnO3EouHpzpYoc9Ev2aTdTG5nx7GX5bmPNVyBn0tsVZ/KGlOniv7ljxMiUxesYLsdGXbPfwShQJ
I6wHtU8bFGTL/q1bl/r7hDXmtJMf4mq3vdr6bUR0XEMCzNb6adQ4tWRXFEKN4XQm4zUyN/kI3fjl
9i2KohdYz193Y5usEFA9gug7wOlLLMU3DovZhQRqQz9dpUls7nRXMSYYOvNHBJrBVEcl6QogXU1d
Pf1Lr0VqGrRI9ryqC7YIsQ0/Mq/P6VPuMzvEcuWl+pgGjPzWj52gBOnG0CrG9gTQSKs9L8kL8AMy
wyag0LNORW38SMzIRfV3rG68cdmirok9rZV0IotBytu57JPtOOoc8y3QtDOd5NxsCgm/cyBeTeHQ
CvoOEd6mHHiz1E7ptqNnsexEFQXZ2989mvfufEKXie9hg/RQJ0wnYA/KLldZPW+9zpVcoryYuljA
2C/WSdpMqPf+aE2MT4rbd17W8r0HIccwQ/M/hGhUdbu2P1FpHVCiygcckTS5RM+VXJ+M1LQtUp0L
OXcsvRHcwbcBh93zP93XCnbfa+ABFORmquRAHnt+WMRrA6sHVDkIZ92Ew2n/4TFA08YjRHU3hpr9
o6VJiUfk1dxFe0qLEfoW/X13cc5Fb0UzFSrDiwlwY7obPqnotFnyM8/inTz1OemIvP6pvfHxTaOe
aZdCo3a91v5CEM7atY1Bd6pgJDSzHDlX9lV+HVUCB5cd8lXp6S8osaF1R8aQEXBHv8KDsnByaPdk
r+AtVn0G3wByqm3NG02Y5495MT4ameGk4TPQTZU87TYRMo2L/H9Dpk3eKKwAVe6w7NHTPq8SkRq/
aIIj+gH99cWDjfLgWzytPFKxJgNaCckd4NMimerLxCUGa6ksG+ZiR4eFTmGWSVbo7BjMhSrPujGV
F8bReG5CTvape22RhnagyXC/sOzfUp1YS83ujx9G5Mdq1R7MPxVng0n5fRCVMky162oOiOClIC42
ubULtv96I1pFbXpTAp8rDHeF49QaOhG808xBw2/mKd5wtSubaIV2b0Z3E6GJECbLg8eNP1gCVzDG
ZW4hNzE23akiFPJeWAc7+OZueb7qbu9C9sWZE39lyH6rK4fFeXlElY1his7u+b7sbebb8doCZ40j
CpHTuFILvaepSE6TicYyJNFBZQHAvuRrUjBhhJje7h2X+TJ1GAXRYuWgNlpZlIxgf/5wkbtEM7UF
jmdnlodvu0Ua/n7GAryo+Yp9+bnFxPf0JZ5YgtWi9cq9dmRIHGEYJEY5d65RW9g7Ma2aUCcOxSM2
6jxxHuBnVJaK7JuPck2Biiajvp/LpUB5xI8kZFSdh7DfQ2mYLSfwHlmK5NskD5gMNTR3h0ueqKk5
I+eJDY4zYo1uzjZTFdXZDh6/x/MWG3lHw/9ZutVCTm95PNnKAcTO4pSXUUNlCW4YwCr7frBWIjUB
AZEsBIRJICgXdRlsLp0p0OldqDbUp6t2hRj7KA6SPYwCorNowex2r6NAIqVGF3jlkS1gXxN9rT7K
763Ao3RlDwexidhV0ExWsL2Wf3a+l/FcYUomO8EoGRq3r+FlJCtuva75pxgt8gP63rO1CoHy4VqN
avQPS9rfH2lZaRFBsC3ngbY+KCzgiOu2atMM0FR3IjCMm6qEWqiMdCIp92imvFBFwcjlPT3fmG+n
BBk9LnEkM/yhJJMpZIj8/yJTk8qkXzuFRPrFpvA7A3ay2ES7200t5JWgzetWElBX96Yl4KqT114c
gs8tRT3cpkgO8CnWdKzhDc2smxnOd3KuSLrvZoZTSVJmbad4rfwQhOcj4CCpVVD5RpP3X0mEyTZA
DLuOVUOYN1jfaSEaNZUjMEAvAvHtA4Fd1QXr4EG/3AijqmlKNO+MhHCIc8VH/xWn7ujGoykyykO1
ZT7SIzJj/NiNH/MjbZB1kwJ23h2FCensANOYyuwM+sTeBUNQZx5hzeqzF1d9hWWYTZmhINqvpTAL
5P5NzIYPhk68Ct457NL+2aR7RNlhtb2gcAbXRmrQGCfppt6FKX7iaIQvsLTRSuF6P2CLpeIflDnc
j1cVUKS2mn9jP8hZjdzDJuTUplYEjQjibI8xTzmKOj5M87o+uNQe2xXMyPkfBfkSFDndQxMRD/JC
DnV1N4bFpNoiep1/HTX2uWcCWA1XLpF5sfhvO+wdu3BGf+Fm4E7Fn9EsOz+rBwODe9GAG6zS/sk7
KunmLIDPG9sXDJYoTyp566XS4gB+pdtI/0qOBhMqAOR4VllvFfx9xG9fzW8LfEIP/QwfJtthFZ4n
GTdcxgjHV22JsqwYNOoGlAdwa75moqg7wsP8GqlZQRYfY+jFnp0oAZknCi6Wp5+Erw/t+LjXt2Y7
tSYuTfjpXOj1W70s33LsEpqyG0yZrSv3qOYd51MUwwz+7KYyWFldtsM8uecu40sJ9Q9NIGuBncrJ
W1wJeh/jDGvWmB13AMkg5n0Z9C/PdOiVwk+xGxQ78/OQzeKm+9k6mc/e+yvEsXMuvbidQFWUpTxr
XgvXrNCG4PzRGoON/qZRENQxi106a0l4QwdHJTh77OpPY8uF/gQUaTy1f77GHcfpQNQF7ZRWe5YT
zb0mKMbmOxGT1xsbKhCXel9ZFzgPo1Tvi1DpIa9xZbUxkjqqOGQ9rFrOi5gFcCl3FRtAC0kZFpwx
9nR44IL3hP5BTQS82fpB0JLmpzCdCBuiaDbMehdpsG2B3XjQvNlDSbdZlSXFhozKwx2PHaF7Ugte
sECOCjiwI34xX1HHwf/KKUkX8lsdum3L6C/nxGph88b67S9YBGaQ/5niNZo7BWMfE/YKvrfHGIEp
dqrtlvAAcODexdxPrY2uypXrkQHMiPw94OtegSMOO0hW85AXc+8uc38OFTv5Kw2q/pYThUgcfIxY
s2sem8+Tr4piRsWcdOilGS9SIhRoYYV6NFiergDsdtXu9cqDKhhWAUkN3nDJTXfkz5B6SlAcryVc
gCBsNHiFjJME2LwBA7rOnFhcn0rUgyBwV1Te5VQ+kiFSw+saV2HZVUj/6Wbg759N92WFHHIF7TuQ
xXUgnNeOjbvdZlNzBFgepcbgE9m2l4yEU0Y1gjqTOwiVU3eBntFaVElgG1tVuS9eanF3PPR01BHp
Jc+JzxjNRLbuH/ypCDUCb/AiTpN+cg9P1LokEagjGBYcS4X6vh2TAdqGTfHC+2VEl89E4Vvo412l
IpxLUo0yGZN3g+zH+mOFLYkBVG9dzjk1aSCYnNVmI5lygI50Pm7yDI8P3sZUOuRVCWFrawRoUvWq
/du+h2hUMd6PziVNjU2MhjoYJJKQs6G2DDEuU8NFGA6V03MwCXG6s3Rejr87v1bMDO8bTQptoF94
4pOqEDlQEd4+iIc6zDwJbYO300asT3UwzZ+5PyDpxS1QYC7as2rPxQJhizCOBp2xmI8STfSmdyOs
gip9STbPCZMgIKjm921BICcOs2+hz9nq238oc98SqYrqZstzdAjgauEpNz1TweCpntR/PqMAOghG
PZeiLg3QU4WeAHDIWp4CfBqdT6uedW4EQP0dYALZMRdUK6XQWxSgMapFo4ogZFKy99j1T4e12T5C
93r+O9SiApTimMYmxKbCFj6xpwVaXnntPIgM9uQdaZUagvpE+yWNjD0Oc3QCZsbbt3qsUegPSC6w
faW4gw4UNbcymkGy1iwSSV380rCzoOg4dIMoIKQ3K1HtZc0hCXUCa1H4C1EGwaQYQOiGW71VK3oB
2eWNz/Y4qxutS3JBrBpCvC2nGNiK5YN+YSERJlMwtwQA4VjM753yq0N6PwsNqVtPptENeYd5GjCl
GiHnprVEoey0ein6U/iXQacLyXCP/0XTRrkzgJ+Fn7XUv5euOC73QOshyWbBZQ1t/kXgL64lHAK6
+vaSTKmqAf/xpgRdHEWoM6oH0Pi5VTBa4dm+b1i7U5ULsYQl3IpZ1JJ/bq7iD3CXVCzXMSCWaN4x
9pm3iCAC2ZD3M7YIuIt9OvoYQ906E7iHTh/3/R2LNacR7IdpInNIxk8DaiyvHJhQ65Hk9Wk5ahyC
xje79xUQHGP7H1E1BVExIS3upaReItT4W+m9Mk4uobUdtbj2rfrxAak3m+0kIgHgKHwj0vxTvHaW
8tXFfNJ7xmlFrcXpsOOkVqv4Bd2mid+LWbztkB9hzT1sGIJ2tFBD1n905FyWhAXdKhYnKZDBSZq3
3GifrpvoEYN99ZWy0IRGeaCsWn8Al59oeWUeciGcWREleQeZxNQSFyRXzP9QPKOsqfokIRh6Vnqe
YLOGaNbCMp9KWMxS7yFw2HwBUllN8Q/IsrjcZmO6t8W6nrQKtVVh1vMNR1shCcbuSoPxXcxhOGuS
9pYUH0C8HdtgfjBs1cKzyaRrcftMk0FhrGkHXGtrJ5lWe5QGm7N45pNipuS2rYFV5RQ/w6uWca5k
elT2osQrrDlvwJoRT2Jvyw+Tly0YJ3GcMaRUUiX39OPE3h4nBNODTe31dUGEI7Mh060kuuuIpgoS
+A9THvX6nr8ZjDf0qExoic75h396QdH0KJPr1x5o6nIBeqUVeQ4u/xxcQITpw+HzdfS5s+GXrf6n
+ffqnr9QB+jULAthIU2euIhw2oDEJt6rmPjDf/jrBS5Z1n673B453ZdtaiK+eRwOxHvmLYuZidN/
93zJW15piJdwQBDnomY/g1r9rIhToSrNmVPBSt3EeRnjRwpLKjXOfQm7tXu87GuwVSUGp0dZ1hTr
PZTDL/BUouvyST64duqnzNY590cDGqEHeAvERgY2OanMQSkowGi+cs9MdGuj4kK9WVZbFJcaasbn
uBGZj2EjxW86eSVb1b+pR9lUmQWRR8evf6rkHXf9q4CJJBiYhsDyu2mo9jzrIc7RAQShYsHMrzyn
a7O4GGF0DPydPrl5NR8WzvKisUE1dmTUMw8XqtxO0mtgsLyw9fF3yXRqRoFQR6oEo3AnuWBBOPO+
U6aZxtPkZx2qe294dcBy7xnJhNmo8G2adqdBweeYfMd5d4PVIfJwE+mW6hI/4GrWGP96ll6aS8Wj
9FEbqSTtswcox/k8wSRHxHRMbK496kVXjFoJeps4DmLVIDTUBRJ3mQGtv17PXmu4mVTrrFqBjJbm
VHdLo+dSs6E8nYceOQrXr3AlypepUT2EozB452loNTp4l4621xcCghMvA1WVwrZ4r3Igdy6KEHvj
MIDnxn9PWNH3nrnq6ke7ttskiCS+nJZKZNblcXir9WoWJPM7dl2xAjac5GhYQ+33xgfIUiKLHs2e
khHOm2uOi/DeUcxB77qPAkckcK/6e2Nfi10MJ9LHqNE4udZS3gVMgCRy2hzGRGLiE7g/7ErZ8y7h
CcDFPUW4rGA4Np99EOu/BqX9ixRuPH4t5PPrZAlKURpOHTXW8w4oYexOdR1iKaqWuZayI/7HAD+f
itFzKngikqVvCxyWwDQYA+1Xv8XvLRUq1DAu0aPsoEIo5DOAeo21frj3YvFgUUYqrekbQFx2ZBkY
uhOhAFjun9uUkspn6AELxgUzrMcVCO1cK7XS7Sqpv3DCWoExvG0m0HvZyKkVDShQXJ9oeNrhka3y
oPbKtxnO4DEUfFzLWK8UcEkahw4vtWPAx7IzgxgFN2QTZTTSxUBRhHtuD74Xx6oPSsSptiFW4Ewr
Y6Rcd8XZEuBxQCQ/+Udm55oZIV0/dHQe+2/qb7MwBU0K5y5IXPHRyXvCDhZiVPJAwixjliNCodjA
x6g8g5+XydKpYSK9XiRS0CNamHsh9gKLndJ/BfuUHc0nvPmjl2qcCmTaWbcdbc92FZ3pPb4g9uPZ
ix0/35WERuzQh39v5QbMj2mTnoB0CU65iK6rOc7s+7jXBfkqNzkwBmPh2EZm03nDdAqw6UuCvFwQ
1l55SUZqINM6+6Tckr0lFncdmikX8kaanClbAqyvKeK+VjcotV5+07P6C3esL48GeeobPx0JE9xQ
gEKBMSCeA0nHg7+/YdcRYTTcqnULTkwh5utB0y1XDIyuUsi1YB/2Jr4NKi9RJzJyuX0SnAa/oP7o
kSpeACsOwJJxacDbs2g/AucEJPm+VUzcbhwdZ/5G1P9OAMEWJr2leYPQZ9UZ7XxM+MnzdlshGIOu
rc08e1G8JKtl6qTB8aH5LcqEr2ZJj70v5pcgPbPdF3Nd2vEd22WhukwNzNp9XedyiepPNN17uh57
YjrWE/aidFM7YX+p0KX6GPcR8QH2w25tL+gAkF/keQEezMyuV2yRJUbXHg8YfR24dMjuMHeOAhT3
1BQ0yuGu85P6XCo38ivGCFRm5pk2shgOXFBY6GvWWmembtq7O4I1G31X6g6VI5MXCsPBYfaPHOQq
viWaOulP06CYoZkPeLNa4jXMK/bVnB5HSDy6RdVfUV6gPTRuSLq6rnAZOjE3JhyzRqkPFtBBxHiT
b+8nu5eOzv1kYdodhchZc6jNLO3k0lYuCLVRXmIz2SytEJaBSZVvC3dnhunXkR+k5V1hCfp+9ObN
nTTgzYmzzEPYKluVSjNhjYAyY+aflseoGPUyCptChoO2LY84AKcFjkIaOhCTaEKkzof4NMlrXKeJ
ihDx0B2SkSpI1rGAwbznQoPr+lW8kCEM3xDJaf+HYhLGIOnwkIM9v+ZBDvQT2fRNUhbzQa8ETCgG
FXGp16lurZ6HBCfERpaDjvffOZu5qfJgZWsQICYimkNDWihGcy+ZsrmGGZ0l0wfapZH6LS7lQcT4
8Xz6mrhP8WE93QajJIvI9XAYKi3UJNgg9JWKW7mpYuZ46yv+zcxmg8fRePF/xWPxC8JB0TCoSp1A
iZqExq4aPw3oGGwoL2BJhPfD0WYyn3jod2pAH0mIcVjdYS9ux4CWx1PczS05DVKnBlRdYLV272kR
OQ/9jca5uG0DGAQJ/qVBjD0IWibLDbPkrMFIZoqEpvT729Tl9nso8qZKu6wXggrEQvqDvhxp463j
3XkNTgnxZTYL37B/h2osBTd1+Fzqycq5ai97HV6EziHR/zP/m89B9Edg+BFhWh76OPscPq592nyW
EkKaR//XTlCY6aBX/Vh7eFPRlbVXyftr4ZaipBjX3ZPwA6tNV5OeUjycF21159bDvfTUYZbK2Wt7
TQkBFd3vrpnB06X0x4dkgwtBu5I/tPvu2StgjW8o17E8TJ7WOAjkn1MRYrfAa3KaRFsP99hEV54k
RDMSga2orLsH7iZX/wzxpaZ7ZgCQyAEBMappj81VX1ept6E3hCkgPHJw8cZFrVG4BkF90+Dld0gw
edNZFl6mtf6uuif6r76CN76VqqBZcI8Nan5y6wXJXCOzxq3Cm99BYVBaNXsaK0jETdku7JUkaiRd
miLlxip1TW0l6KIda0QdpvTPf4DOQMwWhY4AgsOERaxEZJDMAWGG1fH8lc2xH02rtUhjmKfApBhz
joXpOw9siHrsrizitERxY0FeLQwdujXY3EkFhfQR2q/MX2W611gtypl5I7hwFtHId7HeVt+Ef1TP
BIhLHyalpWOffmsAgGK2ELOZ2z9dSFZEokOCgnHBZRZLy3rE0VRCwHSkZ6aqLlCzGtt1Yg290QAt
nf82/TEBVq1nO8c5h98fAABCufKjYJgOsGXTYud7mtzObFyYiJwgOzBJ3xyoz6xONK6ussirsuMh
JL1thg3tf3OQup3iPYi4dBBVfsnJO3SPsIApuFk9CoLM6GIOIuNWhYVzy58xxr788xc/pPXsb1uw
5keienmwM/ZWv82iJbQD4I4G95lj6Li1sbk4/VIntdYEdrTqemKc+3Vvtvw775xO9DVIMTV1kMrL
FOnzC2F4XpBoouYijziGCZdYidzwkzmldf68JBs+PjDAWpSEto/lePzLWhleW1sEJJ6v4S17lzj6
Ct+susVetNKRhLvjHYYB8nFFVNGe5oj6KX1S0WbRrDLWNFWHti6p7JxXlh4/24px78PucIjOgrat
m6tA80kGVEabDYukhgIKOVsVdtDB7QtaUtWunEId0Flo759aqghTp1L0Ug0TF5oKXBdiPwG73VIl
qtMeY5an5UEvXMDk8fDizTdm29FeRXS/11+oUKUSSi3B8PJLG8WcKGYs9Kp1IKRoBlOFUcRDotkg
Ez8NhaRYMji076WMhA63snaJ6EKrH6biqI7WtRWg3u1n4rlt48OMOXtS0opOB+/gP8jBrbCaHoGc
k35O+VE5hEh4qJLtq3QX9pmNSNKNfYldt+ITv8S8B+QNP4ZirWDLiPuaDyIKe0A7ktvM7kuzMdzZ
dgBUINZfg+lxfwBPSPi8fHfDtWGWqaG0mR/6BFMX33m1N4USDGe5RgFoB1iG9J70s3A4sprWyV0T
C6bPYNS4Vo4R3r+Meoj56Aq5NtlyUHX5jaUPlUV1r6PC8z7wmnizsHA4Gq/1Px5kDi5Isb8w9GEc
LMX/XE9RyDkoU2pqJ0ighGlhnanwc0D//UP7LW+qHgu1u7IgScUgOt9bPQyDFngFsu+xxv2ZoGZj
EKHEU+VCf5NqvijOngEU44WULoIDgtxMvrfRye/YSIwikcb4XA1fP/9RQBXaDUgwyeri9NBQnrG3
xvrf2SUCa92NWsqIHTQ9BVsnvCDDOIwcqD33TeYsGK3x25I3RGfDeUkpATT3jz+oXXnUNVoNO/L1
6ur6MjRXXxGMmp86wSsEfin8LIkoPlUSiougdZ262bHJRpE0ZwPRMI35p9GNXdLwqBBnoBCFzeQS
IYr48zvs4rDx1Jfgin6rFYa1Oy8hrzmPndAX3wphNij0atmnXFot9Mqf9Vo9E/IYcgGzHMJLEBac
joaAIq62tjFuOYCIl9bJFK+w9KGk0c43wCKDrPYTHgsGbV6iv9JjqOkaZxDjT14CTW1kfoe4GY9E
cxienUQ/J/VY3As79BcZw96gqbiW0l5GY7dk7Tts2Kuj4Ck+ZOQBJ7Jg89mfiFbJyv4bmYkKHc4E
Z5NaCBE4QaP/eDoZyVe+kAO3X0rKdd7XxkcsV4TKwkm4RIv7CcvLE6fkcvbCpSNpsYqVCs/IX8Id
gzreidekOcFN/VUXLawMlfvjRsp3jOUoqEMdELptLV51m1UmL7gcJpwxUHrvU/qlfT11qFCs+dDt
wzTTv4IhnJg6XrOOEw4ej6bjSda3+J8Y/3mJ0kRCpZQwViLppZ7KjyECK+FUkYC/vWVvL3VfdK8V
2jY4Vx3maa46ZSnvRDPJGxxqvVvesn8C7+XH+QueneCsj06W9QZJRpVlTtJjpHZvOO1D3SVkQg+T
WBivDEKtB7M6Bh4zht8Dq6YyKp/smGhXZxh5oNFuZ1uaAnu8b50448S7eWtGfaQWkJuYDGOJmonu
62ox4J64GriHdOpqHoxy1y8E+WTviGYrUfimdRfX5QVfWw+fJCWeDLIYBz5DZtHNhQJNCT7RIdWd
mI3/r4YyesFqXePE3VLA0RD1SyisAr1QaJKU7BTZLhZ1wJQtCMRc12bfcFUxv6zgfdd1Fx9ZM9Fy
U+5abSAg1D1wtT/FHq9OiXe9Sz1DCfOuCQVRu3dEOifXrzLNKpDVcjbd3RjVLBbrNcr1cy9XnBZs
Kt/ORy9neHAhJNlt+wRl0bP54wcPSQg2weyLnn73Jr1fZxJYtCkp1iFzP2ay3k4GimhAcfLScawJ
41/Kqo7UqypUyIGo05peted3m8oEOk1IxfOZT294vSxs4ZtfUMYd3XEE08aPdJx9D4xMruHsjXe9
TNanSihJPLhJbA+RzGalQgvmqqj3nk4iAad9sVowd/sEATGB1ZYRXcRK4f2ieFVvFfB6qC0zsOa4
T4XjitVDg8dF/olkQnXUuDX07y1CJNBqz6mCFuwJsq21K8Bv2lE6OzxsQOWdNm8qwlIHt10ih07i
OdpoDNH+HEX5MIXuerMr/9ELtRWkjCUabLtzPsPJZM9geappK3bn5Pu3RpC5e1+B4XMk5eX9YxKb
r9I4aTNPhlqJHJmup2a3joQrnVzHe7dnh538MD3p40dB0wwpI/ImmP0TdZRmb3AjPMTuC93K/3j8
FrNM2s1lj0MZY9wecdgEOMP3iV3YCZCoNE9KDw+kwvIgl0ouKzyDvf/yrwoMiDuxZruphtkd1zML
kYx7+WDuUPJxEDG5X5UrZZCEUpRVv5RZBnRAhz1blDK0RPeg7Vp7pMxG5ffW87VFgYchDG6qXnfB
P4RvBxES4bE19uNDRgNN5OnB3t0hUjLGkbPh5r2v5hBpUWwYsnwwGJyeswp5vjOGv5WLa/9gQ1fT
3RN65PB0DrhoxeJ7yoFK1wSO97P8fvu/+PW2TKwk4mUiGChFLYKFKiz6jvwFdolR8OxR8p++sFeE
TdO5ad61hVPKpsnldBYI0w9ZbRhlWgOZOIITXGEsP4ntw6jUT3008k3LZ+8M/JKLExnYpD4hVUwC
oDEk6IyzzMYp1ODFlu5xHDyhgl+7WUzryz7QjpI/kx3lYZAyTuSHvsEDkUs/ARAYrRt68nqE6D/S
khlHOBfUlBa13gukbshYO0rD8E0IZPgQhlf7eg4lXw1hgrWwcTyIxYDdGWso/w4vnl31kQU2Nsop
d8bEGlgMD16aScraVdM06Rsvv+hxJruhO7jWQrsddxkYknk05yWQq/9pSqYOkMgZxRtOjkunupQ2
N7tKrcwckEm4aQheSTqR45+x1sK63UCgOd4mmU0aWYOSEUPlrtQBwbK+0AaXtKr8FX2COxBuMmxB
DSiW/GHGN6oltb8RTOKVVbwP5Uyp+8kC2Jg+lvUQd8a8D1ZOMulX04nH1GTC5xhJGIEJq91zKZgd
ozfNsupNukRdsLur8Xy3jrB5bBM2tNPWFOYeMAJ2JZwYbIJm4xHGiauzdzyIGse2Z7vhVxyrPqvD
tQ80YEyEXt0R1j1MC1KKf3wZ/S62rVxMH3ggCbW3sQnpwzN8RFJGOK0B+7AVn6RZM2LFfaChy9UE
B6xkokbzDgGNd1Fbm5jHKuJeX+jmtaFFocT5qsZu1wRS0Wt+6eFzKQV8c1AAPVLAqHhf1mIqWRoJ
C5f70qwpuUOH/AG4mUGbJpZyQe4ua4YaFR8WTWMt77jfHpLCHnM0HFQxPPZ0ikeoS4sMfdM61YAB
fUIF6vHIMmJEuFJpuoDfjLgiShqvJktodpxMNqmC2yemRzQsLmmPXfc368FWdvM5m+sIZRgZxexb
pndDNgS/RJ4rFlOIFmIYiX+8wTSBd1hYrQ6jlpCGfEEQO8r4IUdH0QLNHTlcBqtFqrquLC2vxPy/
d8g1lerU7xAPcKtK9pIDPVvPKkjEx0dbojiaJptGOLlVWl6n6ZMPTc4xzC+ErB7XhTY70tu96aIs
531OMvpuHqyWdq5xS6YeIHaYDKQHCDiD2I+PoqmKI2+3q3i51ePcg64XwHyIuPC62WmksQULBt23
wmPz4MMd3BOhCCqdJIRlmjXDXMisiSMANX04VayOOMKCg+BRLexr+SPV+sePrnpUngSOdR5cEL9o
IuRcs5SwLVvnoms2AO7YSEzTFWRwlJrqsIZJsZs9cp43fCYLsdcS6PubbMpzdXKkbvKtnJ79uMzz
+9yX731ZNraIaPClSklaP03aJw41ezG+ZsKzRoD4Qqqgvc7q0VFkPQD5v01vUMQJ2zFd/bmxyhbh
Nn8915HK1BOqLAkCsL82IQJq0jcN+BffoaIcyCKKbRMzp66xV4TLWv3fkcnie8r5zAtm6+Yz8PNr
cSV17bpix+U7ioNl/MqPcgod86kU4DkywyMXEp9F82uA3bQhWbdNjKWFty4V3gwpVoKBQnvrCA36
PxhQh2UOmpI/+VWBiFLf9OnZT0EAhUYS0MFGq3Vylq0MO7MxlM3yN6bqCrgPHfEoe5b70zUlXI7r
1UwccfPX5HXmuTSSPhkHxEA9AWge/4KUI4DtyikKtqiodmqCjJaAp0jH20kZH0Pwtg893Cpl0Yy9
wutbbDzSEI4xNh+mvg5/+e4zPaOtkM/GHa6LBMHVG6gZoVZgZy8+dAtTCk3nVs8vI0bZbbL2cjVY
YZTLXCzZXDmnZ+rPZSfDGJ8dMgvpgdonjBJwSViYuBxpdR7Qy8RnoW2uBeO32ipyjIWcV+ZHMRzK
nLrmhn0jdQoIsb3nxsE8rJyIYtqXaDANKUVkI8vDsQ2VjWW2KZ3CpfsJdDwsUJzP2g5XrRs3HO7k
0ar+2jWu1Bf8cWmR87vb3/TJb986P4P6E89tMXAnjWDn0neN/LMcVP5MmJbosmad+PE9Z1aDTmdr
cviClfLg/GpU7ue2HfCbVEMu58zvg+394STCm3K7G878raAc0pjyzhT9L7lvF0chYOxCd5Egriw8
tgt1R24fXXi7g008mvf1C1Qk71MDn1GCsELIMQrk+RF/aEx2fpBmgL78d0GQSwdoK4SCqbLfbeIL
GMV4FbjALPR0V+s/KNEjfqkLGYPuvF51xrG6+60bku/XbdtgtQYQuB4ABNuENWzAmbhNipZx7n2d
CxNzX23twNELXEFvHnR6sajkD4cEZiN7qkZ+HUcBxEl4eWlYvT54lTgpVpu0L3eCTfIISCK6wU5l
qlAjotl9Lwe3GxckgyIblkXNVA3yFZO9zF0Nj5DXLcinLRUzh99lVLvd9sqCDtcINJYXdFFNIu4+
XlxYbf0AJkmcBKPInarX5mFE3RcF3C8GZbYU0q1EH7TAhKgoB0evTc2gJskRTRXsXeSVzNUXNKXM
QcGjlipBhju+wFiIhZHunCNCdlr3OidgmGkpwa3xw+cah2sYcRasSmYpdPgm3ANxpMlfD1vI94Qn
l0hWQ36585Q+oztKfYp+WaY0OSC3uEghO+8Tb2SiQ0hM3PhVNpTlx29xtHWnVWmHn0rH1rxoCdZq
6NddbjaE02nttAeFDrPWZ3UwwCy3NutTolDIYUVaC84oBD0tkyuWU/uI7sOUccXtVoLFN7h8mIoR
tA/6eztcDgcluwbr0RDp6bCdaUCwInHAa3xn00EAQE0xh8tnZl1O1lpjCbTP9q7KZCS38MY+Erw/
mnPMYuAxA85F1poc+cDNv1PhgbRo4yp0cQL7wU78CdkrfSqQg/q9KW/oHxBot8uQ+KKkr/6yMbXT
qoMr/COZyDm2tcALEVkeQUXfuQpZfUPZWgxkLXgWksd8rd00KGOvJK4cu1hh7BmmHZU0lmhf05r1
ClXH3hJAC4v//xXAqjqd94ldrfiV4mSSx0nPOfYLjys8ai+GYI53RTzb9YFPdVGwNk2Q/4WaPVin
WwqpRt3j/ttTDLhGg69dz9l9yi9GZg/B33leSK1PwpesR4qgygdpSL539fTdpGoRjz/F6kN+LPXy
yMQAwu9mjKJPB6/XAVFV1ndC+hEMXrQy5fCkqHXKC8yG46oBGyACqMXTAxyNB01UXsasb1fBtOIH
9jsKl161yhHVfv+TkOI6H9fQje+jXHL5djsWxQynvmwBYve9QO/JVxpXWB6xV0ONT541rFEV523o
RkJS9YvbEgWMseSM8bp+88BAq2BMCvgu8FQ6pFzc8XLhs7HRk4rLvjvlvGV83fSr+LPeu7TV4iUB
sLBQtTqwTtJRQtByf6/ah4wp2ZlS/A50XzoRd/P+IlsgZzDgcyCfcuXeoGD/ns8TmWWo4JvXGv6c
MeyE/3knzXboHirtK76P4OnLG0y6lEitt9ZFMKr1JDQDQw6nOfvjub/pjbi5vMhgI1cLPQmXN+mf
d+bc9+ERJ3TEdTuWeEVIbCXbtQfgGZkEq8nZKvNyNysEkaFpf/hbhINXUhkab35cKTSJH2PlmccR
0dqgHGQK3WVWuL7vVtVBuqKBFnMCrS4ja67ckxc6TIbK/Q5GaRgsRgTtgcl2JFEE1ESgqwgF5QRW
2o7mIgrAmNPhg5YgRV8byDDfiKuGhAuMGPpcGGehxhzCIh3bUpfjDn0UiXHeM2bu1JrMXPhN6ZVE
XNEF5G79LdTl8xUGyABEdV7iSXCf2GCCDmNq2Zg+O+YrJ+rLDvIDnlOR7b+NMcDxbAXutphejq2S
Ixh0kSk+JsDrg+TP+k/Thu+mEzzHB6Wq3fEYo7gYJhEXRvtC/1UmBamPEFE1IqDlCRVzY0SdQ7Zq
JpFlwmTrDKio08Erl4OMVb7z2PhOC7pTj/FGBoyI0Fy2h6gIScK2EhhETRDlwzeL1ZnH2WG93MwJ
Y3z0pj/N+6l9OZjCRkSJPuD0QJQdHOo6NYzHfzJ01OUO+zDeWdHpnCkMgToPTUaFTNFYSfm5CFxY
Y0S3hgpTVp2CFrkUexiBJ3AdvIZuZcG+Gqiqe1RJiKJ2Qe07klBJhVtuk81HyM0yAy7IWUbUmlC9
lkB0hCvcV0fek3f9/ni+WCXDwevAQDYPLzC4beNliEeBt21MsO6Gq6LOPMIj7EPjKNH6mt04NeNZ
TNcJNOTTjdLFoXD2kUEuSeMu6XnIKPWcW2NRF58NuZGx5a3xX4FZGE8jXLh6yDi3+3GxR40lm7sp
9buJ/kzQ4k2puHRKHeS+1hiFqHrKA6vYoEz9anEPQKYIiJ2b1+GIB+e/bkYvKGdTq2X5+xu2PFAZ
Po+h9jWa4OjzxT9Y4GzzEP1m2iKs501DcyH2Y9ibJvbj5TGYJGfZj9dVgE4Ew7C6RdsXJXJ4sfdy
PVixHOdfge4dCjaYkGyC70RIEalB93G44SsAcZZykwaCh5F+ZE36kKPozh/n9G5g8GGa6pUej7aM
BaYZznJ1AiybOE6nBEDIDf5xS4WxknRdxtK7yyv9OU1WQftSg67EA6Raq2Zarz4FQDciM7lrFq8H
LfO/hTOEATJqyTrONVWPvZvo+biyX+JILzwo5wLW9sQkkHb0MRoKBHid8B1G7zll4rQlsrYcwRFW
JtZBe3pGjh/Nmeu6l50JcpePkTWXv5MZBMFk9Ioy9bIIGCd5v8saO2b4C08AOkHAmzyMPi96LfFc
O7wItS5gZlIJuN7CFCCRyChIeKlMGTjT/rxyGYxXuzV+5vxOFQwmRC24gotlC0nvMj/htNENo0ul
f3eRquhCAMrzwch8GhrL/lv5zLIZeJrkU0mw8GusarLCIYqR1rGrPlsQA/bd5SHDtH5Zs24QJ7ps
1oqr4M+mUX8OW9rskU/Wupcu0IueOjR01rr24Jgd02Wlgdbc7Ze6lrLE5mUl2dcisoVslMe742+e
g2OVd2ue8vEt0mpUtycNA01jAGrE4BF7/wwdmAcCT1gl8Vcr99ELgRRiLd0uQww78LuEGQ3bRthR
QH75XAl2XBjOSV13pq7uGAmGY3BC4MC9uZVlG6F+JRHOSAM0XCOZqwzXg/7h3cceqw65c7lwOotK
zPQeVth0HNqMVUAfoRPGrRfXu3IqY+8U5xCc8SSIwJ3Ffwx7Wgamav5IMAr7AJXsv9VGln+t02GL
a5H8V9iIc5505sgoQIN9NSo3F+uzWXQONhs8wBow4YzYvSWmvGedKAL/rEqk+V41fSIvfoXdjRTE
Xjhv1nFPZWtPW3Q+lZejm6QfpVWOuAcQdl+t2FcsyEIGJh0uz0O/XCo0+7czWBP3lSYrdwmB5UXv
mUkJeXnhRXKrt1ORoZPsOZbjIvIONYsxdAp8jm+BhA0F21ZKyGyBv1LeGDOKUevXVCXEEe3ZUW6G
G7xB7rhAUn+VGznvGwGlf417OUE/hRqgUQwSQMRXwmPUuDpio0cZIBTLwvtVUKa0wvi1DOECek/f
VxHrE0m4/7mtf/FwI+cK9D3p56KdcpoSc0FdWcwWrrrgvBn/my8IgpHI3nOAwU3SjWPgwC83DLx3
OtM0WKK24OMbo2u3E++usEJxHT2xxecBEcM03uDUQCJ6caqTU+sBSykDt+4oQWVDWSUliXQtkXLe
gggadZRGwBiCzrpY2KWcxJzkFLRSKyES6YqTUOEoRM7maBREqYbIqVS8hMPxBPwKH0sbQyn+86Yz
nI6pi9QosTEEo1XeI7L1mwICxTM3rS4juesVsQoLKW+g9kT2434spIP4FzGlxSdSz6o1J7mGTpWM
7RlIo5eFbIGTGQRs/bfqusu5IrOJoorno0ex24U/VONg3Uva0W2coAjhJlGM877aPlFXheLlEIl0
yZsqNaon3CmIz+CSYQNnMvfdvqdwZ5kjJ2Jcdn5yVdk5aRrshoedfuC/p4C7Wtz6Dpja12kRajy+
re+qNphY6XD3eB1WeOlBMiAlw96Y6DCcwsoWFHqRu7xYJswMHGTa6XKnZBhEIS8Ja7HCG3cfKgvV
yhhOB8L+WOS0of51XYdt0eRL+9Kb5VZZlI+OI6Z6gCJmWxTRLqXmQ1uGZau9OHR58OElzvodA8Ju
4JegXkcyABcPfGxSzlWYMa2SBqBPLEUhr569H1AMZF6/Ku4XGkfZBhjaXLAjkEc8BWWqn2spMsbM
hY2xTgB1oryT/uelkBEjczr0ricYVtDr8e29g57g2gtEtLWumTIGrNJCzr2CahByxVGcPMDLp81I
+TPm2u0gzsTln6WayU6yRrCj4/1bAv+wLBMaurpapO/i7YhD6xQJ3lbFeSB5jW9/8MaOM2jvy6Mz
R/zyL3MoG/b8XqCIGDwX8r9I9cSZLaqh0c+LGzpBkHFDkCBkec2hmow0GlGCHt8baBa83Fqkirp2
BTJ51RQzCeEEJs1A7ize/5b6OJ07+t7RR7r5LbPsWhO1daPV7C/Nrv7L4f5IZtauKslyAbbJbHCd
p6WYjLEF/qn4bzcvdjYwP3XmTqYjA0y67Um3am/bbby4uYfa5YXEsEi0XfmKIjAhiq8Ub3eSUIz6
EuFM7FuWirgWV/DT9CmYj4QLHNGaVuxK8woNjp8LKqkjAi9+ZDGTwV0vCLDAR9MFe2+U1FOFFjYb
70pwcRYGPK6ckPLSIlfbXKQrcJdzfonY30+rd5D5ONspAgvugN32MtMzyo3B7aR+dzJ7GMaV2hgN
IsV44Q4KCHTwck7mfKRt24VLNVA4rRWQ1VJEZAQyHBcmwpk6FvVRHjtn2v4ZIaW1Yn9MxGybEqVL
2DGBOc1tfiluaqkZtmbDiuTVkIKQv9IzU5R+XXT8Nfs3KkNG/HyB3zFOGe2dkKNkRJCJ5E4KgPol
iVpR2ZKPf4y5zOgJ7++CK+ESOA2JGCA9/762p/raxvrx98xaFNIkjxZqAmUBa+zzNrqMFhm5s3K/
hnUhYvPWs/1oM3uq+iofbuGDQ+0dDjCBBpvYGTV0xUuEqULualcNX50cKGYqBLenzJvjFGY8RC8d
HptR1HX2DNV8mu863XTq/5xyeZqpMuxzP9oCoKp7yNABkyf993lfcZLIx+vkuD7qWXQpsy1aC5rN
TOXGDao/wjiCYZSemncxaqX0yYm+48W3q2IcgKPlZV2h4MbC54mi4y1YdhiuehKiOKoAEQGxBy3s
OICdXGnM5UoZ2fZkZe1xbH5Vri/Ten/asEnFSujo/q3TqWkgIMJl8s7OSCOg0OHPbrqNnV5adYZ8
1kqECOzmR0huNY1wDuRSvX6gWUBQIqHylBiGS14NwHvyK3py/S/xPtBvgD5VFCuCGn6T3xHRkdNB
4LG08O/nlKTPgCdbq53PnDDRIdfILQkbzfSWyAI//cxU8sq8+AuU4sZXPFm9o3992WPNhjMsBH3C
m4i6T670C7eTuencYkiyvAsGLErEmZ4RzVD8PU8FYOBiJE6+j7QF3TuMWxeEMdRcyY6NMwdMH6Il
jYkuabFZbW9d9vtLYTy8nWS9Eg+xAZC1YEVBNH4nNlDs8Av85U5/h2/ZrYp0JxFVNTCAG3NUbEeU
614XODRxktyajiObaFSfskhyK+hLWCsEngdE5VyXn53yiIuBVbckvnNFXeVLYJSn8OaE5fbqtgck
1Nwbo/zYeJZOjCai+ulfzIYmuUyhH37s1lNg3E/92AkjjY5rBmN/FhPU3OfM+MckMaizx+Y2Dzy8
WMWXMoDUVQub5P9j3NfSFYST0CY8TdisvpSoVgy8yVI9Zy6VAWTBJYL9ArOpMspyNy/Y8sFagu3o
GW9xkj9V+6s6BhaXCm0A6tPRbwHZv8el0uKRu9n+/6c37fdgDkBjlkYo1+K0FqVpf7kTY3m9txTE
g0Qm4QaLoHx8WmQTl2FzVvDA8gn9fiMi2kAw5vtMhf+JNDqoTZxHxD0cUTa/vVDvFDwrmFl+39VZ
3sKqaC6f7u7ofGFgKwsJqTH91eFU5dzIURcu0cc8eKGf+cPCf5uW3X+/0TEavLh7zsSIUiJw90YG
CRZDyHk8u8rvzwcWjcXNXc0JF/Tm0YnE+jwZdmWcU+p2O8eVvW+OQ4bwjRlxuQBlOuVqKKK0ZIpf
SZ8hmuI7A/nf1CrvgUXhfb2V9ltrvnKNRUDZgE3f+TIgEA0PbcIeGz8qRrG6ngv3uRME+Lnml/Oa
SoQDnNH3pLSWWL06joOduUkaaGbOJZyCPyFXA5I2jJQYg4eaijIvvc/Nbe+1b4daAbMlbs9MjqCB
l/lmY2xr9R+bDDMubhyaSVxAOrPeEwTzxhM3qjAC2L3+f+1Kj0A8E3wRyiFS8UE+zDNs+QT7DKSV
pQq/7gWlXY61l96CAUhHRuyu9MqMpOtFZi+PrrORZeBBQAuClo7JLJ0TNXGhXkOrw6rzFXqFrnJ5
g5HBTK4quZerpcuy0K115B7ePRAAVSgbrrbtgoNeguppfnthtICrlBr2wZzq0eehOZupT2tYMNV2
pvBTML0hqGpkoeFMCd09EW8XMApGEjqb2+YoNJxBIIfvjTQYfgaYJAfuuJowzw5q9bA1cpJuSC1M
Ii+Yz2pBjSHJdQamAwrjvVn7BctuVijAQ1Pi1zZHevRHjdj9RjVN7ND3Xzkw91YVW2ofSnv721hS
903Gyu/3oa21m4xx+VJ4bAOG4NxxYM2T/MFHP9K/oaUe3q62Wh4s+7FPAxgpKXGRo9qZ0+81Xb1N
0VnWk8MP1hhim0rrO3y50ReaETWUeAsVNIdrr0Vhb+WnVfiXjfFmeL8Eqwq+K4UlEqfQO/pBnJTq
2m4RW23jiBoCg2HPVdmT5lo7yIk6XrLf4ErzCSS9RBBRkJbmuKDJSGZul8dxG/Uah4FTDlhg9eCu
yrc4LDJ7rKWN4LVIDmCaq0VvOKderOD/EdYrvmYjcfajwG1ok6Z3gtNQpuvVDkwdI8eNqYKitWST
vkHNAVq8PbCoDY376w5jw3jVKZmQpyX8q7GW60ww39yVv+vBQ2xNy7JuAlZYLiM6kVdEDTOV8xEE
NxJNGStG3+vP3WfbKgRb8ucH1Bp45gK8fcsgC2SJ/wm6h+ILpH+91IBMeGDnMzhciVirctiGGNA8
FfUCbkYRIwJ7f6h5BFvK99JznjqQ6FE4iagm6JytAWq1sXRY2L9QyeDxcgIsZojPv6QNknZxsLwp
BCfO3bjfWvVqcZHh5tXsnl/ZWNI0RaRDLuVihgQ1vBit4NI/KgYVGqOP83IoPxBQXrvIRlm6I4MB
CpKDWofeq9r79+v/0FiedYrnwvvKqead8ALmsR5/qTDwEgSj9EEtIApy9dLFBDpPD8+LiybB9IxB
t8ULrgw9r1fJl7bmcsqveM72ezQHdXjk1zjiEmFrfB9bNggxMC1oYOTYUqYht5fuYR/+myyFd1dj
6Fj2vS2dkVA0HaVX+yFGZbpGWX87w0p2gA+u5LBRVbBSz79XQLBTsOkXpx3vyKsjsyo25Ubbj2Fo
2wquxMHBwJW7cpLeyPWA9Vhlgdfmrloap1al6WHM8CIfIZILpzDAItQI+FuX9Ug/58mebIsBhpA1
Y1uJKY6xgO4xFmb999CoWIQSht7XiatQIU0rYNL+QFixafvSDobmg4Ox63+AYZgs2/5O9U0m5cKs
b4Y0onGfzcEj33fBnqzV6Rz9RRMZxgrYIPLcsUt1RuEMICu3NqA8W2qURwf1HtjRd2PwMkIEntkA
6vbme0pGJ+4Bd/u1xInX0R9bkts49n6WiwkZ4L6lxztw4VBW9t9rVdm8EIv5lE4A4SF7MzftBQKv
Zn2cwcO0f9oQxVa62NeqfTIt67TQutnhWuF4tXFZM4s/5YhvF3pfc7bl5PRnec4NYWyeHm0DzHT0
mSBzoulGIgFRWkQBpqPxmn1chrFPERDhJjG/c98D+0lc3XtvHchi/Y7cR1GVb/HAwP+0MknnSkqV
33FFQ5joJgu4wynzgJ0PgbjKvzi08Ml6Z6sZLvYPPUJjeDJLoxPnC6xqsLqqj9IbH8C6vCrRlduT
6tZGDgNm2yxW6t80LLVfpGT+cCz6XJ34ikzpHUz+1nZS8uWg+/o+ygjChfXIJcnKyVodRVrKQVpd
C8DCk4JfGEJKmg1QTVHqiRWnMoVHgooqF+wXmu8wPEgwMtnmGXNEPXdwALMZXPPpdazVGanq4nHZ
vMnrUblNJtamljWet/xUSTJhegnpaFx5Kg4fE/w9m+azzPY2HN47dDvTIgq1dXO1ylq88uJy3K8F
QUfvxHsarrWcqJXH4HoMzVQMNM9mtKAzq46/axpu98ptmOyKx8eWRUmpG30929nnwPJMhdpAHbkv
mWERWkxDc4CpKVUYa0Y4r+UQQDMhSJl9sGtkNc6b+mZ+H14sTAdhTMwRUP78x1aSRlhihB7TzMJ7
HZGsmXUVmxRqR0Nd++j4bwLyQXnU4mdAbfJvKWjaqq927PvbvSgTEaNASH5RpPmQu4RWObxSZvB6
AhE9hWBmQEoo5aHZVk7J+rAzflDgxma2fo49otIOBdFkaBPGoY3RwSSAr9rHD3kehDOZ+hoNHN2H
K69u9f1O8pTtxheggu/JawhTm/LxxY84kVehwe1NNf9T5Lh0vzZS/JtMql0Jz79rkpAsJHkAszCu
BdT4i9bUM6o1rHLDnvVgqBP3yfU7SUm1pbiQCbb+TAYBnt5/sxrJbmbq72lGdfZYMIoGREcai4fz
SE4pFhRyt+k7/h/YEp0ubF8Yvrq0NCTdMk96W4yG8Xo/1QRPQTya+I4WPXSCJUV7Dt/ctcv1Hwey
+FhY3qClaOh/2UXsAOn0ta+pbreUsc8ZVlngPFOll4+TMzSNxCTDMxOpH5nJuEkUBLs+82KL2+RI
AvPTuPSvfGosGos4ITnFugeDpHMTqQNGlLh7qFg5ZkDzvR62H24RBlvjurvf9/s9rYJ8JTtNFjf/
N6jIeUg18WIPrTQd49xCVm79hI/PFlz0avehTuYz08UdS9KtzgC5aQ4MpLmJmaven+vrH4tmFeYD
1+e7y2db42ZNkmj9yolipWtiCT+zY6Gw7V01Cg6m+3uBSo64cPExCmUV497NKsrTm5oL9UHA8vtk
ZGeZX/ml8MgPE90qNwEOOkt9/1PZfz7+l9/j1lxX15R/wZ2cxSxUcTqkuZ2fI20aW1ktY7h7DApp
DUOo2s/1MMYLIIJ+a1zbgTJbbAn6NGMLSDPOyezjEkXw3KepMK7BhytVo8herfHc+zQEtG28t2kx
XXG+k3304lnAtgq1lGfJWMiA8hYUlAPBIVQmEHHaLzj+iqaGoR2eMWSrU8u9kubPqvCWy5bk3UY9
IyGrtxCRhwzGxe3xnBOsMnFY9RmDKV5jqp/cV1wI7lT59K6OmKYHaN7l+dksQjDg2HjAQtrA7vEg
CgmRqhE4HWavzaiAmX+ZSZR2HfPMaCQE0YsichEVQCqltEZaJzK7dNqnVLbS9CkFN/kDvr6CmMba
Hk8ViZpCArtbVrPIyDjBS9LDfms7y+qGEa1T2d27yFbIXJw0rRBHEzfB1ARaqGjW48qJXFJrJi7N
j5fMYLUpXctUNIQhMnDfaBAudDfGqkNjHfdIWB6G23PwRlyAatX4KVSsyUDeXbARjDVKhYjVV6jz
61O8Yew4DWh7WQo+NYuGm/6N4pdoEVSSEhDIq+7n/8ScNlXgkg/cQkOm5gVz6iHg+/2/vIoWkqq2
PjhSJMsSkzKAH2qHPAbMxMg/uidY5oeJS11X40+nB6fXqO/VMuEQyFLuejs3EJeyV8xdNDPBVR5J
iUgGqbjvdWpvvjmowX6F2YBHe3ar+/a+hK2po60bqVQ6gWtDQ8DZauzqWmUyfuJYwE7lxhAVVfRD
FL7x1BE/AL1dS3NcEpyl5A6Mttl1ZMCoNQvnt0tj5oGwQJDnmXOXYATdfAV2Wh3rxR5snuf+JUg6
E29S0FtdoT/EzLNQRbAk+QUYt3cphhVJeHidmzvK/GxjZ+XpwfTKGyr4i9yQniVanLZvxdIhDf4H
iEBv+Ay4SLIBSFtNQZAcGmNUvf7kFY587sQF6mqJm7eJMo/LxYizjXYymab5q5HhqgfWmIau0k09
L2W0TpYuEtU5d2qebK+En/afv4BNiRPLJ2BG5KVTskfhQEQKuFlXR6j+9ltAUZ/eh75Yjj2Pr4dm
KMG7ev0WtnwBcw5h7ltyY/yyoKaNny4k0a9VoZVjX8E10RJqGcKQJw4J/49ZukH0vH7HLl7M26kk
uqajZZ0KhVo23SgTV0V0F8tqnI6slUyvGZysdVe4B6aiI/0maojZdkjO5JxU+SMqzFcuDNm5TziO
DH7W9JHgUW023+Aug/F+OGw9x3qzso1T0jaN5bqmytjhG1/6HL+cnwBzzE7ckyuSsOWh4bD4AfdN
aMhuKB5plUuvL3AMr42Q22I7YV0jzljog5GmpxImueVW2qGmbZgnYQ9Ue5ltVMIDvhRjA5B5zJ6R
aTQRsnqXTfJUfFXplQ8vbKdMNgGcb4ImTvSyNbyzWFcjZEJOKcEGYP2foSByXavqZaUd6wY/bEfR
Xg19uqBBoEjTBBRFMICS8YePRfIChNWgxAvXBjPHq8Tzy9h+3QLWMyd3FTtnMDv7IfJu8ToH4jbI
W7W10iJIWjW0/teEdkTVfU/robF/t8Uvahw/iet3Ob2mFcVGb9RmMFpi0YknFg+lHYG5SPhlgYwq
zwl3wc79ypLpEw9AkQWpvwWSmRbY+IKfkl7bv/p1CVpyoF0vxvkuZz5bcgO/lTV4Uu79tj0wqClx
Du5kf9fGTL9ys1aED91g6SPWg9wEvOfwQ8IZGpk5+uA0FtwgXAUwaOtL/ioDJpbrZYl93ninA4+M
A1nOPrRZMByvECoZpRQVUoXT4dJDKs6DAPhmpACEjAuTB84a8AoVDrYWlUpP6J3mNViiEbqkPPWt
tsp40TbeZBnLwmXZQQlH0tS/1UamE4vfjoM9M6E+r0EeK2GK6zCxuEU5NiuftcF/BSWO4lvPWLrx
af5yFsGAFjeNsflZQqAMGhPZpxNrtiKifkKVhIFmXXvurv+HRbg23wm6QFshRoc0aedmXF2H37Xk
rDdYLSzX6J1wuzE2QE3qzpuy+eWCo4WeS0x8+S+KvW8Yt7y+DNz03lq/cpsbz30nqUWqqlCjW1d2
owuw2n9IwmLHoFW2kWAJ7VWhDgoLk5cc5qe7AjnwTosuUAzcsxlAJt0CDwj9+LZOlI7bSaBtCpbr
6jq8Y4TlMbSnGmIYNMQjLYNKRDtGyKs+MSQYOc7ZZFAHPjOPOBwCIvWvWvryTJNMi6ctEZ/tn0YT
U8Xjw+22Qn7Xs5N8070WpqMT3uA5/LKMfderrUHK6AOUa7SaQI/RkuRXOnvFZOavEl0p3LieLSPL
JpUpyzzd29WEAgJIiVePtRHmdEtsM2DU2cciS0QAOTsyAMUVTzp99dRjOzdrkJeRo8CnnRBXuNoJ
J+W2Olbv/M0sEVrbEwO5TBwPwwDzW0t3urkwAeLDOd48Fs9jumpGqtONiB0YSeNLDAXpJnwdauBW
+zmRu9bVYD2hnvbI2lkOj38zinwYVJavB9BDTAKrQf+Kb61b0UZp5N6zLgAhbi6dCf6UnDzh6Uvl
m2lZOf7hjwA5UqaWyvgJYHO4M+PpRyMy193Z1vCzacFritUfK5Ea9IhSO3R6k4FfpmV0+F3wkDHr
lJr1qzVcSheZuWS3ZR1159hS68K5eFdd7sJQV+a6BHGsaqYPrjE6LCmSVV35a9WAZ4Y9uUoxRuov
+gYQ1YUDymasA3+OGLCLdD1hjHStdLHalKKez7zDTiZIJ3zzcZ1EUuF2b2lultg5aWYJ4tdxJZJE
fvygS1amDtJTewmUU+JPN9pGGe85Zdm3UcR/fp113vZGielMYnkOmn2pqb44KusBSLm5VtOcSdhi
3oFUxyYQf0EuPI7AVzfkIjwGSnHsTI/Gm1AhHMMBUOoiCeqiJ8Dg2jBMZSoZ2us0iyQHcK84xb4f
JC6KJdxzy5yKtRpa+ak/fM8EO9lwD2ZM7nlDXb+I8I+/jTvj4G+mmD9ZodjwboauXzuBjORepabZ
f4tEzhv8aD7TdXrxdpGpONaqtnzdomDs24tx8c/McTebGlQBuwltt8XLSwFG2MpbkcluUNdzH8nU
kbQ/a6EPO4bNwGszvDjPSpsx4Qc4eVWhvonzl01JZ7qBoaLoO38lv+sIE/VN9XExmC1f/uURnxbO
WjeXaw3Jxc1Ojsa2++mvOa/oTE2T6eRzoJGRPp7m1ttwxXSr9GsUDjf/4hs6ZU8CeHwGvusG14Jc
LEbHl4PM8Osc49p+jdSUe+9j1MDPpek3fYceFjjqw9HgLaMkVpT9OZnYimBbgd1tPQhIOoihyg+j
bgTZEjjedUpgmkezjLPB3rfe/HUcpNrnRei4jGNs3zE3JC2Qy0uKyZ/fuy6IMvqc98MsnTqfGyFh
W7H62tJwC40eRIrP3PkI6d2cw2HKpF/RfrPj5MAVT2czENemRjm3jaTPxdA3+90LlbA9ZU1kPiHr
aBcLMSW6tmkNUwpuxIhSM4rQGzreHsmYf9/RWRQ4g08TK5oOCd0uYUVdOuTxG227MgXSEFMqzf2u
xyxjYxHwXJz/cOaMIopLWBf/Uo6Or3RWyW2ZsqZwhilky3x9q2nrIW6/V3RZWcyr4hC6QVhfVyom
zW1qooO4UoJWurLBFwY30Ql7XiYsraZDieiEnMFVZALJKR3THiRLpnwnXyykakP0soZCDKhsRhuO
BdCBeqIMP5XxfZn8P+4Sc5AR6X2RKKLUXg5H8IlWfzPPGmD1H+0RsVwp/8nTSOoJsDUKelb6Hrbj
0CmlmkEBVV35Wu8r8l0fTzGqeB35fUS6d9JfDBwjLj2WVR4gbzBIh6mHHlRlbjJbcRljOGg/gX0J
M5mYGMhVuG+QXDQxItUKlqxUiI+HMKWcxZ26yGa5sDHuVgGOaxMTZFmFeLrgp9gG7VnlHVDzGW4v
0oCznMd6h7ezthbR69vhHaaFqukCGZ4BvKu9AGcmXKohijHuWQy8Xkmj9DYeZcXF5YO+bNrSYbB9
Aw+hKvwXouYYKegp9H/JDUwyfKjuAJRFGjrzL8DeHoIFIrqJLhO07q+OATaUvnBm5+O+rpsz4C4b
6uNjl1IiqhJoL5e9Q1joVCYS0MZZbobhrkqpx68M7ksmXKVPy8C1PB5Gw/zZ6i2UjQrV1sHLpoUA
m+Y6up1uFGfo/JCh7bfK5BDnD2IB/ahNsMk2t0KKTmXNoyJLGrsLyQ4gINlxumwRsBu5iO7zTBWe
maOjBIDPX9oWqJaNa13c2FX92O67DsUMkt3Ust6Tv6Y8mzwA/9KgcB/eUZp67GTs2qtDq+rzPuU/
Nl4HW/OBvFB63CR8aV/YO1wrwRHFqaJDDYwMsDQYbMmvbeCrsyvGyoTTYdkex+DCW6fywkIJ3VZL
NNOnzNwAWljsAaSCFDEN+pBOdD+6YQrIat/e0BP2hbJF1VmCBE4VMWuL5j4HxOfOnWVtnFNCGVGl
EbJhWu6QgJXaFk6lHUqbdTfywEYU9gZuP1az9QBOpOePR8lagk+k2pOsUtxIbrd5VBLt9xnIxYC5
L6vs8NDvVuoT1dP71e1sSoiCuUzriuIvOoYcmBMSnt6p+ShqGDGMEx5Z2fhhBfjfEn/6o/6XxTxs
UeVv6VGiPdIIELzNU7MOoosQn5gtrfRuJPi3VbNiaZ+OV5HwQ7tCuQJ6a37skd46MT1vb8/QhGx+
VHlh9odxZFJsZCz/7xGoLFy8OAVLEdVOG2Xso03GeaFSVZGjjB+I9KKXpmkK4t5rCX1RA+6mYK8H
lrjTqqq7n4ezmX9bqXlrjONzSb5Ak1BYS/Si/BX1rvXs8M12HYXqxr8mWYQEnl+sR2nHBT8c548u
XOamQO0kwRS0q/hq6ON0/8n2dZmiZg0gjf4kS8KqnkL0i4pTQP0wNNbBl+3ydOhVfov5QW9XuFbR
p0b+8oDv9UjhFmYqPwuKhuawJV9bWDaBx9lcNnd/bqbcaahPM7r9sX84NYIjB7Yytafe6gKg4vC2
ubVBXVsp5nOB53fEJreW4nYVNNrOUetG2vgPpjVfCAqqvcof+pBnibFEiAg1Hy4tnC1hUdXvB4Rw
E/uhNHcWK4/7sIqoYTiTgWaJNultKPe7rKsJo/DSAVSTiEBTiUAwFejbAxWckWuIWw7fisL+17Nb
QaBYlQylzG3nX1KzqRCP/YDz5KUm8GNdmoZ9sMsKJXWksbJguoh8MqOa5FIVujLWDhMDVJi9ukv2
UcMaDmlDUylMp3qv8oxUjEdhupr8fKXSQidPYUwo/tcfW13YrecTmDpwFRy+Yvqdg1r5Al6fFb7Y
x1eujH2ggI44b3WNKpgzdLWNg2qWxOUBUDnuuFrq9w4xp1lbP3jsuUqpYiFgphXydyie5JbqISh9
XbOzlak5PFu5g5bmihE+9Ht5VPE+90+XgS/Xw1CdH3Q/gQ7HUIPn7xFGsJq5D9J+WvLAaxmftSN7
LTBDSoDvgkPzfHqukSaIcjn3hCwunnBJxiCv1/VKk+uUKW35SRC1br5kKrKtpOdMtM4HlajAc9jx
gBC1eafp3CkZiT1ztUyzWG8CWrpZ4qP2xbKTyKmApy8QwgB1c0oP0dWebdXXiDfpgggBnetZIcKX
b4P2P8iyGhxiPimJbf1Hf3J4amMe61O5sCFxYAPIHkazg8kE+7ELmpK2OLN559jS3hrwDW0+LFUC
FVWbS9Arzz3FDOHoKPJwKHl7WWqcbka2btfQKC/smUU+yJSI1Q5l+aUdDIcqvT41NmjR04YCO6QB
BtEao+oDpdfRq5iYtKx+k2+RHFoJHgYXp93hkiQjSUjbMtZC4xdongL5K3EcI3DQRrc9KqwPumO5
sv8fxNMrGHunkplcjqHjAuqwvdMG0+XQtf8MKYn6odkG1UisPAMh5LsdD/G/Ku+iCYrBZQgn2Jnj
V5Rx3YqqstshRK1Crz39doNtgjqcqrS4696tNbYGRrIkzM+M3zakgjBFkaIQ9lNg4rQxQkJNKpkL
zqvtcc27ENXa68+QL5dQZR5s0rNv5dwHAh5JazAbkU+8od8I4T9/blzTatjf+YU+WZ0kWtFjeF6c
mbb1PdzXa7WUHYsAeTHs3kiJCc+sKfQCM0hceJVQP7OfQirE6T1euhvmFuExUZDlc7NciWAow1jR
TmthVwfvT7i/654AKKINVHM0x3ROIXCYy7ptDUj5mj+XSSt17utmwsq2ctfknCItKEJO8ucaj6DY
yuyXAJ6tvJvt46tbgjkpWfm663jyhthoz9uTEVo7htpxVLD7Eoflz3wxAMIpwpO8on6EhX6Z0P91
Ln1as2fCn7fPeHhrYL7UpTaHqA2fAH+tUTU6sA8YoQkTBm41+wDlg3XzzLPlnpGyFRPAXF1wE6sS
NT1TDAEC8u0WvLOHsg+P/3M1GaULriOvsYq/PGOXJJqpAQoIEWzjGXGFj06njeGNddEAmwtTLa4H
/8YTV1kK0PCOTZVggFeUQFSDmkmztjHxZzzgtH+LIEucen/zm3Zbo9yGZ0BIrUVE4o2UbFf6CPb+
9CQf7ag6xPkwBZjExbioVxdNTMjHOXUl4ls3X5KpMPYD77frBDpPzEvHWk/FBcwYdDYqDNb14lEw
d8QinGxvGeRVG3YOW7BvQlNRu9qzV/KVT9pu0KMcr0NEnu8ZYqTiDbisbsCuAPH2hQVBHPQqREo8
tQcB1wawOBNf7VDdjLbbw5MXgY6mwcb11SefbGvARmnUxNlGpDBKV9C42P0UxL3qUIjb5HFXGrnY
ajDl+7R0rtysPS5A5M6q3Xt+db79E1lsZ44NAcYKSmT3xiuLhqaxnZADWSUKWwmUrAu5JHYqXbst
TjeAEbhwhADwnvpdNGxS/ttdlE6LqOJXJwYfyK/0bWtSKsmACPany3jn1zFGfnP37Q0fdgIFqyrc
jESu//JjfPE/+QjUa+4hJllLSDUPyvZONFx/7Y1H8rhujCrFzVY/m8/2EdTe3NDwunZOHIlQJ3Pj
8F2uZOyU+6Fb7U/MiopHw1wI17p8qLtkKEDDfeCIwQHa53qE5m74I+7M2oaCTaG/N939ZlQyx46G
MOFrmbhWO/bYhcFbBMWhSnWEmBXDOpXrI7oVZWJH8XH/uUPE6+YnNUWNncwwebvYiaEJ9Ghi0C6s
914147RHJsHqUIDj29Pm9zeN0IlbLqJE87wI5Tww9IpZE9qqzpWBrRidHQeizaYbibRp0HzIiPoe
I95+3SLv4hLm8yyGAbhv6MqmuniO+BhUhx0NnbmCa7fwlOjL/2MwCrnYC6qfGsFhoReRBlANmxrw
tRug/nnQPZYHJCx+3cxLdovMHYA324Hf/rPw8iNtwh6UF+a/qrtqK8Q90uPZcPAORtpc2Td9Ge1Z
H/IKrESuT4dBxooWKWb1J0NKxfqYVCmPLf1QmTtRcGtMprKj3xP3aLcnKzNKwCQqhoc3p+x5ChgJ
ekkiS3LK60HgsmSuLHHZdjYBIm+Pg+xUNUfYgQPE4XKV3e3V4fnjVcFvB1lTcop9HzzCgD/s+ZTL
fxngB1oKzDp29QRJZo5ylZ7LmJphRBX4tb3JKqrUN3wTvXJHVB54x2BYaZ3+IhwabJysNXQhIiq9
hE9jJIq3y7y00ZJlf3Ttw6Oe6uETvgBnkUJSGA1k+1ma5oQyZUT586UvEAcJsYMgW1TVPATbPZyx
nrOthhelWeh6E018T5h1paMGThkUy7Kx8KOa8BVOJflp6A4FCuzfyI4mdoRtjEf9yusTgSMHFr/e
t0HoFGNuYN1QtY6QlQoF4RARPY++MRkyoVH/P9pqBX9bH6A+u0FlpSjv//ApqF6SlDHpDdNZHjOi
oNFSi4dK9f3+Gikv0UTGRn7pPPiPWjRQ5ns0GR8BGHeyySldvSTPqqVuga/MXSKrYV9i2KhKI9IZ
jeNvIH2C8pKpV0BFziVRaKqcFKqFcYQrUwN2GLKDJaYF2dGDI+XzPG11Zrcqmn8JJhI7F2jsHjaw
ngo7QLxd10KmTo7TDpfrAxvkJCNbKCrzgRacI8VszvGVATOgCwmAwfyKNcTvXVa/XsukGWjAQBTy
9rlxw7QIzdaruHE4bRk7c1h4xXfbOUdaFr1JDFmqJ9WBTHk8zKbJLdzgVt/Q+EtVNicmZFo2fUlD
6JqpK/ZNkJkd5vwnSLL5nYFJl+BcSJhwku0u4gOHSAt8ncMNTSCzcftGKgQgm1ZTakWyZ77+XfBe
DBIISgeBAak69Vef/MxOlJ9ICp0cN90i5vpLcjT1gAkRSQ8EIIYjgEqOeinj/s3BGGVW/HIKdcej
l2la8actfFi86+dZbwf6Z0a7BJ2iT9RqyToU5ydYSTwoR+WuuN1ihEBhYk8KtAe3/cIqGu6q9lUS
yKMuEu/50PZXT8krVpPMe73abQpeuhefaZ4dQRD0NGH1HGPaaW3cDu4uOxCSD/hzWWf2rlk9y4T/
uWIDVG0EL3dWlpeT008riDezPTAkULLlaLNcSTabzynp8zELVEQsCWSvihhx5lwZNKCtZ8EzsZw2
c+M0xCeaDltcl0G5O3evDTWBL6TgKCTSH4aUacdhtiIEHlqmesL5NvqCjOcKSmP7hp1G/UQjNh8Y
kBnYxWR5u0NsW0Zez+HFgmjdQ7BMsbU4Akxt9MTNeJHn4QanhVppTmyE1w3VYHrNMymsIBOB0Ayv
HR02V6TeiMQFvCVMxx8waExMPlydvDDl3ztaQYInItRwmI0q+LciprWGwgj9+HDWuK8C7kTU79vf
2dD1QPQ53QondGygU3kzEfnzzND9ecqCO36uDHM2DXixA8nd1t/OZWSUqbqpuJoW1+w3dy8YljQZ
EoAthtol4St+FiDQhy8tlxM0rLv0jB4zlgMQI9XAP0BKbUDOAiTTcFrjf9tAXm4aki70TMz5jgxE
wRET+F2/fEE79WN9kx7BjgefNxwa5Rm6hLSVJCmP8NrDmp0cY6WrhGt8riYMX7skNC9kC5doRJDh
+ZfpYgFP/sXrHGdIu9oGuylorABJdP9I8vf7vYsWyqTbWAZAxQhDZfrmD9+cw2dI27BWptxCX4HZ
bi91OSpQstqQNLNWY1j7anE+CxreK8KLmwJB4uusMnda+6+QZJN+H1fYMmn3awrx6wFMJ0mHbRAo
oCzhHLvs4B90DftKH6eMA0cmpm2rWhgvN5sTI4dsku2MhN+K4d6m4/1Moujrcf907A/KD9/oowTn
+xiiY+utstzD34fZ6VpOlql1/h9kHGhcIxcgCY4d/Ga1JewG/1Bt4aB6EARk03LfirCJCvpRXFhn
xD3BMVH9FH9S0M2Fg57L8rWY9c5/aCRqjtCnrZ/y+75hdhDd+gV9ln+Hg0GyB4Dr/jvZo7oGpdD4
69gpPwY70RjNBQdGZRT/0SLquHlR6CPcNk3hn4qbo21xChV8G3Z/wbeysxQCCECsawKP0Z+J+Dt3
WCDWv6EWSyau/ael+isNemnHY9MXrIee0H5QVLkEwVTkxcUenShg1IRyGL7UnrWhd1wtS/hrc6v8
ChIyBszG/Jdg7FpYtU3vXy3onBOoQPlYVC12U/Ir7Yb6NLyjgrrEb6e8bi5c1hDMeM6VQsMAWJ/I
dcfsncUrwRag+VatQ4vR6c3brcf0CJcPNrmOvlEOjlE7KrrHNXK8766i+rlPT19F0Qzb7TJDfASK
pEdyS2ZMuNPhDXuNSfc2tKURZfDGi0eS3M8hJsEn7LI/KL4m1Nd5pCAK3SIaGNqeue2kYrmuW/6J
EW8uWoFGglF4Fu+u95PkQw3dG05OdKTaQMvp+TUeXISWHnfTJxaejG3e2Yv4NKRVLkrSzHFrQSta
ZI4ZSgWZQiBfxowj8AWPleHyMlXTbXVPPsx52ga7Yo1/VIlsViAPiZFQlPWWJCvb979dJtjrlnpj
R1bbKFTVtUFAz04xHVrXVtk6ah1+8AqZoQirBkxNgx7TWvQRDlgsbIUEch8E3mLVta9kBflV24H8
oY5ae390cmCEBJn8YTFzjPLcJmon2DUlL1/LpkdIk0i4qJce2DWybKpGo53Le3ADece7xIfUEAbx
koNvwZEyWRuKKaxxTIIOxzA2KLidyHihEYj0vkeFGFbHBp6DtuSgIKA641Qyuo+7TlnM2g3lDhdX
lZGbx4OuKNHJS0Ab1A5h4I2KADV9gl8i6iS8xND6eLTNQJ0wfXnoqdSA115ggBcJUTEBmExmuEv5
Ihfrp9iEZ+Jh6eKHuqauZXQLNm7CLC2Z5ScpOzY7Sr+hY1rOI6PKBoX561w2qJETY1QlOK0EG0dz
zSaTLba8+4mOKUio9qlEWvO9qAC6KQ4pIW65CfSA8O90wmo3sI1r9gh6rnCkJn6Gz/ZOhwx77AS2
2JOWYoj1rHd6y+oWbiPlNHJfSs1+3gBWv/WCPeJUuTaxoI7YoEGnzV13DcquvDpxQTJOL3KHVuVS
pobeOC8HuXkSDyd5L16vSnjzhWYcyGuhB837Wt/RT4y/zJODilvrLvkM6Cw1BJAmzgvmO2Q3NJEP
dCePcI7g8iomuQwGNBwIn8lshokjTbDYvXz3dVkNBhXKKzmL4FBCupyehdb6NpPLa6mCAn1AhOXj
Zv1EQ3DEuZwOGaPytj1PvoFZ+xIJt6/MkBIq/q9PimCPb2PisbVIXOhX1KqqRrgucvUvfA1sqvhM
CVXRsKcm09NmMEAN9UvQKtTV1F2PgQPOA6GANageySnqF44SJVphBn3ipc2ylC9aRU6krBlXHzWF
sVnEB0KtvCMWbkkpO1jFeP8jfang9BEGfW3rN1jweMlgT5c2ugLE06s7OzYWuxPv5XRtNxAL4x3W
d5Ukrs+jHv/0tRNVZxkN+adlQaHWW3ipBpp+Xsw+oRMA7mioL95mVNXjmb47VBlIuOoZmiEtappI
5OLJ7zizX9SLiLGuyBh39uPkdZKiL1dR5kSgG8T5h2RE3dTaTDLOqC7cd8aeef8avFMnnmBTAup3
UYrX5VHPHLn+y0kQJDbwqiS0VbEZzTM83TfNh6KIuEL2VUh7lwuswxPFxrlcsMuGUmWqBf0iL3r0
Smq0EoNqpQjkmUMt0qGPxFN/4IacSb9scABnFc2OuL3QC2uKGpsaECfSheindK+nwrRH9f0D+w8D
ajNWOq8NKpfriZJCrksr6I/deT6Lrfjc1cuOa+EnOtXBdbxe+KiwavO06L7uQMAKg+jpdQ4MtNg1
0XtsdxR11emfzr1Qp3WgxaQcEZi4dbYMSdotnlvzfyMHq0pDhjY7tQcNlpN4q0Bgl5t42ZwpLzbs
5E8mn/clUgyyjc52yreEDkz+OyYQ5vu6AGGgvQyNXLJAw/L8Jmy2xZYbTzZ12193Q6dEaTxuFnVT
QKaoy9LOpyth8PrROk1WA9ZH1Z5iQL6vc3qVlBKqpuCGO9IngX9FMnV3Zwtpn8+wZy+VF/GI3toC
58OHx8OMJg5QRKlkDM+LV99xuX05sliWXVoOftM3WBx4P7Wy+rxKEnaeeRsXpNbYq+/ca22PDFvg
fnp/UDoufs+TCVZDunEQuHr44P5Zlhfbq2AO1m226VbNE7htyjDkcV2f9KmCZ7JsYaMGd+v91lil
AKDHND5TZU3/a9LjPIkR3jLJ1eVxbxYY/Mm7efPlQiKQStog/XagrGFQ/2KwkVPASP9lhkbHTLS7
IlkSrRl3zF9vBauZThZM3VVSfjrzinHBRI1T0f1ty/E9SB+L1+CS/xGb0X0d/NXWa6s5/1TdfM/y
5fc5sKfvJPVUgWEXhA/38wPGurZz6dQOx0cp07nBg5jUEYfI6HriNGYgm4+CHaUHkq93IWq1HtxV
rNJ+LUJfLfjuv+kfu9ERoiUSoNkJY1HVqF61kEFnlzVCjImZVNO5um8qvkz/dHjvBRfn7IGihyLy
wPkqgnM1EJsNmMX9m0Fi2xx12+usOozEH9jiL5lTgCEjrErh4OxcEszgvBfv0KN5NjlMeutiOSxX
vXjOJLdiDfGptPiSyW0zGEAyh56QNf2Vhw+QSt9KntE8gmxs9EIBKUdBOznMMgNIKzKAYvmXX+s4
Z5N30b9ht+TLS51JS5mVAXpxxiRmjkvdvgeHWDx1pWzfICLarJoTsRIsrQ1zQLEkgQaPC/5PsF00
NX6TXH1iohj0k3n4bfwz3Q5DW48rDJ0dyo+Ry+rrNk2bdMl/oHiTPZ71/rHNAlEjLUXBLKSj2HBA
gfmGFp0JeS3yu8zQ8eXECvTOPuTK5/6mIpfGv/vJyGdfRNqQ07Xzlyg9BJD8tHNNzwJXIcnfOnKt
hd2GpwNh2kIcdlfTgyMcYGfBfGjvZTyyfXtZdwGLbbpCtfSV/H2q/gA8uCEjjcLIKfUDoI7eggdx
Iwy836FALLouM7jrTgwa0VB810RjX8dK/h48MffrO5mGDyR/ISDJOoifS1XwpdrsZ1DZRWS8Npq/
SNs4rf+yd+PfY7/w92LOeigeDoyR6tsCuWx4u5ASLN37/FCaiAOJLtbaGhRRIRkxkdfOtWENX7Wq
dOko8qDCWEv/1Udt9qL3xjyLKydSOlb5DoIe3TcbEsLYCOMlCb0DuEk8t08Ts6FnJChVXG9knYAR
L4vvIEmhTi1M5xfji1haqfOQQ4jbhekhRQmRb6NCwv/UjD1UHgxRBhHEKok8mprVvB2VHw+qQaZM
QWTK6LaUkRhzE5mfKrbEUDSE7uF/DGWPNOaKY5zST/vQIZ35FLZ2HubPy/ojte18/VWGdvObEsmO
8HJNBZZT2TM0rrBOVfQezuwdtf1aLydagBLlykMt1u8fe1GW8ma/5QVJfyxYy4EGOehk6+vi+JJK
b8IJRpswAmDCGwt4yw0e/H5OcbF7dmFnEeHgHuwNNvWiR93DDO6oaun+gyDmPx2fsYegrmElZ6eB
0SibPsVmYdXbO1soSZlGOgDb+fBy5apH/hrQ56gwPe1uD9jR7hc/LbWZP+BWU7ODer8Wq89hCdoA
bPaKH/FlqAHCzfNeN5PRssz9taEP1/xmiCn4cngXOJTiBy4yZeETfxUGoc5epS3c8+iFiyGJR6BV
Q99czYzJcRXEOCTgy7BkHf6VE/+mnjOmySUR8VWRg9rETJrbSzEh+hcaYhK55JUCNhpW1Kj+GdZ7
tH8ZHPBW1OfH/6zfuM0LR3Cg686YFMkIeUDFsq2NqVxKEZ3MXiNldjIMSUpZvVhxqVh7ZBuaXfm0
B3f0aXNRPeo/LMCWC2B/+IDh2rxefFbaRatFIDMFCWTZ7Ze6x1unDbym8sKGgfzk0EsJRFaSx5Pf
FimmPsphkv+sOQa9X7PAthlTiQx7Z3y7zq3GAYXxOmsI6/TujqbKgsn1oK5pY8z6h9nYf2Z8Zv21
rbQ6nxHH8qokMFCHNSbkUsizXU9ilUCFamApQG/K+/0DNjht/5fWQtU+gBtdkwyk+YDD4PnUC6lC
WrMmsiCkX/OACCrPKDPhFI2vvaLenQ7d+jqLLDUwGrV+B1cJd45quHwC9X1WBa0MW2QFdJ8YQxpf
HYznyuTtnI6kB4uDhEDqCgJxXwFQuRBSZnm+p2Rkc4/0ftfa2Ivy9t2m7+WE6PjdI98cTiBkLRGU
IgIv5F3bLWU7C8CRI5OsDlK2uxuCQbjMdcE8O1+H/xbpXsO8OVLoyebrxq2lEzIWo9kh0pb3QcVN
fK2lbXx2ouG7Fm0opAUJ/LljBjhh/A0TffEdcxUntQfPhjR2IakJvhiYWDYGBRYkJ9/b4bL4wd3Y
BNirPtxotdamcaVA5hDn5T6U+3djCOv/X5blsQ6P2G/GsAKEwO1NsYxmEmTgnyqh84C9LLsnzr2i
6kjOPCVTtTHhzATRmgTOcpdET/b5Ga2XVEorznsfCNJf/6RDXE7H4SwIzMsCeS1hYhHfC6//X/6Y
5XDNnyLNiLPpiTT4yvY0tRuVNlvmYuejS/z1vNPYvx24N9fqkOjplrbWs383drAgIZT7bzOLqHL0
UIwpAoF90aQd3fFuLiaS6fh6wtBL8qeuti/iWcGkT+TeLaM4yO1npNEGeRWHgGBSctwVQQDVf2U1
N7BhF1l2VcqXLQgFMBPjRkgQEwZpmXtSpYK7S1muW2PLvYTsFeyeGzTd2oSU5DywXnQ/4FgPbSz5
2K0QDSQA1Mpmw/mE0TJLZxa6dw1NCNJ/e7TbywaMDbNPdUj5tvFFw4pjZd9KTpk+ocjNYJH/6NW6
IQrGDBrCTqLrf2F/42TJQdUE8oS4Vbb25UU9bRJy8RBGX9mFKnY2kx/3mm3L9Hz/0nymDfWmdnlN
o3tbTpHUsHe7Xlwr734ejqqxp7LF3RgidGW3jUtN5QoljcVYp9DZkRCX3QeJu8WyFEGjMJRsItvg
MFYmuQONRAnKToRM0E1+Eo+RAQx9zLfBO95gPasWo/prTdWhrQLH22tzqawVZHaGFQa8ZnSYYMnB
ekml5zSJrhQ0ZH2gtl0PJwUR1dQFrWPVkPcLwKtM3HTrLtsM2ZiznSYxAPpEXKAUuxkx1lV8ddY7
2R7j439d80W0OPM5YxuUS5ItslrNkObBjJGpQ0UK7JKqifmVhy2sWShb7Tp9RaFYVAXNVecZS/BX
29JZ3emjI3UIrEEqMjiDYNjwSEoUa3x807Dw7fR57R8mQnOTUGhgBpIGf0O9P9OBIG4ik/d4MsUE
OSiOuSkwdg0Njsyd2YnNgqWO3wbi3SQnsvDAoVZnQ6SECEbk380KA5ecoo5BkHSxgxfER9Qq5UKp
sm3BK601agNVbwN+ncVBXt3iXxkGV4URWSmxQoYKm9XrK6F9WbM07I5AhOu2/SXAbiwpIMFy7KxM
MBOOv7HxMqANSdTG+TGOmTDJpsB2czHmqD1tamBfKlYw0g2F/E/39sO/Vf4I6gBUi11/dnknRKIw
jOyjE0zKwVqlxeSmCQ5hqDlGXs5eheQYjTfdj9x9O0lIQaU5RYRWL4KF8YN5wAeAByDobT3eCTdw
MYfN4KB/MkYfC2wiQabyO27LoWZk/LZ3FXEggWN+pjpOOzhgb1ebm+4K0UdjCl90BVkha7H3hsaX
OLFFlQvhfOYa4iOGDqaDZaOeqEgFKjVpNg6v1LS/Pp29K/ZeuDx8Nmx2I2VXMIkKGFmGY7lKc9J8
lB3sxgx0VumnTPy/hZLhuwav6aehLcj3PZ/t9er6d96nwJNooA/xH5C2T/fy0hU5H9AR9hQJ82+0
BeS27dPnG88vLBc9JZqZnB/0FwpdfYlREqRqWjF74zdMvS/o20MFuK2Xup8O0sP+D5yjU8fjZpui
X5nRPXyyVQJkyyqHFJsFiNOg+jGuZyx5ZX+5344vAYtipQxZT2c5QqlUP6+j21bcVWZHJCNbMkaW
9qF3I19WkiiqfYnQIhEWUF0iyvRryk3bX4ungX+GE6Z4ZMAcD9hfxGwbNZYNCO89kRowfeQrmIx6
Dy6H9itYI5ztrJyYg5g142AjHVYmz+okkjgs3PU61oqTl6I3zkFLxRLduGjP5iqv/+weqOVKY1Vj
930xcrOMTti4kLo1PyB6wQVHPxOa+dk/LrGanbMi1+YrTEQdyhqVnlnNip7tHJjdTys1BN7quXvi
Q/p5W4e7CRkZ64NtWPSB3oTK9TDyUrMh1grbvt3VIfG0sFc4ePZNiH0xQMa4iX1XnFyr7AejxqBm
Zz6GmrvsXHXydOk4Noo9CoGtlQ0JRzMN6BGxN9UyujJN2H4rdNn7SAGi+Uj8RSpzqF3VxnSDfIPv
FnRKtbvnMSDhlPvFQg4XefqoBpTLGBRV/sbg2RFRoHIPwIVnKRflcCHtD7ns6ivFTw5MyCbb2b4A
U6/F16JkBPL2Yv06lIWvaqZKwTeFU+cws6okTHm61MHtnyMSMG0TaA+Dxl+xrAqsCHhKqRnQCaXp
Lhm9Jj4haICo69UexgyLWGXaQMxc5L8VVUDMUrUoLwES045txWonaRn01oLSTZbxsZIPq0wPAu3d
8cgkc2bzrUo2Pxib7DCrmyRcNBc+IZvykouSj3snWItGgMwSyrpVxN6E5qlG+F2CaBRIPo/Caznw
4zDnGQCn/Xq2siL/KhqzmnxzbmyPn7A9hw+w1J1u+rub6B9z8jpnIm9wZ8uzs2RxjxyphW9lwqBw
cZcTVcrZ1igNX/dFrEmW9fg98/Qr93LXdKwhd+8PuBQoIqRBqw5dSbyX5YxnVLatjkIcrDMdBzLu
E2g2RKLkZVBI5cJuPynxGjygvB9Enrg5MSBJ4Qiq4NrSXdIqMQcs/4IA77bBHhtGXt7T5U+YWFLT
h/jyn4QktlbxzKH9OjAnH7mK/38lrHj50cqEE2WlnvmGyHa4dYoIRYBwAWiAiYGLxJeG27hGEmo/
xXsQwWqbcFS7gAbIvayaKrLdzxrCIcUOhq/7Ug0/piPc2BZ4cPYl+G6Bho1c7p+1FAWpzahvVNoN
8vEDpODnVq0VYoY7Nl8urTdoB9h8Vqm8cutzxmQtoSJm7cVm1WIJ3VQA0DRheDsFvW85ZjTmoSa3
oZ3WHW0AAmlrpATkoUJicBvJbV0XfywdGqKvPfx/Pt5VG4FmC9ucbgE9m6EMsqWvRmJFWDDCxiOi
WbcZJbQT6pmQrERji6aHwf2eaQdCTFhMEtkSk5P6iDR4tt0NNur6WOgHI/tvo6SsEyl5WiZLXuyB
7Pt1EW+PE3jM7fuP6tCc0L1AkNnKL4naZp4rGlgDW1a38iBG/dOLYZqfdw96QO2D1Dzb7XEDLj6J
NykMN7FXWEBaRUQqf4fcNrWlXe0oyiA+hG/llaWKc4vgX0CLuawfc2XtXMM33iz5VKeIxStAgix/
Vg9lcjZBkiU7cLGw9n7EZg4E7nolZkj9RrbH8/JQkDdhuf3I1bjNbp+D3CmDNSd4DuaVxNl4TM0H
egfAcWAnfgnTPmfCtTm1RdLTNxZ3lSS8gWy9ZHEPF8P6HxCOizoOARUQt6HExoxcf6G8oDLqR5As
ZxLhn5XVaadf/xK+YPCWkRyqS0dQfQXCwHQZ+qnEqJkgDq5KpkH7zEwP4hEi1NqcPjs1uXKdJo9Y
/LOBm/+a81z+SFHYOPfTpSXSLj6ve2LyOu0MtleC9vzxIAonE5613+3NMxfSqeooXlrvRei8CKZv
IU6Cjp4N2ntiK1Ey1hi0bAMQCPS/zpVyZTVwdx2MBFYC8exJO/JSmovFSVRsiVeDQ+OV+igRe5ur
tkVTcdW1HWAEWWPCEo8zqKK10cTjY4i+Al7IBmcb9QA1Y+XFOUtwsW8bwNApIZ8xuDg2nG9E34Xd
oIDR7+SkXiI/CTuGWgnueIOuEDMBEodqxL9mXaiR9o70W+YHg+kJOYItO3KwJDrH1q1CuPs8INSE
bCewWLbNe9GC8B+EDjgcU/Fsz8ClhdaIFQYxHJSqUG22vj1SSp+Gttuk33WWO7n8ohlFLMB+zUVu
FqyilmRa2HIp035q5CO8ewjljsl6J7EbiOMdt70nbY/ivOMpXKHt+8rTZGxBu5H1SiIFQEzUlRBq
K3rqM9JCeRjnL/suVPvRUhluSj6XnzatGTLid6IFQVGj4cByqbZWESlehd/ghjwuK8Wa/6ylGSjN
MT/j5nHR0SmMDMdlj8iN2KMlxSn08mpZnfSr/XSJ9f7Bu2QR4M0fqD9voDcguMQhnHzWKz9cpnOK
+rQ+rwa3RY6+zIJ7TjQOAkavHg55R7XIUSHEbtJYBtzZCy84pKbZ5px2w3Me1cGjJOjChUvnMFz/
pZFOBLs8knOnO2tsNwvc9QsLlMZCKsK+5XYqjUe2Z/Ol00hREnx1ND0bQe2u4VhOG7O1sd7u61Sg
CEQyVsDMEZ9/Nru51eZDANJ8D5ZXupS/G8MQsqVgHE6dUveYyIuUAQSvjqCqph1v7ESsTIPkN+Ul
cDCWmcE6iO9rN+MAoLf+W4+QIfvp0QI2HCniWYFe45e591BAeDThfHduh2lEXfr2/05FYwR7AMpX
nTjHEfiYa7wD0hbTN36jsRqY+NhvQec8v94moCKVc53xAqBLPYtWf5WJL9whPy757OivtpRMy0+/
A/I6SYR51EQT9ypNrKh8eyTa0Hj39kc6HP53MuhZt8auRsC7zC0R7u5auh0BGfkrsnFiCwGVCuFj
q2yGZBsVlYfv3SuikpbJndpRNOk6eOd9VLuJCUmzAfF86h0bpUUf+lHNeDkGU3OulcI7UFVNgLaD
IbftH4nCXSIbY/DbADPIiIG4Z8GkKwfe9Hx1OV/rzQf1Dm+y1KvXk9baKf+gJWctSnPh7k8kW9g9
s2nVDL6+EzduWDJk1jS1quzbZImQReapjTNx4jdgme0v6egIlfROGOYs4U6E5cw7OihkBKDNzXPm
l+LYz7SGLnMgWHvIVwY3gdyTLltqCjstMQokep4MIUgsYd2YmEl/7EzksUQjBwDlingVDPQH0gFM
yU8oWQtNZ7PjlsyAn7l5dFkcXz5c9071ZRxscYPQWdSUbjIbatohQi6eZS3/eB2lfoCFIYr4DLd6
evUXy7gUcXmIn98R+bnEJHmnGFhmZ3ZCRQgjsKiwIcZNPMhRNcZbk0aUBS+ZS0r1R7pfcErj49aC
WeerriD7dP6nNwkzKDP5OvXFxoG81N/+wdFoWVGZmRliQYNKZ4yxsjKmLrx3F1OHmMF1NQUC0d49
02zzkPez63UCSs9AK1JrD6GkZkHBcaIAV/D4SBTDljXaVreCIi2xT6mreHCGwQvZsx6XETupDEBC
3jAieyLJTaBsXVSBFJWdwqwBQnK41iQi3AHyYFHScGphg4bc5xvMfL1AzDD59arucNVHmY8v80Ge
+TSV3YEqAqXdHgK9hGj69/9/W6hRtGryBK9AThA1gnAQTK5n/qfMoA2DXbUxS9F4kH0vxnw8aPf1
kMgJbVZeKNlAMLkU+d0c9360UM7kuJQajzGUxwjRYAFOPGRjCYStrDuhKEO0amZjFCME7Y/cLxzV
TDlVCEBQZIaJkMWey6MMp1N3PaDRmVm10yaWQSwQ/6h3xVBWjgoHoJa3+zkRKFLanh8TyhTMvFhX
IQBYBq2vA+HGapd2R+1JdO2VFBK1a5HR+JPFfSHBea4AsE0E71koj5OJ4oXj0678JJI/WtsOcZsh
M4u3HoTOQ65nOtqjKarFOXav15SDMSVGIYnBj+hXgyvWF1OYOHAo2jszfqBL4zPp1ZmBazg49YYw
EWFzrGsdjL5p6sA94Qa4ptBa9aPFyOehSoFmF+yNtzfHdWsu3iUGVV+Y/OFF4jRXZ3ypRYU9sa8d
Q8PnxhLmHNdRRqDpUUfMCYVIXGGBxyHafJ0w2SRgSxutU6UgfTTRs3TQ19gzQ7Zlf2g3PWwwMAHC
bNYGgHaLQjx/khDNaqrYrNVY7/1PQrXnpOO9N0+oI4XJtOg18NRL7uW+J2ZUrAROkJTbq5y2GLvo
3p0tUXuxuSVj2xXlbAUK+lMYe1zy6URyODMhCH6lK45iDv0cOXuViCDAXaNCGOGNWRGcm+UuBJWn
SaQFMUgpjGYEmECY2yRlM9QXGsGeS0c8nSYkAQKjh0VDxEd7GniHqaqcX8GL4WZPmf3eICzkeSJT
5v+BWxoFn8XN8kLjTdtue580A8/0L6RMtsB1hEiUrJ6TdsZi6KVxZkckPtCwErFXDDce2mRobft9
hDHI131+hxp0wUhlk/ADssCnftLGdXcJiKzQ2QjEL/+fQ65EzZNr/LzRIALv5cD+Wjkg9LP3NCB6
By11DLAC32HvYUVxGBnrSl2nSVq4mHqiOoiHOIpl7GUe1DG64F1RceW7AqkLsKwMPbeE2bbS/WaO
zboRBvAfPJBKwaHsL+8S1BK2dNzF5MXYztMk1tnOeycqZ3ZDiDZqb0X/2hoqOkLrcIqUXvoEM2pQ
xm2SQKyJBhVMND4EMYpZXrh0ZHwl0G7t6p9c979Vvcpn6dTjeDrLBpZ5lPK45dVHt5Lz7YtD/V9w
fsUYla7mxGY69VKKH+kQOxuAffdBuCgmwcHPupTNGdb6e7siQJr/N42E/9+8MRkVQZILMSmZbcv9
Q2p7BfEjfztcn9ZpSfKsaARQO/bAh649vWQ9ZisADNNKHAcHuLr4j9GFCy403tsAG2FE+50VQIRQ
uKWl4IwJlY+wF2ieV5da/jzJ3w0jjgjo9pQY105YG3NQVTv94hs+t2D0ma2E0Lrx10xHEPIeqFsH
PM/1AJzSMP0T7SOMgNa7oBZl7cjyHtM5WD6HoHgx8YR6pdr4CLcjtTdK5/YHthMGulsm1/NXvcyW
/RA2PNqG3ntXi/mgF/itFnrWVqEvw3wi0WjDC/7eBeIGxYbt3O6mMeF3NJR4bm5jstMXtNhNM9LW
/tKbNFxMscPQ1EFkhr/vobopIbTxVsfw1S49Ssg/nxPoP9nLJLlsQFzBtxNTOqIPN/Vo03iTKMzF
7YtzGlVUfYCPvYoVo+chs49BbLT13uiRteB/KY0oMSbbMRRrUBbBLZXrmpEa5gBio9RfPSXaQVPa
+zv9m9GCh1pg4XcYCGiojhFrt91a5kP9MVhkXJor9YNpx2xcJF+DfdaFt3WEO5yWqFKkocwLNnp/
alwSdPv+GY9689efGpy4Z4YlAXKOzNp15FpegXclEHaldRpiwYXlDvQm8nVSVy9eMwkMeT4yre/v
RkqweZHNrJn9tAmohx4PjNt5D5JeSy61xBJVPBEMGGdm/R6sUcX0gn9fAW8rowIq6RpkMoHJMnfl
A039dKBFSsrsf7pkNqMd2A2qrsCkzJKZZRxdG3PPNR+MdIWtvfBB2oFHsDFqj9IiEnInZz2FPOe9
eYRMy1ls5AKw8+j73dFAJYK8xD5HuvPwwLbIyNP8/AxNtE8GNFJwpXWZAw6U9RbVZIq6hS8sPC65
8DxSNywyv/o7Eu//JxrmzkytYFk/6KpqxEy8hY1kxgaJ1fTnjvq15Fd+6yesHy314JwF8/HZxMk6
ayB8TJyzu4pMIUvtNFvoLMYtK01eGz5pnitPh+7mCL+8CisDLg3sPZTxp2OjwyrbaNK+5pIi8Sty
2Kvidi/k1GbV8i7lsTvxOH2So3b+B+lMyzjASujycJ8p0lXpUXnokEDdxXU+hFx1SV3+mJ6shsmZ
9HHH33tOe4OkvpGm80iDCiFtSdsScsXMs7tz6SqqCOpNQTWZRx5mEfDGfF+QSjpxhf3vfEs5ZUA8
CI7VEkI7jBkOrzPGAeSbZd57dNhkOR3PwoD0tsiNXKRh9UFjTYRIdV0Us4t2ruSKMAOTOZrqhiRR
2HtJB8B11IeQkJd01wmdek+yMG5LdTz6RbyVI9+qwQpOLr7g5fqeSc1rtQxliHfZnqeWlL83HXyw
vmke73AYSHhq32ag5T0JqeFaDKMgFeb218E8uV0E63AMInhJ1bQdYkGKLRHKVU2BeNwqLMsAnbU/
T3dzZ6IFSRNYYtovQhhNmlv2hSB5PyzVrBGSvG93xgyGsUir2k5cuz5Pck6qayVsXNh8eElzzm6x
24Mn8rhWtTB/+oeZYESv0Lr2X7PSP6BuPZFwMRJiUjxEOxKAuz0p7sWBzc8q2U/80kqJChFwm29p
1yqgGYT2oAkgR1vUF40NvoIIgGFWFjEsRmdl01/E2CR0pYVCa83rQ/3QEypc8FOVQxOgeZLrL2oI
8w3HRCOvV8qi3QVbf1VieTnoufsPbtT6rcUjIN3+HzwsSUeqk+RxSmK1MUX/nQ5Cic1DBTUgJnGr
MM63Wn2d3GnpDZ2WwsFnuLD9sOafcOfUvS6fPYGd0vqZVrxvfwNycDrzAbb56C+GOOa+0B48feLZ
Y76l68HadImJeBbW2ePLBdGq05H8kWHM6Oljmzniiy02nwYYhSTyRN1MKaEnRJsy+0crh9K0bRTi
XHU+XOcTthAa42yiBTUI26r5Y7bS+uCKAD6NU1Bu0ogVPHIR8NeXFYBLUIlTf/1oESG2gRj70yaO
gmZXYJaMHURxqA+9VtGJOFI3uDsqHIWZIpzasc5uHEExqIogtEEzPck5I6b6jmj+RA3B1A5LLOTL
B0ju+QLK4T3Y9orv4J219ItFhlG3yzGHCP8LWtDXNbO5ndaiPgUpGw4PVLsejJNnRz824Vd+eKQb
hdPQLow66tB815hjaOd9s9hVFLkVpoti3pULPoz185tYjfA+ByY9jwr52yUClXAk35TDorxC2dOS
8LN50B6P0HDLaqRY1rf8NkHUclZ7n9N9RlUTk9nQwccZgOGGnPgu6O25zRTgG6eYt7gn1ymLMpLF
sZSxbSh9P1uCioz3f2SsJGm2fXI5RruWqW75kSHJchY2oaBDHVsy5ha7srh9u1kmfhF3nC5jIodu
ADUN7Qgm6FECKKtb/XheGJgKyhqrvjlg2jqhLMiK81qRaD8zHQRolxeUVPjUMRH7dJy7iGIbWonI
AtjGtiNELVGkogifpVRdT0yulnXY8Js+2ESSUPQ21tH/Vt3flhCqpzaZzxF9X/FNbr2/tTeD9UMS
4XWEa5iPIMDJ6rVVQ+NTDC51JLGxfZqcZGnlDCX/3XQxTlFxvXT1XR1BUJqyrAbfIcHValeNam0e
m0PWewFg1jR32wlyjQybNOqDFltvloRjY5nDw5MJ6w25SmzHVCgALz+GayFbYkUCaJOefCegEpAF
xkR7sMG7qrxA8BrjTlnw504KZmP+thlFl1maFW52iqFE6IlgSFpM+Drl0rfu3C3dVi4qkE8iKabv
xsfGaXUt/G2PmoIF9hEj2ZTqKTtyxQYTEZnm30eftXi9Al3z05bsvE3jXAuzmE+rqocgUvxCzT0n
McVNA1nPnb4tpMTLRsYh/athO6Si/k6CbAHQJ7PlbIoNLmByfqIqhMmy75z3QvSvpXi2NILIn3Ig
kZb7uxefhGdD7JRxQSqFJDkZYoBSV4rQOBhEt/+YOd9wFAh1mY4HwQTrHAg4VyyURXmRPE7mb/wq
eeHXwwrRxeSavd1LLc5V6UAmNZvwKl9/4dIkbpAXprSsSGBpsJ02rXvjTM+67O4RVIn8M5Z/mbT+
d4d5yeapD5mpivaql9gfi7d8QEyCnpy9zBtE7/mfVsjdugrT/vtC3NjgDmn6xes5qkwn3k7hZQ6X
0C/Zhyzuh4C8K+zWls4P67bk1BbWp5XaF7kCg7Frrk16skKrYK1FvwtZ+NmMlPuzvXv/2U8D8/AE
9b3yuYyiMsj/tMV4QWtBi5WCYE+7L/UyP/vni+TVmSvlK/83K+em3S8x5WEeDhLVirIMNANvzLgH
G7Sih11mvEHfe7WWHlPLlZGfTRFTzMi2Fh3wP7rT9q7P7YyaOd+SU8AAv2qbC6jQ4391l+hDZBNc
zidXBRZ53sSP2ygRL/vHz4lC6qhsG8dUBgWAlIk11uS02em+H1iYxZFNF/GZCCtSnnLsw6VRujIj
npoKdJoUch+kHUTeDMUKgVVLvOE8zOmADTtv8goXPnBBwZYSox1z59N9fAaHk/a+lWablSF3RSgZ
XtWeO5t9oksh4yd4t4wcJSza1/tjQGVnEIzKCf9bntLSAR0GzlPN9kkV8Uvv9xeWMj3QgIHUbKKs
Zi5fQj5sDjyGnvYjNmzMz1VgS7U35sM/gF+FctfjKotkndcDBRM92XoCg3n0QRYDUIbtiGU+IcvO
LZfO5Ar0rkVpChxsV2EI3PAulMWgFH4ihfcLDMUOhzYafOEHX5Als10/Kq0dzknWvh14ZgSSJ4Ko
M1XJrkw+9GS/EsLTOdbBC1XMn8F1BxwB5kOXoUHXL+/Y7wYi+dNnWuQgVaXn2ULmUQjg8kAYurG1
DO3/2px6Gz6Umc7IMFeZa2McfWyzsm+ZAWoIjIdcOH403tEWtEP5On22utPR8Lciiw4LrRcIu0pH
lfsqdamYJP/mkMe6TrXvS8hxgqGEwcNoClY+e5adcbTe/tF+r+fTf1QqxvOrDbyGLdfLyHaz6Mlj
fS9gL+Lc1kXlJ4EO69BM1oYAUlM6sWbr7Z0d0ryq71JnDwQYyJGRUxBF5t3gKGpsTOFICHE6oHsw
aHsfrOngzsqlofETe8ayclavmSXg+ANXXV/jIjnsNOcoD0p8iSw6vCtu9bDfbjevqaZpU26kxsYW
JNyU4zefLGPtd8sV5yQdV6029RA+3aZM3mMibeudjcL4YztcqYnkmElRTiJca6YMnVnY2p9y3J/c
aThKt1/Ik5jyIJXrAJbLXg1x1T97gXwmsHN68mOXIbS54NySAC6QDbDH4aEdd8O7YB8SY+vkmNo6
DFUTfxpGLNOrCSlxE4W3IQ04OOXIiCvsgdNu2XOI9YHc9OUU4YVEIaHroJUQs79AdfrHcrElLjPx
dPQqToURx3vwhmNJ0vJti7jSenTw/xLp1a+MXD+BPZ4xXGpIs+57bpEBLFp9y5kr2DAnF1Gr9ktd
I5aVGMLE9oyPSQ1VNSXGGnqOaapcMn4a3xdBQkqlGZlc6lmUoeYIoT1VFy27BcwZCyD88ZSQJ7yN
4FFWIbBMRGiDtZ8UltgF8A43/Y4DvvREjQByhBnJ8Sy8psb8Iyr0I1tvcdD9FrDVjlsctokC3A3s
z1XGfdncti1fZmZTbAhKgYchsRbm1q1bu0nh26Pb4Bg6YjCgt9a9V79ES950HaQAnSQ5j+t6hVkc
XeDh6KVIzi+AXVkhb8jMjUevunoQZbg1G0qx9tSkA9mHB5trP4H0axVU5vNuZTLzaHkfhWYwdjDO
+hC+1io4lJjx2Di+s6zAb5Elvf5GGirrEoGn+78fm6nEHeazXhwem6DtDPRzhCY1pNSigTc2nO7h
dSo61zSTaYtp24QXLgIrIusWNKnU2/hthcFKTBw0JCCPes+AB0f46cZMWUjUF53IbY432VEiClqM
ov4uy82hoLO3TY34MgtL8GMgwk8KjSFrgMvXNq2gIVdXoiMQUdrFQin1X4rwu808t+W109i70f58
xYuLebxfN4AlWbfw4ebwu5xizI6FR9+gxk2sPbiiu/RhPaZiQPPSga8WrO5VukFlc62wyRXpp1G+
zkgWDROoDPzLefSf+eyuL9Ts/WhIR6iw/wExcvetxsHb6WP36+Pt0XEModl+txXYbftX8y/ubstQ
kBxU2KRNQ61rd3udeVAieLcQb6Np9B/KRDAW7iNObl5qQ4Bnnw1Ddfa6RkTYMgVvwp8rsX5r9w5P
SuTm1tpiUHxZci9n+cI0o+KskcgH68dP5i9l6lsD06yLtfbnSpP1Ty0vVSdYUIhS8sFV2ByIhGZu
nI9e4GkWJ+mMQ91jeiP2vUaFxeqwLEzBwBB14YKF4T0i55DE9qTjHOh5satsWKy+cR2c+IjwhK+i
IPu2+jjB5GtZS0BVUuHMNV6JA6HlUD8tJ5InozbzcMh3HHbTDNsjXBdDVxlIcpTgkFEXRohHTpx/
b5bxHtM682a3VJdR4y8mIQun/AuoGo2zYW3F5bm+aSqUoEWaIht3vcdqKGl2akyU3nfVoPpTS8eO
pdfLbUsHizgnzMUtu3tmhHgnpeUnLvbmLztSGSDS/WcBzmJemAH3II33dXy3TMRsejueJzC+eY8H
tseer2/SYi9kSOaMjFTnn7OXe1XnUgHXLC26djolWYrM2XsEQruleJPjBlDXwL3YZ/3H2+2gnKIH
vRlb+czm8/8zGYtNjf2YWAqcK+22XnizN4Oq226G7buyEpWi5jMRQ0mmOxY5pxjdcgyof8bkwKBY
jm3bSCKUyMFhph/3+FFbh8N7n/Ya6VMYAn5x+9WWNsGGIu0iJdQHvWjsGQ+3iI61Q2iSMcNgUfa9
BAjvSg1Mi/31KUqpd6JLBr1xC6GNxPzjF16mmuqfP4XJUWc/PKEfwMxuyZGskdI1xjHJNJVX4LWc
Hbv1FV4NqeFS/7RG/XJ40SvdeeuEUWVh+TlG+IfHuOUySEFk3BAfbdzHEwaOw4sxzQmO/vCTKxkl
CR2YtJLiEldUOP8BL4KV77tLam06p2QnNeQ4CO5RC4QOH4XopD/Ty0W8b9HE31/HZx1JFEkjpToX
MGFN2bsBdZPP8EP+Uj9ZjyiX+3TKelwNwGBq0xxl2WUyg61R/vqcSM99wcRhVpcy5px5a/nhjKBh
97ZbsosKOQqLJt+unch1/0nVMVTtP5RYUz3n3t+3Ptc0IUycLnOBpzRd5Rrot/y/OtX83wQqNMfe
BR97Y0tpYW6L8H0SD2y1cabocR9gzp57yrdSfbWuoc2btOL6McNR/JnyqTe17cBY6JmOu8X44s3Y
NEGJehFXF2BSZvlOXdLXpdI1Z7X+f3E6TkLPvvR9X7vy9OgJHemw0+VY3NQGN0P9j8mJj9ItEnas
1rI75gQrPzn0Z0mGRYb+I75xUd+4M/3U0HHz6x1f8I6GTVqEFIzPH1d4+F7E2XiowgdVlVpVZUVc
PsqCQ5WTqoeMGxwj7cplhfYGmwY7JnHl/C8nqwktXbRKVGRtG3l2BoKXEB6vVpnqR3ioJqwglmMu
RHrLVWiBVAV6faVFMjjvWTtgm6CCSh3ieGPMzv9ME5Ji7UNp5aQnpNddc1kGYc830Lm8HNLOLlb0
dVpmnVjOfomPAaPUu5hcgqJyaoEHWjELR39HWQCeFE0WijGX0FLQgFhviT7KsnM8iV6p+zY20XI8
LFvFyauq+3WcxMnETG46tNQ2sJPWIoBz+D+v0nibYSvnCEOzfaKSTrQ6MVNZFJFUzcVf3yctE3aL
mHqJUuLxiLj5TMRldvy6rD6jNupdOpmF7p4TOlX+EnDMvMEm2QiawLKFtfnq6OGBdGDqlzHwe4r8
EvrdyG5AILSWAFWXEgN019pIa82OXxU8NqEL5AXz+VyzPMWVOpu0LWND69TXtgqlda8/pmSLho1k
ErEK6Wy0zXIZGpEt5DU/bitPFxY4WsxCDgf0gPSbf9E9nGUI+AL55mF8pXfJJKC9iOP0VKM+HhAm
+xFb/cDiA/GHamgPKpW1Bi3WX0F8pIy3h5+P2yXC/cbEl+Y6yjjQVI2Kp06ZX/L7nFKAb8KoRIOb
KEJ+ymWwctzVuQin+PS2e4wpGKqNaS/AyR1OFSX3AjhbXXon+MFaA7hXNo7ppp01c2DMWx1h0l9J
WdkxLGgEJzYpSsfQuOv8STZIXLrczl1Bw4POGOq6HItnhYenc+MoMKpXU9p813n9HKW2G5AFCppM
6UJNdUyKsXXR4nOK51PaCgcHwXNBYsOys9fv/KN5QziNI9n/yF2NjpnXaHc3cViMq6mZUnT4aFcD
BFOx5kD7zgGZHyZQ/9t2QCTpxtLRgHlran4KXqwJGgNM/z9HH3Dvo4fThb0mYhiekic/iAcDeHMZ
YHfPzDbwASjXBH9NBgyi36176QQ64voe2ziJAeY/ZYjLRt8uX0EwK86r7LyyDyyJ4Hs+awk1UEcj
abDOwOjSS6TN9WYBl/cFWXntFCeblO6CRMsbW5+QgDik96JYVgj4z87DMO0W5Vse98DH5bhOf/gG
FSmBqZTBCuhUnvENFmb1ma5CLSlp9/k59n75AfmJ4W7Gq0Rhv0r6ztOSZKtTD81f7V3eE15cAccQ
ayRC3ueRedTjCzn88tbMH5V4iB4bmBPRPk52+1hEJN6X+kapMKHlfKzKHRhBfj+v73fnJVyLFBaZ
vyiMXtqaQzehNSfzPbltqOPy4P+h/JKKjJ7VKLZIXz9iBUgcGro/swbybyzWY/lyE7IlQoW5TuEF
t7CcGoX8MMMaoXw7RIA5rZsqjzDtQ+uFwthcTqmez4IXEdd7gXy0Hz+i+/+MJLJCtQqWJeL1KKUI
z6VhFMRVcVEX2x46mbNvNStino+ByQO21ySZcpTvNWZ0w9eaEn8YR0txo123J5I1XRUyJA33r7jm
hGX3IJbP8jd7egjaffqJgWc2bBdwICuob3PWJwHZsGTiKatw8fQWdtK92ngNnDyN4aTRTMG01b6M
+hVlGW0jhkxxU5jqCaisgawIY4OIaaLVQueVwMzquHCdwUA5S59Z6bAPCt60bDMnWuej6p6anu4T
Gay25z1SMxhpvC7j7BWuWvoVEpKRruWVJaa+ln2JQ7gx+TEJDPPP0menY7GxSYh7+Pj6HfInXbn5
HsYWmosi3WA2obQtZ2rBEhRqTgo4keZ/gXgAi+wLTneDb26LlJAIwu9hzbTwT2bFYUAopzjEI+wp
g9w3oktQzVzrhQvMJp5OmabmWH59ekm1qTTY8zYq030m/26JcF90kgKIxIRSW+dYe5Q1XAXBWpUT
ASBz0qdj6QtCL1w2Lu6rT25c4sIBydthY+gLvTNBF2Cnw174lLfNnSVCwyH096Omg/jEYyvxWpmy
H8HUdeuRELHfMUOCCWJj7bqItCFxryfY+c9C6ZYqseNIkwXplIGAgTWuXqnj4eU4UBe83Z3vc+zM
oJzi4iuHtSD22cTbgyc6CvIwh+dfua63ATDKJjVOAtpMSN/VUF77g6w4trgzi6aMCiVPT7+bRfUx
xUC5/qunyHzjNjx6J21+mTC8PVGslsl76fLDUnhyNz1qggLgBvA81Kir/jSc5Kj3L/4DljHI64gg
ISdQ/9d5F9pJZ95XUjBOV3jVwLD/y1GbSagRFbjRxF5GDtF3DAlDzjdLa8Muhl9c72mLMQ36Vv7Q
jye14VyZCmpi+HEcJ5rCOu4luZ5frcidA4UuIx7e6tUWRHOWAzKZ7Zw4mMbr9nvfH6Yg2uicMlzW
y6xgIAyhqThcNU10e8c64dv/XpHsf3rBvJStYtuGRJQdem2aqjoYoZkGZFYV2bp05q+SCJ7pdbEj
TtICRDGcjfIPYA7U1lYfrdUNQhSQ27hVzijor2pLZCj9IyilX+I01MYInKpUDbGtxEKTM0CJ2Vkb
DZPhkkEmgVkkSdxs881B5EUv8fnCliWlAfUek6FexG+4IPPcn/W+PqukbDjW2w9HRIl3PkJG9gkG
Gxq9UZSfjEYFs0Pv6uxp+J0WOtB/r4IEV+jf20MkarP2iTqAnXeJwn2jCUZjCz9Bw+virUQv//2f
LNcHnTQD2qU0LWcmqx80ArJV9pYYHC6lEmcm+cKcmwX3/Ow3NGjHWFLSz8Xhd5MfAyWEcy7cCTi6
2zEuG9WLJtZPfT7BqRiJLWCdI9g8omyUkrt/cArZeiyW1i/a8TV0lGJb0gTeg0Kf2nJxLm87ULx+
kvUdrwtNW6bqUna3ZDAv4QzNL3VVRWd//KbJWwzBVDr5eReay/USj5EOLnz56J07gC2IKsvUY7qS
oyHo9hRvY+Xx/bHIObTEv+xiMCMxMVitWrbrioJ+/bJOnrwirELKw2A/di9Oi5CvyL8SpwDMP41W
uy87uzAqQApGjuQsVTj462P6BVSSKgujmKchlf2UiqdY/ASbvvV5sOXbGMpRSzZBPvC0mMpRaf9f
pOEskAgjRxgvV3+oPjpdCoIpViV1KAvdg5S+LNrBEJuzYXjfUg1ZvgsJQbCcMDiPlHNCzxB/b9aR
Jqn/wwWUefaC3y33HE9oafcKqrXP+MQsJi/z4P9Pq7bz9NKkQIBRUjiDY+QH2oxJI06nrNfP1E8D
Lgz8kutmZtUNU4zvy0psXacCduSlBv0m5AwW6Vv2lUfR0d3xLCLD+i7STukSjVHmXVlFyBUVjdjP
hFj/LwK1NIYCYuPSiWkwvopGNjhGuZMiaIWhThl4Pu/0TFUzulhR4JuOugDtKt3CZSexmsAwD+AK
n3H7xt0FgskIo7UqODcQvPZDZKvQbhaMHndSomqitRECtM4hZPWhpApnppB+gUsd5xUjHOcGO7y/
WyT7GTs9w5juR2bii59xQIQUpv3RSqLk5aD/8k/FUYjXEzzN/HF3W4L4j8ixQWlsvlY/q0+TUMfz
ElJvLfgrovh0Ozx4LV3GIMXE2enoFdur/4VAg5TkJkTIr0OYOwb/weDfz6YDGuUGEPBAKSvc0sPX
Vr0GUV+fmSkGIzyF4HkNSxvn+CdVAr5vxwzC/76akD2WlOhDAZudBh1AIiQ+I3DzeLhvYJ+zU1AB
XmpIoP+8j6eslwvCeVxKsQZ0V7cqKKKCNiIrNA9kklCHda8gS0RZ0Jm2uyAIxVIi2QvKGr6Jozzn
tDU706CIFKn0zYAUwxt30HwHUE1Tj/XnrTY/Bq09l1egcgdP8vGfLlXDFneS94rCOA8vaSEoqZ9Z
7vf4zqJB3VLmLwKWx8yhx8o4pov+x2SmHtW8mZAIo0Gts1ZNlNW2eZOYdqO26CfDM6FjNiU5sS8z
JlkoHFxltPvLJ11gCo6CpWhAeGo2K6vPE+a9kXusqsHiD9hKFnx8Rsmn8+Jh9jh/I+cHc6VDNUCc
C6mCzPEQj+OJkuewzYS7k8T+Ls+TatHqg+Hsp5Ab4x45/WaBCT7g8YSXXSC5RVZYLi0hNhP7YX7B
CfCnnK10NbMx8+GfBQWnX2FjxP8wHq5xXr4toNd/+Px48l40QSdidksjVC4m+1+Xk6oVbUuoZ8Nw
KDCjDFvpZDe9k+QTmWTDnNzwSiDWIjMASDmG7/ZbBD2qrKg/8KLbizdHO3OipOTDM6Jk1OlLEkqH
0o0EXHO1Kb1LEDRyaVMygoFQk8+9Dq9HeUWDRS+YNHZuvyZtFOMCP2dFASaGNejmt17WA1M+rSiG
7JfW7eT8yc4Zw0H5U6vW2GOl1s+bCT8wyHhKQhcBn6gb+aqV2+zOUVA/eqMFHvpICZ4oFHJboq+i
rUhrP5MyWi2iI4fQiFE0QE7HEKfrVpL0FQVTpThsnHHDjj6f9I78aBqFwcPP2XsBCal3oSc8TJ0g
bNo4q7bSb504X++BDb4KJILcAOXLBLbhO2QWC+5kKTPXBO5iWTif0vQWuy8/meRzRi6XviYx0L66
anw5Kmsek7AYUq3iWNLdnQxazSb9dtYkoKrzv6mtmzLUo7DIRlOf/AkubU43P/PnSWj2RelZk8Dk
bMY/Q19XJAt/xhd+QoDaQKYCXMeWG0B4B5XJCGoZMKzQ7iEdgZhskgk0s7LFKnLnORnCo6NI8G8O
U6mW4c4ZCf2YdKWb+XGQYtnLp+ny4lyoGDveaeFWaM971WsjIVnsG7VMqcsbd9OtwVC1+eVt52Od
GnGciys++foLkP1NTTcagRw6+eMYmAo+fLFmGBUBk9kGmHZpg12WZQL+n+am4Eul1SzF+WI2wf9O
JWl2YuhGsCUnmY0BmPVZRiN3bcxBzfelXThBe2RJHDRA+XlfEpQIPC84ObeK9R34ws9wkhHGVnbb
uzw7gXGUsnSbXgLAv0jUh8aiVLjOvpACyRcUC79dTu8KBH7RgFolo217/6/rPxTssYOrXiQY1Cz2
hWaCsL+DZ06WtYB01szsYJ76GJDT7ymu0x5lVwIOFoIB+IekMqWG89wEHjz6dvNCLqKLlJp/2Nlu
Qf5cOh+//Io8tpWwkj21f7wbKhgQVEqmVn8y5aOm3FXUKbzBWegAcPOAXkyoi36FXhlzaykBLMI3
g9N8uFmKm3DE5YjUfD1mnkMyeStg/zJKcLS9Dg86xVFKKx/MAwlSfAWCx3Ls4jdP5NQSXPUXW2gA
2vZm5MNJNrk3b2ZVV+nGK0SlH3v0b3wVsZMgYv1tgBA5ZPwOtGWYYE3FShTGqgiHjZlztznrTI+4
t6dj2e+3GX1tA5m/k1f6rfq/+pyIm5QFGiUb5WLC2a7x50mkQEkABUaiWJF1UrThLS5/0tBbquAW
8Cuqho/OetXd5x+kWdv5kyR+YQ7RSt5X5gDQzytXYYN5JY1WU5z0aRJmHue3lqG0Bq78f4Hm16BF
ubBuRZBQmiuHIHJNB2CEqPpVQhWbzJrmOTh7AxlqFQDcx+Ratpjxhbl++9yoqmrO4mEgrRMshhjL
op8mJAd653wuhbG33acSq+4ppOiNhVd52SSsCQv2xTqJ5TrsZY9ZGE8cUDwKWvWV6hK1TMHn34GO
xx05XafY1jaN0EoNdN8qm32CGiW4LvVNUiNLJfZr0+bIzT3zVkxqf4X0fXc5H/t+2LtPkoZ6EmYu
5k5tux/HrZWqLxw/xSUn8JB5ikWoMfRElJf2jvI7TnJ8tBSJ02rIJLTy+Tr90g5doZb/MrAeEiJt
IFaeUKgEJcxZbwoa0p/O/Qrf8/vI57VAw9YHSX5P/jVTru0jnrBH9hGNXxVDO15hQGzQ01W0/P6M
tvzSobzvruJUw+h23Yb35EVVZZQkjjKDfF6oK1Dh9KfgBWMqHo0xbDy1Wjnfa0DiIaU1aLU/JK5w
0VFBoxYyQeggvnXAGQ50+P2ixaJgJh3pn9gZpNuqJKtVXMbwJQSFtj/rUrxfe7XlgYstN8oUVT4b
lo8T2hYUHcsKii+pgZezbr19qCnr3ybRvYQbGBO3ClY+dLv0knaGoPhALSdXAIy4UeWYgjINFWKL
TE3XI3qh/aCGkWBRBP+bxtBq0HqL4uIq4Y6BUepzx9cz7JVeEU4cn3LWxqGIff1c7L94ZKGf6uFm
9wgLyU+M7znmKlKcogvhFQvnbU8Ij7bGKZ6MUlaMk2kNe3hDXADWUMhDkgELeo2Gukj26ALcIHR8
Gtx7LYiiq9Zxzeq8UlMxck/xdZAIqacwyHWOJ9uU13ku3LO42KeprLZUk4wh+MTrJmo//178tblB
YJ3MnE2tpnkKWS9IofU/ycWTqPPW8TeF3oqZOw2GN24FKqVissAGzkCpJRmCP7voKzGcQ/AqA4Yy
5IxnPdWt/aKr1htR67qWfhHWrmWwuU+fI2bSCUlA1DgLkvR+TxVrm862ur/cmXhvIdbRqUWqGNbt
Gn8sb16wX1H49aLZczWx4rqzG0f4vsfDUTkH9f2E2ZpmAunMj+uH+i7gFbgsfFqFAm8DMePqbJr9
ucTSqjOROPEEhbx6UXEcWaAiYSg7+va08nTeX0OxexCBZbehzOBMm6p68cBOxRMR2WGcllfwe6BR
xmv38VgX4aNvIbL70Gambg3NQvTjLaS9I/slS3TEgKmKcD12tyFAnZYnbiZR6AkPZSmAQ56zQhwg
L/SqNB0tzxM9rgUsmvSQLN9dgoh8mdKDOoZPdVXDOC8GkhEjl1L9NmCgHXDQLZBE/OdsAL6hhgM4
I6/aMyvft2OTZahydLixY/l21JxvQf9yNZcdoI6cFGcnz0RbIYoxuBnLJDn0gjtjU7jHwqwcybIs
KaA7NxvB2bScV5/bL7kSNmtbgkrO9PLz5HS37v5UAwJL5cpswnY6kN7LbeK0I3/2ODyNzeDBHU3k
+XZPvA7frMwfpgBT3skwFSPmFwhhGRcBg9ruGYl8ex6xjiVbO7G3TdxlINxyLgqMalph8d0kckFw
6IC6WbWwGtIMGhba50T76A6eN5aB3qfTAkxnFVbH+hq/l15m63gYYSdlPeiWGvgfnT3iFd4Bl7Ke
KcjPv1AR0EnrvYVhq6I0fzKMzzBaHedrDBYNo2f7kmoj47ohSBEEILLVldIGoA5LFMkFgNgf4+zx
9/eV4UHPhJV4TEOYe4vQ+wuqJWxmFdk32XlW3ude1v4x+1QNjV2EWPGzKW4kv7h7l2Zuy0QgyMX/
Iah9EHVPJqqIPwdADKVh1231ZqxP11SMvdnK/WgVoNeujItv+Qdr3jnL8VB0VBlpXEdsC34BgryA
cMhB2UHsPNC0wg3g9EyFLsnhP4AQ58kpotanct2HDESFkTdIzsD9BHx7d4LjVvBCXFtcr4qhnc5a
WB23uPeiRupkHej++OaEyiPFOJenUdFh/glbcrFhqhKqCRSbEozzfDKbrWkVP6xxuy7DLVBAeQ2+
NXZWGTrDNpWlgvylKZJOgOmaR16K7ydJFcyP8ga2ujOJMXrIaASvbWJPbPjHSVa1N49yzZk5ndlY
f+zmTNUJRzwZCAsqI7pg/ty6PDisyATOcZgA0br/oNgcG+Ed3Lo6mpoW8YFfhdpEFQz1ptX7GVLK
J/SUxcu3uuCEgCq5NJvO7R2/8da/j9jNZ4h6CrR+xUY3dYod/R+aRcdAqdlRzfDWRvyaWMPyhFKx
4Me+sbWes1bfwIPMpJZBRqIfdMJjZzxhDFrEaE1DjBDdOq1XajfRrPb30QAAWkP4OFcqCCIAvrzD
PSQCRfCUilparTgNRh8RI67ZZb+FtuXThQkCC15eFkWJvMU7WxnP6896qx+LLEUWuE4UBpU0zwV3
N9+13J6j6SImjr6EiKLcdCiPqo0WJqfk/H+kTWWc0OT16N4iUVXfKC2m9n+PZlev3rp/HCPBaDLM
8hXqA4cvA243uUUgH1b+QNfO/m0Mt9c7Gub9GMy1apRNGuwZMOD81wv1SSTJZQG/TWM+MRHglsOv
0e73ZzAcWrTICKDQ5n01HV66eujyKepYb4zXeI6F0ZlsWSbLEDmp2M2AvbL+KjmWr6rdfrb5mwKT
X5osYBzjbD2T/rS13ryouZDioes5cjXGrJXFpB7Ydf2mmUm/PF7o7urkTHP36uwFFbaQ6//3JfuJ
Hty3v65IVef10Y6jt2jUPSOwN0OdAIa//DyX4FGwM5oPpy8p2Dmu9hUEYXZV69iSEvESO5NlNZsK
ZTOXjowqBzhtzXjxFONFaGCdoz1yoKtcOW/e5wg+xNO73bzHwznGjdqVUKah6bFzP4zS9PO/GDp3
a0KPsNnFhLZLGnwso6I/cxf9cIUiTmTGgxVND5GxcC9zhb1iHtwH067eifX7fInMqYq+5Eb4KLnP
N1KDB0CZTpHdEH5dTKZ1icjplgu0gJGadjrjFTSvo2yjR/lzcYJYuZzeJDcSRgjLzBMfkndPhhL0
86XgzJEXgH44TPjvBiRV/7jn5CSMzgrRpK2zxQdp08s6A+mQiXz3COlAC+MW6OeBQMGnx1hQRh8I
g/QszDPNzrJuEXdfIb8B5v104i85gNXJsFQbGMCwt9F6DEeN4eQ8h4xft2ld4jIX43PgiK/j1l8j
C+8YhituoSj7E8WMZRvTvUGvf1QG5SG2XK9Cy4rF5fjQqeOARwC5VTAf6BpVy3e7u5L38ErCz1Yy
WwDpdgE6/Ik/p4PdBteKuDDZqtrYxOa63DwYEU/P738x4hPvfrDC+4oojP0QH9kwpyXyY3oLIZCE
0Bq4+n5XK9F6oVGdq/Gw69ajpxcU4mnTGXFnNRktHcwGNnkAbbbP25agPehY1bwkOW+7E/CKFlSY
kAeTANoX17H0TE0tM9vk+slhDIGqFwkf1XusLp+VMscK5B89S+Oh21UC28l3venJtTvFbXEIeVVJ
kdx/KUsTSJF3qSKJy7gH3HdoDLqguEZu7o9eM5sQ78YhEv6s+G0DWjn+27e+I9KZgTMoO2okMXbZ
om49VsShr18NOQF4VW7eH3ycSE/39AqEj77LhYSlM9NOklE/H2kNAQ+TqDhJS4PHf3L1i7dPf1Jq
p4vA672Ej/ohpzMgK0tXxP5se7MgBEPNVmSxXZHwbpSR1Ph5LxGxPf+fUo30z2f1ZGovuhuP1xwd
o0VKklg98SY4flmfaLxACUmnIGgBYAMTGyYMlFRGZe1zcljgQ1vu5W/fRNMJIYvIQW6yz8B5ayV9
mGY9ojMAr1eUBlH3wtCqatREaPmI8ovxLusX99SMNWGIatzlw7+jSQFZEV+3BVmeN+cmh8tSBwMs
6I5gVoBsoE0XY/vVQBeLXy/mA4xBMnLnUPZ+uailPMFQQt8hwzC8FtgENei7/pK1WpJ9EaxEkNkI
KepvBatFycjItCjo/HV3Tyzc9ff+P+FVKhbyMuJYtN1JndHD9BeVKqqR9/SWzib/LeBHENz9JsNf
uRZWk0awdqpIlty8lmayphs6jipHUgM39Lg9Us97LYvPk2hwCyX2HPGxCi8bgNCTL7dGuYMpRnvm
RIqs1MHbBoYGcYhJE2tddJ4fMOpMYa/3v4cg0s5KU5RxLJqmWHvh3MZOoEusOB4qnAjtL6np5CX7
iu7caZ84XB8iZRBwJUCqoVuN+Aqg2IK9t/sabrcpe43CFheLN6V0dJwf25hvc7weTYbtxCYW16xa
b3cppoiIEK9l5G2gclPfI8bqX3mH1eOg9ycAdlchbML4A4dIXf/kidMC/kC8VcSdbLT9ExqiM+Gj
CeBJWO2KIVVY6+vBMRuCPNnCluje7R45KZ//zaSIRrjb/+8zXSTunKWKsBu2XHsevR3X1UTE6SlA
Qlpl6rVaX+BXi+nXb5e9r7cs++j83nQfCfxeHVzxIcOxzg6Vb7xi5qsRLzgs+Y0Kqy5EHddqfXft
3mX8RCpnDNDcHMjjZKb4sMaHUWyJ7hqWKsS+f3LFePXLApMn8BGAijWeEBIQwrPeX1e7YbgY1hF0
p342pUZhexvQ2N/NCWwZQJ+dzrrvis3Y8zVk6I/cUw9tiBiZyHsBn/YIBMhiCPovHd3fbZkPoFqg
zpnsuiZehvU1Qh3jZnrXC9WAJLGjfwZpNKgHpQZ5vJNea1ANjWtBiAKZBBB4lMxlxkgpkeZ4gEIG
W9lP+sAWsh/uWTWX0N3bF5bCUhYc4kyhEpsRfELoDHa/vYsJmeRdKVCKWKC9xeMm0dyBLGJ0xQ3m
cDEeYLi54X+xNv22heylLCP0jUskjPsuIxrLsbJwalSBmx1wWCgi+JgviuJYFAhOy5hxmFdUtE1O
5h4kB7yGhmqwvMUWWTtF7/uv+ged0M0sHBieRGb6BepW2L5kl/10o80gToVYc5G5V6VX5/MVC8Ci
DzqR7250232QBcWNSbxN9LA9wU+IxxTtNkPJqLzHagIb+q2Xtq8QNw+Bs0tIJ43L3VlKRDRS1vHv
ZAUwiF2wlUQxdmAJOCOl0+Hi1sJSwjgDLEK/kTI9qRTcyWAGtcp7ix3quXOgopH47PeL610Dk4pU
aRfJcl7Ju2m7oLRD+XkkuvmYo9SsJTfIVmLRUgcl+4EZfRaVk8Z5PC3tk9I6lisWt0nvOD3J4cjO
zz5x+lSqMkNkdRGg25tApnHxa7StqqlI2ar/8BWQREHY9ZPN/IB1eCsWX27Pr5SIRZ6UtMc5G1Zm
hv3cJGyL9qD8EMFjXb71+WbjW2d8NVqddRV7wui65Xy8tidpireL7qtLnUYuS2VODHg9in2GTI+W
JsSu6iaMmojTIQCDd5B0Z+uBTT7NehBDh3Z34cUWf8AkAeGMCfzQ/FVGkkenz1ozdOPfaYCw35+t
Dlp0PvNpK+yEVnPTO6sS8QCxiEJxfeT/r/9FhELb8A73ED5jDID296ebQjzY88HuGMKgFfotMCAT
m43fgt9azkynASyKTc+Bedt74hwtdaKCRzRKZXM633FI8orRmhHa9F5F6oz8f4/7e5NNMZZ2FFUl
aDNjzSpAxub1PfwBYD3y5bDpgqowr73+NjgBrhrET8zL+ypsVWuVQFjRIVLtlcG/D0AMzxL/X77E
x237TxP0kpOW1Il0yp/MkIxTqB3nnXkVeMHuikgDiKqbCQxeeMnSVn03j2+zHIgckGfjsMU0yk8P
bPs5tz0a90S8h5o6Rw+JnkYTRp5PSxQ0bl3F0RKba7UOavt0Kn6As8GP/mfEJ2OTkVPsBXCa8kix
J+yRr2+VG6JYRA2QZ466vt//iTzeqMBy8877/NtUeFB6mGdpFWltHA5YoDc2AsGNmyt1veWFECfz
3VG2eLIDKrdeuaGSDAcTFL6lcePBNAchBvHTkqSGnUgK7tvKatt/XYHZt6MQvNC5+OrlatPnKd1T
+cpb/maZ3ZWf3YWpI4JqUku3D3KpliuzDHAt5gKxh/tQAeJzJVsmSxfwDD23HpR0RZiQfYyO+D6y
Hd5G9hMcKBgDoOCk5+u7tSHSaPW6uHZd6KTixKupMhVHKEv6dGHYl2/QPtMROWu1vTj1pLYtog79
xoDde82gt5vsddpyB+Tspz6WS7RyMZEbi2QDVj+SC0auvGiI94z3BiulxvUZwUFQvVIbTSBF8s63
9EMQiH0tLIq1gEzYjaZyeUNyt48EbW/obamFVGqqXcof9xhVnR4L3xLdnM0hHehai07RYk7KAnZ7
ytrRh888yjYQyxBjAR8AFWDZfbBWIIeEgxleKLvAGkINTDuxW/qcYNc8ohW66YCIGMHTxKR8mHj/
Y3+PVj9Fr4kM89cmSHH0760XbCkmrWZqEPmvGCkcejjpFBVDnm3WdEGyP0RmMRUUVQziHtkaGHrY
kB786AYfYYImvm1QhltbC34mEE7Ob11CfIMTUnBvjypN/c9RcnEbiaBtbNjhpyoKHpD0mTjXHfoR
ybE8ghPG9Qca99tAbzrYUa0ZuezfbF6YmFW7TGkP9dS8VlAU1aucieBor00lmie2eeuCLVBsRkE3
4OfiD1RvVnt+aoXDjRgsoU6OdFpljPO43Qd2XushpAaZ0ApDk4DSUNfMXWXYQmLV4mvGdrFrrq7J
/2I5hrm5TXX5HiwJHwYQHYdOWDEtDlqqR2aPS3CReTSM75zfuEcpqd+mE50TKJPNTnn5N2WrPMtg
k6Sf1pikov1ZfTzkf0Z85fSQn8dZh3bEVcTcDVoS0N8DpwoZR/yHC67mJLEaWfM9LUhuXZthyF90
RPi2XTEJ9M7C8EmAvyt5gqnCBJp+f9BX8HvVM1khyZBk32wWuJnmiTJGaW7ShwrLwh6KsWZC2l8T
QA/2vACkJc+mw9mE2SXVN7u55mDUi97hb4Cn+HLa9ywDJHdL0vLf14rLaf9zzBcPtHVr3n1v036+
eNCIuqLWa2MVZ5Uuf5AezH3D2ijY/ZC9iHrKcMhHdFriTPm+sM6rtX4RByUmxWrypJ50Cf09RvG7
sLLzRassG+yq4XDn4mImS3EXdhQqXKFhuwQEpsOpeBiWjcyqYpaeTUHaxDglB92Fr93trTiI4EED
+UXBCu5ILnTZc/TW7HFtMHoGHXZvQiysvtjflrXAU2rQYnx7VMDnUsEGOEZL1NjrGq0CS1eohzMs
1WE26HAUPCZQqlOHD2ngi9QoNbNiVkkAQLOOKGMwfLN76oQizqNqE8FLG9l7nqAVRUfzvZU4Fi9p
YvtO+3Nk6t7xSeSzQAeu+j7atpOX8OSMQ8VUaQ7G8osqRjQlaUCGD6uAMBq11e6IhX+FNBlkx6zG
2KkG/HGQCBDq6aZ9+KAfmo9WLFgIh5TtVX1tkTnWmbV0xn/29fg3q6nDyDwP3rHJvE6WHMqwX6Bh
1MLiRMutMwYmhfvEyKmAkj8SFzHZSGwVqROc+48qoPdYiTNIr7RACbnt7DO8i6qyL0z4w7/vprMx
7i2eAbRMJpeb2l4gQjnw2fanrlG6fhV78l0OWd/44CDjkX1M2NTID5KuYJl1oyzl1/F3nADeo30C
wyGZAO9D70coeNH2eLrwfKQnpEc2X4LpWDH/FCZ9GON3ersq1PgTJFxe7a4Uxono347tL+rmx2ux
Yzup9G/QnDGebZplpanB1CU1HmhJjHIfy9XalGg0ZSl0PlpMj1RgiEaQsG9mTUbPA7RA0DvJpRqP
Ocowdob/dxFaZ/uJSK/BXDSbiNJm2FUj97tKINKQf0LHVs/4/pJFNFAxDKvpl6XpKB5Yr5fveWyl
iV+xBCC5TCvlb9gxdsnwA48iMgVJOBLpSrRY2P2zBhLOJSAZpiEuj9SqL0YECyW+vWiZKSqTVRWo
mfK/xz7NnWQEPNuHdYj4jAyFqvoD+AHS6JuvtAxVwC+q6NBZWjAQl//qMHMsqHr6Ye7cB3xDSndC
ebgMhka5g6OWGCrV0vC7mqOfQrHVfDYI2Lpvwi2XkbuEfRNZpDpmXkCHgmetIhSKF6kmuyNLNFJ6
FbGNpvja0GLQqguBjqubxiSNyBCvqHj81dpyg2UFNlDqHuHY1wMhzFQUxqdsSQOWBc66KO2P+XLY
1BQFYtDfstHVWNqzHW+ngE5g/3haYIKsmqP6r3SEN409V1QY9jj721gsJ9ezVv7MwYlb8IYdI/xc
6rFKu8meBfvqsWTKD7EtbvgsXFiK+wTR+UCsf/DBjxH9N8bOvYBlQNzWMfsX5tbdyQ0dgvDeozuq
IG51CzwSKhTAcrqhsahpYsnXnrwaBo7vcENc4a3FxSJC99Akdad4o/MAHFt2y/96WOe55Xc+fK0h
PbH7fe7sFX877lwgKzFen4wkV9NqAbFaKC1vujgn20PThlPhJDy0RyK7X7PbCDUKBmyE2rk3buUL
U5Jd9fnLTZVYnXbCYaAXMzB2oip1jgX6DzCRp3xELMamGKj9FVD/nZghvBcqKys2ym5lHswGK2sP
dOSDepwtBaK67pryAgw8x8/dS1x/AQHVAfsLc1xEVfQvYzCiTNrdXrPZZr5pf4h1moEOdI7edn4B
ww1nADljCzsQ23pi63KVcF+JESUhKDO9AMfIge6U71ByTdhcSSyjSBEstq93F/atxrB6EZdyHrm9
Yx6L6lWMjQiNoJe3semi6fWJO8G9A+7ZzPvFgqvodHB0sYpYV7/uBhq9fv6UCO50f3x6zyKIS4t/
/p112Hmyk2sE9KqPwYMymrOVtcaUnkoAfOo2BIwCb0HQyeH3iNqJnUbxFR51wohIGizG2/D86mSV
NQQNzCGIebh+XTiR8uMUkVUT1KMi95ITU/2FkARPl+8PWLD7uYOMQvp6o/cggU5QuCFQtZhL5B+W
ogdLLiUTCp6p9KJ89Jc/VDwddYNUItMioMaghIlaLGpVBvSVj20O3RapOw8P49RZM6ixo4ibIX00
SPfG8HdhA0w3yvX/ml+PxeW3hgYIao0D4481fpuYK8BS2uqz73IBC56gIrNJQF1QJuvUutc5c8aw
N4HlkSy62guH6Wthwi8lXJxq0unfbfvlRYxUDsSJ9m2wKtWSsdt9R9TE68MKBSC7jSWTFSgBiygu
LGbmDqDo8M3jBgPLE2u5Q/3K2iJeEaBlp5XH40+JrF9x3Wmz0IOtCZxpGuM1E4iwI9DxeG3KD1qr
dJXPxmiJnXBxmJqD7rIbhawzoAyhB/tEQpCrY4cPpyl85eydAWr6WuFh/SxPj4lZAF+5fMyg0T0D
Fc00g4UKc90fFG2I+LZigD/KM0IBJjuucilNTxLFPM1JUpsPgOX2vO1XM7pSmXH2FcBoH8gGX3rW
iJARLel39E+l2BiiLeBWLI+mDyaUJVAZiRhnPpD/AbsFBAQTlh8mwcSfMvRID2VBbm+5IGKOn7rL
7W4AOmGhpdhRTyAib5sBh1lCeeSns/k6ScfZQF+3uqP+5DCnALQa/cnfmw7sb5+hVrjgJUdeW9x9
pI9sU0aG3M6bGnZ1OWex0gsJQKc75cqSVCpqUhmxi0i4GpDU9qCRZp65Y/yDZ1uqNSG8Ud8dGx8R
+WL9XE+hd/XHE9BMTr9Fe/XqcsikDo/gZ0WrTslTFo5/v2r5bbaVJJBwQYbfigKHSlQNrIXfCeDm
S8DgqgIckeWF/UzVRaNAjZfrEESnm9w9BAnw6/1g1nJSa6/cdPwjlV0qgiQ6YSi0IXS9ABLz/HzT
C8M5PCjaj9ipe6ff/0OG7zlXLEo3FvVFmCAjMPzwdnVkcxDOvpuLIzjgplx+rEinjPoC7J4yB46l
9eAGeU85dN8Z36r5Zm3MynjGH2w3ZpZGEGHYsN9Tym36NyuZFX5/Euon3VEiuo7AS8taiIzHIbYa
Mra/LVOI8rs5r9py/woJx1KGUPKxt4HOhF91AyuHTA9Tj8d1AEv26K3Bk7YKNYT08Wz0PIOB6FEV
Bzu36Snd1Vpd6D4zsrL4PuCXDHfQgemHxWhsrZTK9Fy1fK5vCGHAgKu0pSMVMtNgOAW3c2EHna82
E/FpEzvGt86O+Cy9t7oUmOiBiKMoRuCdCaVMOGzn1hCQvsi5PvuwkClHnEvexqg6gVvPere5zZYp
FOHmCu2mK85m5n8eretHWrA6k4jxljQ5bEu6UZadYBxpAelBcmHIrbEdRH21hQGMPI88Bk3GT1R6
pYI07pH51h09nrUGwNiwXjUPXv21QHRn28L6aKW8YIRS3pUdtAeyWhCybeVJNismxRA5GnHC2QSl
CQPBMZkI6brgAln/LaIvtVbbLMIQtEBRSPf+Jrq7PZSauYStH6Bg+2j7JfOjtuJ1UhS4MZyGIqvi
HbZ8mch4s7W6tLYU3XqSW5kCHOzVmPWiw27TWD5qgAMSsjsq8Woi40lEPvKB4zHOZfEgWauxKK1g
1H1QYM3QZ7TPKAiDwM16aN7zDFK/lDFxlIcVrb+tnS/8TJJ7xLg71l0XZXTugStDR6JTtRgZQjBL
9RgA2nH/UIYUPplTx6LyBheHC0vcUEPDmZc3fj8Eofxrf2FvvKWpKgyUFEA2fGJGpLC4WLIeLEHk
8c7rxWapljs5XPPRXCzJczqlyJq+vPfN1l68paPcrBztjSTeu9hkPyVYsjuWMKLxlNBGk0D4kfGS
is8iGOtMTOxLrvRuU/6rvPT45vABuXehP5jw1BZLfah8GymE7arW+frxln/jn3eW9IrX7bfOAJLi
3XjZ5eqGaRX4ygxZkk81cYSMYhi0T0Fi2acMBV6QJulVM0O3OoQ9kibn/WK8kzIduzaC/JIqnYih
sMdivqUhaiB8zxGxRbz9ZDMzQGH5kLFV1ifFlEYxxkjDfgPGZsVAznnqa8K0hkfEVZ0TM71yKvCU
XvQK2o5G9XYWXfC7PKXOt75f9CHhA/nbezwhAwNKMxnwWOFghIqj4Ux/gcb3vNamTo8XNBnxMAxn
CScu0Dtvr5vx8BSfUk6hn6ZHMF+6lnmSgkZL/v7y5pViPEV0dZh6Xh4T3dUBXmEBW2iN8UxXEtp5
BNk6ZbwNpaH3FVg0yslKJyfrir8GpSSvKZ68TdeElMRcOOON2lN6UqA4XJmHXKEV24aBo3KCpylb
MYhTx2JNZDP8AAb0peYcOdrLqm/iAkx0L5+QXUqGoCQp8Yo01ly8K5DxP/KECXwqiF4+PYZGSat3
0fyKQVBR8fVn8KUx7wxrY1S3aF4QdijFNgZ2eiJoIbTFccFZiCUEVu+WtM/RHJTT8jFXTE5FEDxB
h9/Q/amAFhRIBstAUuEHyBpj6F8Mf6251PQFZnMUqFJOWAQ1Jy7BkokigyGfvrQTlnPysv5h83ok
aUk6yxULooQqzy8FLTJdAyOaLcJaH5dcLjU6JgYSYHWzb2bIt/8v4ypiNs7y43Bq5LGxpt/GnR6t
DeFB5+FmvhaGq6j8OqUPPdQSg5GFEjL7tHWLZUyNFaNkpIwVTgu1kX0E82wjpVCwBk4ydZXgR+8Q
Hx/HN/QVOOfoZH0jIrHouzZ4lBVYU0V4v2ZZzEBa5DssR6VnksArRBab3Tc7IvdNkJ4lFDHLjAgf
fjS/+Nq5sS8x5SJprdWoatzdHtBswHtsT0bg74xqgrtIBK5ZnZAw/1usyBQj+TH3+hIYDGB2pNYr
6H0AUiDcoaOrm/VPurAU4HfrDA4DZlSRtm8QH00rPP3lPlrdz/iQkYgvEqgUTVlq4Hur+B7nc9/z
aDeoCpwjLEaCpUqgJ8EE9NL2npG9qY86Cle1MgkfGPlEtifL8CW33N/6VXDok2f7BVvcex4jn3cY
YrQaUqo56sWYboDO0kCs3e575R5YUPfi3t6JFojf5/CVLqzmV423RaUGHLmRJ86QA2c4YDuhXnxY
PBYdTuf52cMjS1kwgYrOaPCFDlqqruc6+DP2y2Wqty7usuO4oOZC9217teS7HWwMD3MHwF/30VPU
UL3iuEBVFBwrRz+qL9n7JojTy7xBkRMkX60uZuzwNjESyw6KjnkadJoXGe9MQ5Fe+Kn8yX+NEuqj
3nSg/0HEfnsmr8KeFApin39IRrT7013R/j0k63jlLASzr5SzhHxBRoECdxmG6QKxsY9tw2lVWOd0
lEG/TuTjP/PWqcc2zVetBxH4KvzYnn1T4cfUNXUmxM6RfLqxe2NeLwuY2NCENn9wSlPaH7NzlgIt
C1dlz5k09ySQIPfmBV1dHhT78Sr+DGoSjsI5WNQTvsgMjXD1t99hcnhJp6is5bP2IZZ40GDp/5/O
z2FxPjSUMeWgf5mcVcwLRiKxnIf8MDsk0Pvikz4yv51RZ/b0kOxDNOVyk/wrP07us+ZGn/jn4X4V
hMh+FyVAUcoJYPSOQo8js2FvIbtw/CrK8pGOvn+oTjzxzq4/Bd8sU4Qta53qhFGCtX+u+lbcYcFw
CYS4wHZEavPopwUQh3YVJSuNT3MSPjvmi4M+XmcK1W0g9lUri1Pe3LrbVI/y4i3gCKdP+8x8o60X
HPIZDI3Bm9L89UOjZz8ZxCv5REVoxMp8hCMRMg4bpJaSXZts9yx7Mk8k19sNXQYlFyAOrws2X9wi
zhz7wQzL74Z72tRmZktq8nCuctv8uWykAIeUSiTR1G73ICrIbbslVWhNtllsNg3dV2yz4g+Pbc/W
mwGUAMJQ1ELRIdwN6wVFok3XrUI/lzpruejWAKFTyIXl225q64oTZyyXbuYQB6W5kLQULNw0F+IF
FyPsozo6hoDzJDo3VJsEVAPi0aJ2LNrveBfHyuRSw2PlklRU35ih65EU3LifA57XIG9b8FAadv7L
mvhOJKFYFQkLd57q2CbqeDkzZKGzf4Xx9qonTESy+lkHloX1Mm0u3//l0euAzWglzwZFUjbEqXAi
HlCIwqD5kltCJY8UWRcBggWWibYMEHoXK58xsGMizy+hBVZ1cJxpHJ1XSw+wnMCHO0XimnsIXi7G
0PVUdZhbGel5sfqqX5u/hJakccVFmnPvwpq1+/Z6SY5DgQ7jsMCD2KkrwyrdwcQKiIKKB7PGrWxs
Zpn2hBDzlcQbcuRL/h0guL/jP5yY83IlOcg+PEO8XpAZcTDlAbL0j+oVSIHcIKMJZ3wz7/4c62ve
eWLCES8pnUbIOD1DA1l5TdbbhtPU2ctrOZ0ZIEK3TjsFgTjuFDw3k6xN2Y43CHvG0cKwQNzhprKJ
G1jLJAtuUY1CN86yxDeca75lQ3aNJbP5gB90OqtiQS0v5tdCszITCrSc4sQSRl7F/vtfkuCDJ6KT
kA9YqGfGF83D9kcNMOpdLaVKiv9v0LmTB3SOxKKJ3ZZHwQkKtDrSPyLjr+l3a/1J+DdPEds+FOBq
B2aGnlzPiMVwe/dqomJQL5C72EofnmEZrrmOQn519xJKj9mC1T3n/dEvonE2he13BHW5sEJ4SNrm
uAhPf/eYO6yZn2bxo0rD0xskLmbzSrvzgu/zE4cK5mF/YF4zQB7ihJ0SLQgZO0/A1QBfz/ANKO5N
ePNtxnM7ZFJ0/0FZMkiRHvy2LzM8b4fauirz03VtaY0FVG9eZdaC3f4DH7PcaIriYdu7AKxQKSOz
sgBTVCemQ77S5R/clcr+h8GAORg59cTVmmSG3hMuCwms7Jcq3FzxmTqOYkUivvMVMCMj7So4r2Wg
DozSpAYLUvkAgX+OlghRlAqlnUm7hsZnxYHX+bE2tETqJkUF5Q2B5dYIXi1g/cLgvvrqOKsb1e3t
c5yvY/djAVd/1c61J8QKySYYBvF3kG34x5Zw6PokP9Y8tWFBIJEjeeRPUnbKUH7rsZ5fURAzNHnw
AJcDLQWQ2ebMv6Es3l5Siv+gtb80UfUDWdoEMSQ92bXfyKHmqbM+xJnF0tZKi0aVrBbzXKPXhonE
PmkNxEwthYel6zjKFeiMiC4ZveAshNf1JCQ5//qyOT19dFwNoSYofJJQODuEM1CsWU8EUredvcwt
iiJvRFt9AF6W6PB1+Uw4RlMKoPUat1xkAEsAP9DjNHv1GFc9DfJ3yjTUChA523heCu+B4uGCLW7L
HLH85khIeujr0qFEy9T0Bj9t3c4iEuWHMtGHQJ///90RlR+z9iNhEpEYBlNsCuEyeAxrkFrbcs8q
EFzdXtTc3rgDJ/6mcYsxkpKKot/QRw9sUZagsGdIBrxWppeQl5zvT/52J/d9Wkur/GzaldFPIjOy
eWvHy0dsEjckx9gUrXz1CML7YO+oSvTuZPaADF7m6Vg6wVcKargatWuDFiXkEsXKaW51q0FSYs8F
1NcmkToSoHCBlPjl/1+epHyM41htMw38O7JsIbdAG7iCDoiblVUL6sK4uwNpVYr9n/4DAhdyacMr
k4NwA3Xzlpf5yuVYVXFwSLR3zIdijua+gCDT5VwPd2NP8iJJ7BaQPaBSIbWoEXFnGX1vhXqEspnK
9ZI4hsnASYheYbrKzfnZTDrg7lOntJv58xJn3d60atjRMi1pYlaDblI/AEk3/SNx1eHtR8mhgag1
cT/UsT+840kgYLjA8OvEad6P8aunFzwtOMPBkg1KBSVzg/1e2BRuXuWaHRB1O3PneZshmLKAZu9K
fRY7fhDUn5DI4EHK4u02361X5m0234T03sx83FtX5mrsPbeV/faQwjGBWtSI4U183XUv7W/0680X
6zp+Gih4N/55A82IMSKiPYSEjODRXwqIsrRl5PfTqbplY34MuJgmNJKA6mO0Z7ORz/IHM4a9G+nC
dy0ssdlq7mXK+kPYpvLEmsY4NHrQaZG5W2KzqdZkoCEBtPF8qUlj90+cVkfl1vutVcgaGfY/6EFj
pQ0meZ+0IFbXuUAC7pjHsnrwsjm2h6wH6d9KRlaZ/HNLKDmKR8IIcRG0bqbiEI00D3tJKcCZutus
36Nw15Rp85J5LGLpjkQlNIhi62mPeDcRU43Hp92bVepssi2tOIjn+DtElCHEflde9eMLwjmMtioX
8xRa6J3YTdSS5s7WgJIVR7j46/4sN0sCbX82MiiHPvWXdJncE2SgHTeYMAp3WHyfkey5cGEk9jtf
zSbHSrZl9HsvLD5x1ouZDAF2amDmw+cnFWwDOZoaJQIrRaLRQGAF0TfBJuW7F/gzs/vdRWikc7ki
7qj6cPBC8uGVQxHwIbs2eaox6MazkJDs84YxAKCM658LgzxQzK+lNTj8APhjvc9CzhP4FWPHSLr/
Sa/QkmZ09ohinU/9SaQOgV623cYkxL/2z+wXWIrdjQDjNNJRyZIeJvZbChL0SchqKrnZA+DrjlOF
mx+NHjfWEhvAwl2g21RCp6xVkrj6W39fyA+MQmpFWinCpBCcRKU/i2kqbWaOnXGCZK4S9ga97GUq
59Wo4I/jz9kwocqLRo67Hati3EjBfB4pTWE4vGtthHTtKkdiJiLJKFEIjMGCoPzpc6Uh+0PYVCbK
qCcgHhx4QSo13zWK3Q5W1vPjfNHj8oIaTo8+3yoVj5N6Jot+qZy0p2IIqYvWuLcIcTAz7ECukrKp
LHSSJbfRAbyf4Ia6lZ9jp+U4aiH19rAVPiU0KzMryKfhw6RcvAU5GYdaefHnBgKZDUww/Vim1xgl
45ZMX8RdtPVR2wQq+d0XISaDquPdnt3CH+fAhCcxtQc1LmObwk1HjZZJ2SaB8K9H1fd+GiY3TIV2
9ZnAYafVaUyOJleL6kd9gs6EZIgHIGvhKcmO15QEYVlPNys04rXGwDI2VrUr4gZfDpelMnTrciCT
p8GwMtBe8SDfJUP+C2IX8LOzDf81TBvFBi1AazchCKlNpYsLoMiQ2hfBiY2kbb8chfdkiVVUf0eC
jWN3l6kwhQ38Olz7abKBTw4Z7rlc/RvFQAkSiHxJ+WYiyj1tpjny5WNIdi6OGlahsvUKopkWBWSY
qMSOKg9tX595x5uLic/TMa/3SR2r1p8zP7yKdQxEh4GPQq2CQgLiVCcMwclw7aydjov7+9za3IPA
5SRhYzKeNWdBhyJRCHWIk/Oh8QFJyAiNnkz2Jxj/sSjQA0IL5WKBb6bZXmpmlEJMc+jwoUj6DcEP
LO3PZ3LBjUWxCQQRIM0UMYwjnT0MgWMlpjJnX6UPR3aROIFdHTPx3bvMaB8BCa0+Hrfi04E4urB8
mi+uvqpKEX4gcg7y5fBgi9CTkFAuTuwtfz6DXzVed8QXqAGPSfyT+TrszYscQK8QiP89+0ZHEQp8
BX7itb7aOKmy0EK98f5iLB9gsqYcZuWsFoEEciLk3e2U3wY45gNaCZAVAwz8SLe1+YJZlVM1HzfA
T/sZ/ZfNvcjVm+BPYgPj63Ds7WdKRHk0iepuwcsjNldVK/vxIvc9H23X+zrm7f4pZaiOh7TaG8E6
5//yC4e5RkVRLR/Alz8k/1Vv+CYx2VsPalCwI5hrueQP/mnncLAdfSXCbTajSd8sv9l4FtdWhmzV
toQavO+LmRz4r2aHMMY4eIaThm3IuLb6AFW5UTCrAg0biqfSC99UqCk29LYVUrzMaLTIykFT1iHI
xFQm8Gb8DtwMoE7OMs45Syh5IbsWqGQf/RQPMEVGp/jETLasyaNyIW2DJV4YIWSpGdYML8QaLKwZ
3V+hr9wYiQmrMpDV/OoHtwOskph01I+4VHnHW+FmYNU8jM2DJddJOE3TuGZN+e6wymxK723UdUnh
VjchpFFbmB4OooZljbcHJJ7iZz2wck7s2ELuFdhDPoAacyawMhkbOKprQObmQz/EAE6vFqxJD4bH
QnRSwjL9PpaPyTee+53Aqrh1I+3yALAGnLfJ59IfrCIO73dDFpv+O6kmvHgdXKqHq5HjockYomXg
Q50vXPNAvl7Xiv4GXLe+9J4dGMKzgycVhiJw14r7RHD8X06kg/luBJvVyGc1gVAcX9mRguWlwHK8
m/lCBYJ+IlG0TsyPlSrCdMlmZsSc5XhMJb/A4TpYiUqDOfmrJ4rp/oIaUXlgSth2MagKxAjxiwNC
hP3a7kXWEK8mvzaNSrjPkFI5jaXWrwfvPuaCr+kqNiKAMaa9uHbVYu5PZYKXc18FV0c/86a7vD2E
JUMuE1tHAIZWWOk4Chn2zxbrYFdVKTo43CwQlut0bVbFPJAD5VlCTA4DVLn7Fzt6a9vSQbFrTN9m
0q68+3L8owWFWx7YJtI4uPPN7F7p1TRVXKP0+r/y7noSQfrkmLImBa1DWDALRzOZkaP+ygNLz1X9
kU7lfv3TST+r2xCcIsGH7FmuiRFWKa5djBq8Q4xWjydg4KepejmJxucK3TMVs/Pz1prFG7G8cVbj
O39FycfAnXw0lDnywpvIUlaEeR4lLXbgjDw1nx3R1CRX532d3EBf8t6T+PSsNiTzRq5ER0RjDQZw
4hr5UM1hNF2hqeXZO7NKftfjOOafp8VgQUVCyJk2VNFN/5P6+dkHNnIzObIDDMd/9K9yiXPIGt8j
ntE3hMkDfLH+njAIx4GeZ5TBaPD1CEDWyA3CcogZxZ8znh7HLh6Q1I0eFDGSwB8KcMr3WJTh2/Bl
DXuiab52F3tcwM72uXzhqmvebhufEQswUB33UCBIyQlPKosuHynuCiWapLOlB8M/Lxmsxjxw0hoA
Kd9Vd/apA8t+hZ/wg+zc/XrG7VoHUzCzoTOZHVD7VzKko1tEgyth+OLAuvAk0/1qMCrwnAf9YmR1
UI5/A6P2hew/HmJOE6QNBJTYfkISaJIquKPOcj9+fVMnF7S2IosIPNhfuJx+QoH4R4fsjz8e0iNa
jcjZ1E4jZXvRhH9cLTuUTRZxlugZYJUj6QJTxwGCGDL76PXMqIdPiqCYunIz1XRcasii7efB8Its
GsO7cOujG9kXzT5KRHZJVBH26egxHxGX71VfEyiWEl1vSCnT+864hY6W8f0t6Gf/7QGBUN8RU3L2
4CJTjc1toFhL4paVQpOtwY8KH9qRBDZ5PVDA7oD6F4sfLoZIwmb3C82fdhWedwhZrrb1Fe3canvf
IltIQEPsuCIy8sqtudfTmUjXlOCCKJc+qMd5/lg7qSCpkIeyBhEfTGoBiLZGwhc7UdA1GfIswOW8
18dfRYq2qlVKyw9AbJraKFZBQ1ObK33yaPj+eK2ENpgdrN4T3/WX9BHdPljFQG+ZlZ8HiqCUQh92
+wwjFkLERnbyNE9S4Wr8p33BXZABTEFyT1xy1cpfDnhSQYlvHSMmZoXouQvicdWh/+a4iJavxas4
sVl2zP+fc1R5dO5/gxOxiY0PirP3vrWu+s0baSLZ+XjIu2l5eCz8hO+0rvnz17Ol2juALBfOMo/m
9lpGBBtMVVbZY5BeATaCn14gxsU23KRppeToLp2es90MR+vudc4SK8ybJlKne0BdhV5VnZNhvzgz
EcNXOgWDaPE8TmoPSYYTK4wgS/XBE7qy83x9zYN8eTa+2kDTVl0ba5NPjWtyeAT6idjR1/lY/sZe
gZnp7T1nPc6/HsBdUc96C4oLvkp8MkWA4MUvrLQEXhOnfktvYHZwFkLT0H/iN2ug5arqCoc4HbIr
OvaSwGuPIazVYNzWrC3YZMmbcGxCg9dxf7jQJWISTp1Q4anGOsmYtgS79HRmDl5qcYkYy4CAlD3B
CASdKT/XipijbfJ2f9qKMtFkO9hNk+6jArLnJL512IxiBLMOHG5Ikwgtau1jo5d7VxPjl5B/THlY
hp6Fzjx6MaOTxujp30uRzGAAb+4lWhwfgf4TUsCsGnUAr+upvPoDzF9tm7vfVLyGb6JNj8/jYi+H
GmYriurM+Ag4jc4R34hZjfbI01muqX6EhHz4GjycCq3KAUPBbicGWbowWV51ipjgltvMpAy9cA43
CDfHYiLxS8W1I0ZfC5QjaVgyMpaxaBJDRTh3lVip12F1W1A6CbDQtiZ5TIZayOIgMKjGr3cJ3KCX
WYafnKtJAJuDQiFHraggLinEWqFkHmndT58/Ae6pjf4sF0TiJMmINu05TeIe/GsAXPjNBE5iEpAb
58uI3Rx5YnponvULIalPMdDhnoPCXZzq1GCliYIj8jQZYv+0NQxDPZDpRBP88zr4uQb1Blp0FIKE
tEeRu6dMaxrfWgfw+pX6yrmJ4XnEqzAhVYs9wmDJd4D/5tyJDb8SaDvC7/tHrdCjzbqQ1tMgWkDZ
+ABuNE/s5SmcItTKAVju7GVx7098AJTXimiO1tljIX0PJErrZEC+URuniUH+8nQMOxhpaaYJsqYN
Z7eTO5m2o5fu7Nh1lYqOvl9qR4QcUtHsMKXJNjpuy2/1xPv5rRkV7OKD8snS5PxeME4C7jF0nyBW
E0D8vdOsCk3T2QC8GYMUbGHfOVBNV/POLcGAtidPneQynCJq+DeT0NAukNwBU5dgiZ1oDKsZ6Lwi
2l2sR09Wnv6PxysbXESnHv9iwTjve/fB9vyoiCogY+3TIje5bmRfh+IeGKksmdNIESaoTKdegHwW
6SEMwt+5n/h3SlmYNz9IE2CXtU7qm0+7xB/nnst0VTUwA97i1MxusFFkY1FoB5OURZs/c5D9DK1Q
xhuQVB5YmsiePnWWVnaxaSslHPDV1AnhyCcFRnnMtmf/GUuSSpD5FqqTmVpw8eTgV/jwj3b3b9WL
7UCaiyo5MI2z4mnv/8mrOwzCdPsXSSttquC2BdIYlQiUPuTdGC7YwwJvUUC4d2csltqdWbUXOkLN
op70ifER0vMVAeDgyS+tpgh5qfAu6rLQApXKs9ZVuE07sD06M03h7V0ZPPcH7U4+Stql3xR3fAun
0yUtEXFkerMPk0EqSb7aNYALJBENqaDhNtXM4yvHureA9+1BpupxUPOQrzCyS3FsjJFfpmX/Rzmu
/6rK711g/TcBYKiv0E7uN/rW1PtcyaMZPWWpwh7VlOSO9LaucZ2+KOuGN/MLHxlYA37LmkcLSbhY
0I1mTAFG6sc9E+yKEEQvUWeUOJfoVg9sx8zjHblIsqFnv7a6wPQYwrQycOa6bH7ufiYDhIcoNH8O
kmyx1/CJkF7+xK2lOfhEcsIA8ZI6eXqMyEGBj+6ZoRe/7eDQS1+rxwtY8moXSrf3lReuIT+ypQ1g
WMxOJzGAep+SvU3SiXrmBP1WyHzIgT5x2wEnbP1CJnRkbidtEvledLSTUU5jneEEcO6XaPACYEma
Gd2ijy0beHwl6cfWdTW1w1dn3HRTldrEi/XvTZgEVNDG8nDDLYKhp151phB00XojNm3BIPRqIpH5
4hhPU6f298SYCpsVOaURSwrOUXE+QK+Gsnl1y+J2Z25OGuul0I3vBJ3baKtm3lKmvZUuJuRbYvcH
drvbyq+/K0grukgepZ8iJDZ5YgwsBW3tJuecXrWg4SQSEmzuux7NYIwmVQNwOZYhhzZS1yIhkymt
staJi3kKvTNc9PSQcDa1Bfk5ZdsZDQN0i0pX/yZAeucmSsOY38XoK2F4nU/u/8/Y+vsK01rNj/0F
l0YyLme2NMbCs8IyxqnlmzlA6IVPHSEpQzHQ4XR8EMEB8xnyPR7DZQ2LKLkO2nNRIWtlYY7c2R1k
Zi0qAbqXX7yfi39NvGvRJLJxU9t6ISl9lzsLSV5cXupQsxDvfdOkaVy6A+Sl5eF8Lm6ZU9i98KJn
fUQy54QKq4iGPYK1taqt5mirz88p1XwykVnQXm5ZNLruz9G+GRbCYstF+w4uL9FNO6fi0jDWt25M
sl3dNFBL7BGKsru66Yva9XOGsdEI00KE5E+dgy6N/Lx9+lS+0dLXANvre3DAS6Y8jsrg8vtjFFK3
mREBqoWvCmnLLUsGxTvmdq05nzp6aUlZyeENtxT88aMy8ibpYP0n4MxA0PH+ar0aszPHm4cntYdw
rjWmSDZkTznTk618zBWPNuZbchHdVecFXzYOMXu9/QS5lVgPdqEeqUAQMXeB7rLqHviXzpxEigck
I+ZytH++QbbeTVJ6YLCJqqAfpVggciYWTJbkaTZRc/UCTXl8GLTLyfRRerVTQ9DHUBzPpfSSQoVa
8vGcS6xz9DOi1tZJV3Fz6il5+uuD9g1ZUJ+fs8FErQq5W9mtrs76oU9suLimPssq65FDppX0NHwT
0wU+1a8d5/aaMTn6EFe1HKQrRQCkE6N5ep4NrYPwa9O0IA2XKvqT9j7LGRZQgkMgRf5oHITaMB2c
lQJ1t8FMF7HsZuKyXszwPUofhv6adpLZNyQakbDVZ6mNF1k/AUK90dr9VkEWkUTKQArfrMn59FbV
oRuPgxaO8iTN/deHFnuH60+9jGbBtifKyO1AAhle6TffQHiAre+Lv6Q53CX4li5YKIevpzV9IgNE
gqJ3tXjET6/T1xMSWKhcXwXHa/hLRN12NQ0xUdvzRlia/LMrKM1WoPtjtdHdeT2sKjjpaPRwhjkU
VJm+YIy5AQpUuDgJn0IDDL4iJY4kczhV9SaXnXj6vq+URY2u/N9dZBjLxdTS7okfvSmvxD9o81GC
t/AlnhOgzcbxUjEiDsmD+gzjCN2dJVO0sOuWonqwHd6dl6m7FANJGTqCGP3Wt0HX4qBfk8oXyWIQ
3IYdwyvgn4WgFoRB0ldG/DoiDjwNpJ+0q99ibKK4eG3owh+YJ3nXI2eoiW+hfETVRRQotbGSlEe3
poyC7FBtzhHKGwXjZHhbvrNHfrCfLEQjkF6k3NQ7TVBUSNguzUHGWBIxqnSZsu/qHDUJJLCiBVk5
Q3FhzJVp9bPyq5fDMzWwR1zuo3FMHNykAM7A2WZojBsqw9W7MUWsidAR3K+9pHt4hNCXTIhzeYl6
HlrOtU/jdV19SAjnI4royQOWtsxuagOxPAHQ7+CNl0TELpEYcz65Cv6loRZP/Kf2E0hPu4LF5LcQ
BGIohlJCvMNJ/dQxG92oRGXTPp8eSmMPoZ3hxEOvbkuwErhQiKjb1xhNOZVzJc3V6GQMrVOufIhG
NhfMukbLDBjrD0hJW/HkVw17KMB1xJJDDngfSAYaFmnc7n4IwNDmxzVWYc4/hz8zuG3JuoaDvb7w
JG06l9Mas9XMl7LGsoK6VEY0JgKI72rsiZjP/ZnfGzdQYjU8duObEYR3qZP3+0jItIPMc1AugP37
i5Po44O00nt3AqlVP1f+FweUfnON5wWfuuZF44/IPD+zAYJvNVdPqGN+r92veKJyCg+LT8ZwyTC0
kTSJRVky4OgHkLUnkNibaDR/17SHaEG/PDazLLfbXbG7Aabr/R6KEkrT3dDz0idrK8tgrjfxqxy9
aMh5+LjYDTXEY2jV5NpsZL5bJWGSKX+6aoUK+y8hwd1TVEUVmm3JoAZxQ8fGSg9yE5iy1eUTV/ti
WM1tSmufkcfu3SaV9HypyBa+b2lVCd5MyDTXPFMC6swBEm4UmpPPfWKfrhLpSRGxFwG0qbbU7h2M
j0QksP27XvvX3dtMjsJNkCxEgFPyGjiGGC5khbZtfSaVsT3LLIMQsCMFZHqe2ZRvH+WBJLlVmoRp
vTMp7EK5FJgGUklT0GSkTkMnIWEpcELIfuQV00IdX4sDo/oeWcCoHwO4PzTgeaFt1JYmZ8Y9LBZU
TsA+D7KSNPXAhkHVj9KYYE4cRNZxSxHRC67ZkwJie9FmmGxk+wmIbCqhvhFz3F2jRzdhmP3Ku7BA
oy+KU1dNNBPM4ES2jStKrktddx98BZvAT1DJQdpwUE0+bDdprjwXzBBV4qbIkDSXdosPwRqnXT0y
FMSAj84kzEDT6C0ufkNFiogj67c/JTy7yAYAL0TaGyg2G5/O3Es8NtzteDoJeLYMmUF1LPQ1pqF1
WVQx61RqdTUQQrgShRnDji43hlRhYZ+64WL/i0QRPEWT47uqc7B7Z/t90YenidBZ+gi22Fj1F8Dp
3mF5qGS4F00cRd4xyLgsGPUqG72gGRsdretH7kQYCanRBHwecMal8qGSpT4dJnhny7NcvjDzoNsY
j88s3FXJuJ/RcpmItg+aCHiC9gBQP/HZQ5erifuC/gJn7NPd03Q4CHukIQ9UCNDBoiQFwTSuqn9r
zuOetjMiSRHYj0uwLxJrVvWVupS4iwx4IyvT1BziE+jYTTXZzUTuIhfpFNjSVQiUH40DT/5+XD1f
1V7nCanWUQkTaMCPqS8jMaHVNHPqSI4YyPIvLgBVr5712dzWKRiNhIPFpTuFlhDM4STwdWY5rGFw
I8qWYisucGjgDUDt5TVumeXXtuKIVHOD05e0u1EkBXGzq2TYzf+snF8NMDn1aTKpq0CzQSRCwddd
HuB9d0N3SRBxJ6Gj6HkZlTorce5aym8Mgu0PDljFL/2l0/up1POGsQaWOCd0J7kQ3j5NbkLNIdcz
5bzaWKVPpi4w0sTZcXVN5WMoXNYZ3zbEhgOCZF7bVacQIZZsQpUYfRwePOWDpWehBTNl0e9C0SbG
D2BjfHl4UNrnCpVoe/AnS6JngOOLbr81pf+iEj24IbC7TYCf8M4/XBBMfoP382dW73q0dU/CjXdB
Lg8AyWjp+p04OCTpwjLobg5Asw9+kh3OLjPB/fJk+TUIwHce5sV3zUNy6TuWCU2ammU7DUNj0mAM
hXzFnDba+BW1Bg6Ks4me/k3d2evFADlTCc6s/9T+yEmPvZHWAyUI/s7oa9G/e75CpWRMlWjNjIjC
pbMk9t+p9+rsT06CkDC9fPF5LIoWsCaolpP4T15wCnHl6UGFx296tKDf/RrtMYExHjfHwNAneZmK
44Dp0/egm5EaKzbDc//0CSytN2uVo/4HQWW6H+E4xIMGcBDfgZD+9+JWphh2Uw7KmK80qBYosnBQ
nqvig6K3jh4aHUZs/yICTDe9HM4gM3Gq/To8ShPkPHX4Ir3+gq7ssOsuS8lS8AGl2tOlUToMwuq0
WQ3pnfi6hhcB1wQQkBuYB6rzeK6GLM3mgmS3UYXdawskB4w90ca2rMDLtd/wu1lAIHYh5sbNWixo
qwjHtPho9RonVdL6+YIURC6WsieXVPPo/gG3xG7nFarjm146EEu3dU2J454D5BB3zU2n5xhG9XhR
D91MIuHRUazdp7TNQjWJZ49KbcYuTcfK2QvU6KzoNxFE+50Oc3Nqpd5tHOZj1HxgQtJtthTwPoDo
DzIyUeBZbN3AsFR/ceWdNb0GdHVCbbSkCbY+IXit7U+j4J0f+IXz6IiJoINQEpVwaSRKjQsx3Yi4
Vq17JCQv/Ho4xv4HHMOdEiY0Q+1AxSzTUixdKIJn8IOTf35bOzuDgbF9xxcOEqssfKdoNbCRlCMu
xmM7KB597shwycKx+TUKrsbqnlgWxFoKdCJo8AQmrpQSI1+aEO5Pb7NJc1Zu/9yH8HevlAxeuBYd
yyL34oDZw6VngP2ilOthXXw8HEwakrtF5sQ2f0K5S44XkqHYf49XkOA/OKfb5/XBjF9pkeQSSZw1
P8xWO2Kc7B/WjTGVSIScMy4pQmd/J4pn1fGoa7Rx/C317NwhIfvoMt/S9V5+X5KGVOqDTHl9WiYJ
XXwKszAxNBCwmUZ3qWx7c9MCUBm8rRFC5iIF4sH51QREpghAhZUMxIP3UXYLrWGyU5E9EBCITFVE
fGUfmlo9OZ+6XTNOesoJj3WuMoTxBXnmpXYTlPw+Irg3npxuHvHsM0QKmGQVyf6jfnl1x/dW1Tid
D1wAbFpLCcACuEZ5vs++72JID1Z6HtxNHvSJ53LfgB3FsQ4XZGjoxr7rfnN/ucQnOmklWDuN9zKF
+wvDm64QSsBckk39JesHhpzfqxHNofKImeP+tg0Og0KMV9gwlZxXfUJg7fm0fFI7Junr94Ysgpjc
lpMgi1aC/19FPvcOLamo1JxbUZ1pQUXO/uCzdtfYhkyBDjIM8BQW57Mw8weMAdPyCTbhApEC1UjS
5Bykbkcz2R+QfGOcpvRahfJNyd5LkCOEkpldnrjpiTQ6R71nTz4h0cDkG/Jhi1Bxmsv9rWBUiSA0
6KgyLrTUaeNFxbvvWSWItK02pBHcDRnUiPHw2gGWMDwSexi8vNu3siASBfrCdA/xtmieen2k6mBj
w36Nq75ZJLUFCGhcDYWCyYkJ5At5wc7410DG6SD5xiVYLOuYa/Tnb1X6W+inBcRxtk/ONhUyfpCY
k7a+bY0aU0K0NYz6X/GgZYvmHzwxPYOxDtCwI/dB/iuMQOJm+a06JrNDI1ww+OKDLgTtSPgJwDfi
TilM0L2d2dQcV4Nxy1JJu2T03FQwPnX8nifq32ZhR4SoAnOWnJe/eMe9apV+r6G4SElsMplNVxaR
T7kI10YIZQSLUJ6MFiI9mjI3yBuGfDbi436av/6WxQMq3vDQU+o1yB644jwgeTG8rltAlpxHchzp
/8fGu/XImZHPiPx+iU4DHCqGSWrVrcL1UJKOxgHgKDHX1M6Bosj8DSeICtbCUKIcBlYWYJfdMeED
NaBgkwjSvldHYi5yKwr5VVkOqPASZTgxDUhmblXGMP4cSi5gI5f+9DQ9xhKorwjXYN7f7GQJxY54
YcMjlq+FGhp49G2+WaKuzoDcNVHH0hyr7CjFmVIY5uWBxitygezjBW2Oi8fdLgShWvOeRr1k90kE
TlelZwzSDjjhs0DVytfKe6nu0ctv3TC9R03KteZZN/aUQNjCQmiWaRFrc34CnEQ+VQirqdV/uTkN
IeXhuO0IXjfrg7/xilJuRA0bG6M+GNFZmMpdgy76MSSlc64+l2YfLQEdM0ZTjrBcWZ1UOKSXyk4P
2MDKEpluqwvn+xE93JUVciAlqPx3sAxkC9WqISN9yP/RtpxIJ6DAac7OGkwQX1kOCLkbiOjJ85SP
wO309aaSp7Ivt3ZL0gsC5F3JgsEcM/5Y41aujF4GNqbz8cMy+MsZbd2aHnfGfsMmmDj7Fm5wRpMF
yuIJjPQrpezvwoLE1OHXQJ2xecVVbpkmdKEa5nEjGrvHN5fHGoThsX1Q9x1qudXOolvgdrUY91UY
qxNpU4biXUYYeV94Q/SOvXBvElPb9qMo2H5wij2g5Sba5Z4hFkCSYA01UUGwmRHzn36bL/5kwT+0
RkDa4ZAKrq2QARO5j2OWS0pU/vmVC0RbvBXrbn/18J/CqrL5pqmAR4yfgMhDSXr/3LTPDStFW7rw
m7GCC/gfm+qX/CqMkJ3c0Ro6XOcy7YpF3H0+uUUphmL0HNHXPzQFZjVODCZMhEWa7Iu+N2udbLk4
YeqMZA5ZIUbnCzBbflkUnPLxOvwtxBxr7XmxKA26eAPI8otZBDA/2b7Inj7ayY6pIlsDtuSFf0pl
fqXeU23Fbr18cmOLkIW2523ucfPFyPVIRyU5kWQ2AN6B/7/4SFD9i8a9xnCVF/X0cAwzt+HOrxAJ
TUtpiD+HRvvmmBNjk9cKO3w4cuQiBRGf8A3Hs2/EARNM1oDNOjnEXeUp88OA0/NclC5c51CZapaN
JjcJ6rdCaMBaupqdrHjyv9P8z4S6H53Kgb1F7isvKbIAN3b0+YBRm51MFRGPHB7r5290Xhn0mGYp
FxQDl0M49qSmPF6etNmlz5tj4bOjb4EeOm5hdrBU8iW6XeLMkziSSWg+lONiGyCVdDBckjPYY7Uc
K9KP5e0oL1VWUbMKA2ypMrymn+j/xx4mtknU4vtzfLnotMt0iGBLxew+zpYh4DuZMC0xH9DFr1Qv
fZm3mreTGmqtYEwTo/pSw3sXBDbhUpIwKo2ARjKayKqqc3EoSYaDx2OgVM/5fmhwxKd0UnuHCpEe
Y2605vjX2Ufs/Ryu5AAqlWIIJ86Dt4RkDhtCc8mZsIu9Lw4d6WKPaTwTFJdrOhEvT99eXR16d3Lv
ZBGGajdA3OLTctE8UsdlEfl7ZLK5SRxXOQYvlbIa17Z6jeT0V513DK6Gj+B0griDgCfA3RasoBVV
3GBZzpESNovdq3239PgZsP0Qs2FM+oPskJwDvkAy1ZE/7HSpn+CPa2tm6Dz5u6mLVA5MyNrP9MHM
sP7m9cyA5/x5/Cd3eFkCg97mVF2Af7HJbvt5NmVQr0b98BNkjLOpfdDaUlYUounKdQDLoaV0BLsR
mYo6p1+snMcRAKrk8RXBvP43Kb9ZFFo9QijBMV0n7PfUX7f0LywGGxnDf1yQuIUyFdH7le/1jyKx
ZZYPcdah4a3s4RAfU8xunuqcuJqnOiVi8Kc47gKhKA/AlKpXre6vXJsuOk1WC7P/JoyWirSQ+Sjg
0x+Bvd6kBOmqfCLJC/h1EI01RF/Sv1jCunNrAjKqnMut2a2WibKuVaoU1Co5XhDpqXGNVMma1zgT
iaGXEJ7/8d6K+1LNYO8ETCS0z9CwJVT/hXWz7C3iJEra873d81CbknAAfKa869f+P76uDrf36f5o
Hx+DTxPXttxQbEHcpLamlltVLL41zOb8XKY9qF2O0qfpCDWkqZDeVny4CXzAJBpqimIgoHB27VT3
X9kyNbVlTwqVcgDUWuxVtt5WGYV0R81bK2iXgr7RHnVhMzZFAlygDNgXnuCJruYx83cSvMEzKkHw
8tGteb8ljXBBVUZtBDxhLsBpJR8I4z3+DPuvPFpBX0AjD7udEE8ulHzJpJmFX9czUB7UmA+laWue
zVNihKCA2Nnu9Ly8eSZROXxKU0VgjNdxYAQJqKDgBkIh3zPNbO++ypmBzeWlJPEPwwtaevDIq8wN
gUUdcfPVoxAUVHHGSUNScOyKwjkPnbEdq2QzUASuORD8icoOTqGBIqzbZCcLYTN+SfkvqYb8ru+l
qQrZJYwnj973WD3wnzgqZBycLpFfciIdjVlcf49CyLrs7WsXyercsIXDTprnYmk0vYsVk9JqGdt+
oYbv96tht3KIbRVfUbWBFGFjlUIx/8xyHXu4VDd/jCJhcTgBPjAM8vTdMU1l/jeiXQZkAZHTeW1M
oOx093r0HvllIGcXRqODJoEAqagpLozX1EGL9y176IVmLd6iZe8uEA+EFscnXMPcpx3wy6jKRkto
jFqQpdJHMY5iKG58/w63heX9LnfEJeT0ysBcwu0Ylc4CLECfihr/7FJ1jQAijr+gZcX/H+46/IQ7
65xyTOHx0/KU8SNZIOjTVZq/q6p27qzUED2T20n8ABRP5D0toTzxstd8jGzYeVlTxtjJyXOSWEqp
9mKzQWin5TUB/wVlCF4qZQZKBL21DeshJJ0FBxissjU2v3nwSfcwtAz7khznqxHgh14ork3SggHn
nPH2x0I5LrjPoEXtfnlmFhGUOGtLRlkFUd+n7AFNboSuSbfEegxl42xnDMDBz+1lGES/XR7XmgDi
QuMUxtr9aYCerXOkj7o3XEVlvNtuIGKK3yWKroMta5rETwDWIbMqiUqZM3KdIE5o4pZ5HQmmiBPr
LF3TKPNB9rmDUfzQInCtPyQq/nSXCQkpjsddiTqzGmijeGBqsQNhSmMJMP03TWPIScgkYiKIp/wM
+xQo1GTf5eQj6VnrRPvJ2hThOcYk7pPPEC79oR8u1LAKNlCICP7MGDM3DFANTT/VNh5kkKcP8XGM
Z8OrgVhzNwpC32FHIY/zZwoL1wfxffkrMt5YrFuRQB3U6fZTuIl5olv8W1AVeFceTkZ06U2mi2ZC
sZTtTPFOhKkYRuaD3LU+xaLReq2BfUdhwuqqsa1qZcQwZnfHNULbYiEkkJ13rkKQ1Mreblow6Gjl
B2BODL2a7Xoy/b8dvG3zqkqkqLGMb9BTvjZMwsxQP/JGpghxaFO7eHXrODPOil73hA7TjWK8ya0D
XAvDqEaE4FCpzsIiigUHgmt8a23FZEfd4SUarGDaf4ezhTmGWrhvr4Y44BngvTUOWvbfY0aXDqxf
z8GJ5m9EcgXHSJe3MUCwuxY9GPxoHy82OX0b/sREANODLc19B/1eQSztxjka1K1OxZ1xZE4sY3m2
N/DBXR7LE88VTTRSRJbhb2d/oDMtFmZ2cple1wh7zVXesqw/b5wgBqaHqJEkFWg5S1DXKCFMPg2I
M8zUQC0Pltsfd6wy15+RaQCrsXFUdElThO9RK9YhUy3zX2JsBAdxl0SwEojIGhn5YUcAPc3B4Gol
TEXLb4MHBUNL53R1bVkR1YEc3g1+V/cg9efeUtDde/X9d9j9I5k8WTYwbF7DSmeB/XF0SqgqSk5E
tGirNk+g3OIgbaR2CpCI++luoky3oAHVs1Yfm5YCtXGzp78HTxQWido2DEbxHOxKnvKzFrDPlxj4
wqHw6eKbd1S+jr60qsogTPZgmlQfQy82qctFbV524Bap38KgQH98Ip4EzG/o9Ea+ZOqcJivU6VnV
QhZ+SlMvjMiS9yczWZ9uTeLKZK4u09jAb/LxaPHpeXE6xANalMteMWNntoq+d2IxqhHpKJb25eDZ
lOVxyKFXcczcHhH69yTDOgqiOCKO640o43uEOSK0cRaI7uQE4c2D08GWFGsKz1yz1+c1bKgRax83
KruTCqz6XO17prCise1Ag3s3KJYj3KZJFv+iZjkNpADDt1ue0aj3jQomg8NN+MyyGZ93IT5xj25f
EN5VE5FbmMBZ3Ri1PJx+66O3XdTjUqIciEMck/ozdfcphAQTavLyLH8UH3cBq3G1XlzW+cdZ6gT/
LMzfnVStO/80a36+VxzhvwjMPRJqRdTsOIWXniJ9Ex0siFfWJLvM3cuijKeMApGHM6t364M3MAuy
YiwxC/3Boh3NeHwywczubzpaSlKvfd9N9BclpwWluzjbF9kRk2jDFm6PE19bPq3OwnGIgcg8VA1h
euCRIuN1vZSCj28e9DWbDtZQYnZc2GVYBTWFPDmLgCO9QZWf0/I4I1Yt5H/M9nC9exnbwRdBpu31
QS5g41ZRX54nlJuX582/84nUY1YVSLRwF3FxVcZSR4IZhJ9ntmKudykskSSbv7M3wx23BLNxHsII
9ZSinn0lje8lJee6XYFf+9av6/NoVlGwGlvORVlFw3cil2Dl6cvM63Z4QHfK8sxS4Q07ZOce3mq0
cHlC3NE1yhdySxWDz6vxebBDK7+Lkn1XFY+pmYbJmqkRYSBWodTpXTzzZ7j0CWYl+jhbljCVqS+P
Za//SDBZLNVK3GJ1YCxzUa6TYiLOJI58p45xVhsKxteLec+QEbB80Bdijk7DBWKSW+EwRhU3RQFO
oUY0J8n6dKzR3tLs1rvXb52Sels5I19nvvn25Dv3Ed/vQVuUs64wmnaTqKD7nXpzNsXl+qP+hXpT
IPG45S73aU96loriHRn0SqrTfoUvDDm6Nglm/GxSSvYwo3s5X6TqFuoRoJpEp8zLOC7OcefqxxxU
4czGINZD8CckecxKxA6IrF4ie7qpdwuq+qmCy+DXhRNapKrQlqWC2OhLMAPndTYRK6220+u54R3q
QJvQEWIJ397Cxq7BCmU2h7UkxKLWYmibORVQwZBlrimGov+C7Xi11GWej5kMAMgbcSAwO6j4B0SL
lBa19gFos18eY6ay5ksXo+lYONRz9qJgBkPZMB4/GevE+3xyELxBa7Zxnv+wCvTvz3TrHfHDkEFf
CJibI9rQzAEmCHVRqiuEDqvoU7UhUfJF4tdjFmIJYga104PNjwWJ3ivmy0Lx70v1YmFU7GD494t8
MELgjmoAHTl5qoN8DoyQliEIbivKKd29jgrXwl7zDXjDwrJ5jQXw1S1JADiG/KEgz0myTcEKt4Tc
0r/qNwfjpLFgKNmPOVEX47dQlhiqoU/BdWqmJPwp7DZIqnCAPxPOj0it5wHZ7QtJebEG3EShBkvD
+HJddzSSs02i+teZvu5b78n5eWdu6Nu+hFqQKnrmFnFGkme1CiyHDjgvRiU+Ao83bhglgWFRFHCw
aXJAqI22IRtfIBJHSjgYsigkrXJcYOwyBtXXj9xL5kCs+C3UcUyOeniwcYOLEYtQ3MHRfHEPKmQ7
gHicNMGJzk1qnujlpgzPv1jLd+lypx1+DO/RydE1qU2U4cONiJGBbViPEdkk/J8nyXg5E/Pu+JWq
9nFWDgghPPzVW0d5NUDt3NVvyEGR7p8AEzApWty02yPdXQ/MYMTWqvmudhwLHuACDxtrZprpW8UX
ODqmsB5WCIKoWwM3Qy/50H/dTISXW6HZE3XtkWKzyHT5yiBlOxKbDozBkwY2CuPMmJPya4+vTQh6
RJke6Exk7s/z5X6J+K5L7MLJX1IFVBwcwHas8719QC5CEomD0J33vrcnzfb/N/mjplquWDBNAAM0
aWrkqndWIW/jJ9WtBgmNCBoy2ixBuwQxHpA/jER05/JAfP9Nki0qdKovaVdkQiKOmYAqbIUodDSm
4q0r/ZPmQ5m0mWJTaX+ozz93lrpF1mczjrrvyMElSwGtukEfCEe1u1M7wC9WN/de3z54gOciW6PI
jf5UPhI7C7wu3yd6+qtDzyFoaqgfg/8sPaZQRWGr9hDfcz6qDz7t9pwiQ2enrQ7C4YEs4LjnKBzo
HsNd2IfRX2wbqlMh36aHIb8S22OfH5sPdSYhS+Bz7xKfGorc+5ehfYMnLFSjV1hVKVvG33VYvM3C
kLHf8ye7MBR5m+80Ul/cKzDy4QciODoyzE9GrAm8dli3AH1twzH1gpJHSYFRN8SrQbP2Xhde7UZE
jlqd04gM+5T97GDKLZSvnNIacXVTJGpvrNwLweiB2M+JIJI/Mop7Q4eIx+SFyyVs67GUFgWIE4g9
9xDHN5jN24yBC1zXs87nwcgcESWrd17GF1rxi7SyaP3ZtLj8aB4ODhoHzHi2ZNiwpH3F8Gbj6w62
kLn5T+VnXLaoG7yM64drArERUd7S6qkJQY9gYAELbE4Wg9yLQSwRy09NNAodXX4WS6Ymzxon0MoE
0A7b1PUgW6VE7IlI3e5z9DiGK7309yKAS9w6RRoqz/6DpRw5SWOGT2D1k8yMObLdo48MdJ1acsES
ZD5eaYySUi4PTWv85J+bDo0bg/PYrtE/S3f4s35Z568MtP5cdWN5Kfj3V/Uc/r+yMFk0qmbwhgnL
4gVXQVDNrHYXSjbP0jNgG/bAB5wLriuG1X9wjCCxyAYoOo+/b7jAtXjNZ3jT4tQ26OQr8hsV0LRC
an2MIRe8x8RjfJC0RRNBdPLbvWLHQI2KgdIwV9G5qUZudGz6XjPIZTjqsK/esXUHxtKeY2CzHwew
sGN8P9DL/WphyAJArNZ826B+ZyRwtlHS6et3N1otzS3wEHkw6dJBf3jfbf+kWLs/u5wRbUBzy8VT
mZuWLv6wzfY3apHs25rlCwgH4KQeYY7s4brQfP8UnG1rJDkeY5jwL5B7VY3GbxejbQqb94z+C+v9
NVihCG902j+PStV4sn2BcZ6zHgzIhd8StAu6OAiy+bxDIW3G/md2vWYuDHdGO/Gckv+xC7U+/0PK
gCV9mihF78Ny64IVZ70RujRgU5rK6FxHhxNJpm1VN+Ay2zlS5NLd8UU+KiqNLL7XMAukYyqMplv4
jq1UMfZPLrBeYkT4glRQEuLNqsIBtURQHtzeh3TqxKN2Qn4NhsLGHVTuSyx1mYLE+yFyMd9VxO2l
SRpg849yt/dqtYvHaWlVjLYZmVY2HLRxoLeOwXUsLiy2+cZd0OF+gyVHMEju74Qr959f+VceHkWD
cmep5JIjN07GogLUw0Bk0PAsc3P2QVWhlfVvqZTh4palgXAon3WTKVvkMIa2i/M58l/MyWq2a3io
DXf96QpOlWqbVKxhituguE33NvWNlAflt5cKdDP7VUyM2vbSqoiVod+rRjzH0mHiXyPkY7FwW2ZE
gWdBh04hjO6rJ5HiArLfFg5J0Ucc8fgE2Xon0HBBTfBbaiFex7+4+gmdTbaZNRtlcUQTcI/QURN1
N2083JAKdXudQ5cqoa3Q8cg4lQyJZI49kFlC6IMz8CbVKgKyKjIhCpzCyHRJ6+3sXEOUxIi0I7z6
nPFuCfjM6qVG2gLBtao6u81w4VeDCMuz4Naswnau9mk+nrH7Qnvm7t9ejwxc84oSRznbZB5gTC+r
7wZOivoFnxwIETHVuoq2CBDsZWHnfoI6TtyDGPK+yTYNgSrIRNYTj+cfHLENe5Lw5OO5ocjUoWwC
cbutu/ALAv+60VADYIcc1Jdy0YLTL96aTKcz7y35ZyNtNvUmZ1TI0uY/ZCCJtujmfbctfM9z2Qj+
MkqPN4aR9e8Ix8AmPiBzvQGBo1Qq3rz/6jg17m5po8073pvAhLZPLPywFjc7t0YXZqXoW8ypgA6v
CJ1XQofufjeZZObz8x1qcezM0tgSFrZn1rd3snMBS/T9Pa7ZF+oEsmOn/jUb6VQ4kz40WXK1OcxB
ame2R1wt27W0HtUIhi85HLTDQHGxjaEkb/D1NbY8CU4FlqXE2shH5VA6Nt75z1Ku/3hqZYYyRjXb
oVByzWR30HCw0QIYaUcbScveKNj51XVhe/WmzXJippean1HsdPu8ANKrOTXj7DMNTtN8A0HL2yCq
XGtW4EyrFJJ0Ep+2NVNAgtysas/E6kD6TofJmqUm/J0bhg17+vo/2YlHrGH+zrvsvCle8+jBFu+e
bE9gPRbb4xZ3ZLZFoJpMQDuUzGsz3mY01CEksdXhfzhkQbVRJpuWSwXCndvPFwUZZF2ME5pW/fBV
DyWxy5P0v68bbdWjy+Tc2xTaRsb5AWGntoE40OVjSpxQfyM8jfcVczAt/GG14w0RwSoQhgRidG3y
uniygAdvj2YGZ9lB3d58KxeVeplmcaz9pyexIIAt4Dvm0DklwItFEXRrITR++eEzj/s4ub7OVLj5
0QwJQL8jYRjeVwLj0nnr6t1+1yFUa89rFhsoTUjUQP6ekahEt3xQPFr27PFrzvUtXHlNLRQ+zoj/
7YMQD7m0J5md5SqYzDI/ImS6MYcmbUydwkYiCRNP0K2qKbLI/vaVdXx5RAfj1xPEx/PqGxYqgTbS
UboTuIYUJRpet6ZT+quYzPsbAvq9x2aP4FPxTNORf+9bcg6ebmA+1sNyhFyNtjbdQbb4tBimh/to
4zPvuRez6CCr0ES9CYOEnaDBRpIxg1FlYAMifCIjL8ngKoLneFBxAKtzNKejrdllnQ8tjexlf+Vx
r9dav6tfLRKk/UFADBI/DhLdP/RTa1TLyZmK7Ocv7Mi7hF5AwigfiXit9egbh8nskta4ObszpXVn
fMmVMWuIFhlbMAd/NVRYI/xSZWx0kjt7sGI+HEZ0Tw6z9YCakzIHfMjVjd86UB78pND9sk08TyJz
dfDpVXgQRKLFzbe8lPmppjFDhevKtFLxfsM0coFzHRsQDP2Dt6eWNlsqPfgX/1Q4u5lJ1a69DmSq
ejSGAOeNVDUyXknJfyzGa4Bg62S2rn2yNhxZJSFbaOy5NGCgtWvHABvXfZELuyB4V7oL+5OIt5g4
ASx3B8kjkha182GJ/+uVipScCLYLaGFdtP8SfiSZjOG1cHKb1IHcd4u5bbnYUKmUSjLOoDKTd5kc
oAaOjBNWMGkaE8XmgGHx2DLSNL/dh3DshNjOMvMEsLIGPKGSWi5KhlDHIC4yU8j/Rojy959NKRbt
vdmQb+2eLdiKuhKKRKdqtvAwiKAL1c1M0zxXHnuKVSsCSr3PdSiPAVUTSXfqdwWc5eDEOhWwxoq7
8N7cTgE4Lq5I7SksiZNx+EtCvwQzQtZ71m0/wSoIxHQgx7QMuGfLvPudvsa2/IQ+OhZHUeoPbAWz
eD01JWTZEqDWjsdjUjutXvAncOCTg28ZNB575m8A9WXrZ9lK1f1AhMjqo7o/aCeBB1Z4DgzI7WCC
APtztR9YMEJkde9JUCMmMtreW8xxSQ795Q5yPgxxxSGHo/RPm8ObEe7vNlwTmE2tW3EH7CWoMLhB
CqiLWzwD1TnyEVWBcrVuTU3+irlUewY9GJ9Ej8CQKGCWCEx5PWL2b8/tEyBcZkeG9lG8Xoaj2E9w
+nZwsSyYfcUZfhjBUjThSCo9DjPFv4IhkJ3XEXczhURkqhAE8XpUsExqQ6RG9zLGLUqDzNXC3Q85
bFTd0AXU9B00ey3AxtJhBYVI12vwhJrKl8uirjlITkKZpRhsyevVj06SLtD3hXaD2mXlN5eZZJx0
aDKldzz1HZIl5BjDwpCLHPOcTtC0lqWtwyTxOakrUOFxMh91zJkF7EC3Rr7E1sIJNGwOaIQlKr/C
tsdJkbBRLHL7Ik7n6tdV+U+WT+iQaaP543sHiQS6A82Qr56J/DHAFTvS3f+cMfLRxIlNfjtrRSLE
IXTufADXjAWD2oyDNLScpicXqWUIK3U8o8loAq9Ot7OfzQDGUxILuUFt/Z74D16kxZvyVCScnlc9
q2/8SuYpVJ6W8xM1WM8G2rhpx8DyaVbSroOoB0pzS0rf6IYLYg0tQjrO/cGo06kaArrzUmqpWNTY
7MZxWzyHaohyR3EnZ8QmHTHxc7NU3Se/lemRIGaNdB92yvo7Ny/X31Ly8SPHoVJv8FrOK1iR0nCO
irNpxTBUMJCARI0L2CR1b19yee5y7oRDzPZcZqJg+6vUYXYKWN7e0lAu9vu2nWL98otZHtvc0hFJ
O4zm6oh+lfDZqlUF22d0amKi2JH3ibww9OipKO5dMWXypR+u69qdQhx3wzrFLqox/n693GE2LcPw
0QcpJhsZ3SXB9vtYeLU/9EeMVmDouwEbOO67YtHO7VmVSJgYOAqFrURxHV19grxmXBuqI5Ixj0Aa
YVOsjsttv2PUkTHM/hw3gCnzi9+ObhmWxuidAllip3mRzbHpVfDVmwxtVKudAOdbgHahrHC8nbrs
hahWw6jfqLPznRlX4qAyxtnyPtYbggDzEETBTNjKDW8hx63289o3fXB+0YuwPVAhEB0SKLJ29vhm
jqV43H7vtJ2gQSW0sV5vBTPGQHQwaDrKiKIgZ9PntPC27K4V0G9zdbCzlN2pG5fV5ofA0BZnSEn5
CyngF72UAfjXjB5cSUnVTnvDYu7p09ENxtoMFxublfXY69PhAcmmO/5qcKHjEEpCt2gUt/mO+qeR
ab6P8QvlqMMUwACJl63EnSH6M+KScypoLE8xeXDpIGGFbewfdKR0QUivyP/EYdJYKSNZZeyVpuKz
bjZkWdSP1PyK9d515PVLQZMxe2QYsfgUFXadWEGr5j5Ep1urni8tt7rf4pvtnLZVbqC6GtL5nItK
o3ilAlfZyp0psL4feHz9NtGTV0f5GTvKCDVeXxAQ7FzN1x4tDNZn7ARpi+yVB6GC5mApXUBgF7xI
YinAnzGE+rJNrqDTibsgTQi032RMm7W3ItcRaeCRYQjJBKS0SmzaXTdFh2nz7aVKQNIkw2017GmL
F7OBI5JuV2Wo/HGqPvZrPfcp/q/mti6I8vi7M5sq7NnfmWt7ug9mPBANXAV5UlWqmEoVh81deQw4
NmlOgtJlX1MCWs0v/wBOkCiSoOCsGrXbLZn6V/mfsbAP6+sG5EppAhFltpzxlLV5Pz8DczuVSUde
ONNfxLu18+ay0qmTFMxwY2GFf/qD0w1xk/OH2jRmq+x8q/D4uYcXRa5p5zA+KqHLIyGZ0d5YVn8n
ivhJ47153cGvmMgdLSs9eS9l2sEbjASApX/o8TOtM+wn8yQHbV4FS/sP6luYslUOIS+W8IK+FRW7
LnUGhVVJAtrbji9Ir5mXELFelSmyaHwJSA5KbtkQwvv4y1uAdZJI3bSjJo0DUEaFFN6gLN6dO5iA
Koa9K8vN63t66oIHAk8hBocMgNBwYo1eUNB8/jU4iJSPRn7z0FtulhyPPy/9QfLCGZ0C2/Tl6nEm
9rYDIS1SpWTUwvEshrq45/zAcQTbwtP/2MWGi3BVEc7w9w3vtcWtFOitegz4ul74Pqg7SUmfv97B
InZ9ZRgSnhS4VtyzqvS5crVLom/IgeYgnn1t84MTpjKr6MF+VApvBj1HFGxBe/ORILUl/7L+8sSU
sgm0qnmeCRdjIROm6e1cupgG0Zd+iMDdpHrET6VJ4LF25k9mVYEo546XYkSZ99wwe+WhXKdxpSke
9LjEH1wjpo4L22eUMgvazf2a4KFNGhJq1nSRuJjARwmA3myJ/ZHIHZizl9PE/lu79sDamhv/MjL1
5O19k2Sssi7aIECuyTdqhVafgUOPmStse53PjTF5/DjmbnBqzrlyh7EcCS153FEVWJZt9ZZDDs6U
2N5pQb8nm2fjVvJDSY+18UwZMp911duGZ6d+xDD/nZd5aypLbrrNQNaSbGce0Kw0U2lovUs7qYDP
JbwEkuu0KBlwiupFkZNOOfJpu2pc2WWMbyoWH3uFwq3/NFOc93EoSqti4NXRFy2cBH8E8rufAbZx
u+2Q+0LSlDkCzPlICVRf0DRCAW+r8tejGS747cwtOc1S4hjyuBkY7StQETJ2BX3AgasHIITglOhC
p1GyzuwbfWFSaINAFV8GWkOP+KHKCcwVIJIYMFj4OtXARKs1XW4WsNxKgtGFa6+u8DXVelNN12kI
So88xIu1JEorzpoJazbWufFB0AEPpbwyhNR8ZDrhOmt2gApbyF97OkSj8HWrHgiLU+zQDpxFzzpc
rukfArUISSZUglUneCa6bnburk7ftf8a0KGc9kqbThLUJ9DjXwZXETFaoOL0c4S8SYrJoIlL2WQ0
I2ok2DQNxngYpfh6ZNPcu9toKIZ6+lrqPPohsWNEPempUKUDez4okXwupiR1clhtGgN8bIVUde/F
az9zIMUThZVdvQUBv0NzhzExbacpPlCV1e3MBDrZgx22zhMxTDKoZY7kYqJQLAWH2mt4+pmTeJmn
FMxAVBkon+Iyv+FZ+vKR+Qs24xRu8t1hSMJPLkHqwqqZ5tvWjl8CVrmRBAjStE5l5eXLk8tPq37T
GqWhAboCMZOYIC/N17shTnU5RpkVWpzwuiOzKZaBy5LoDlYmK6W2/6RL55D2yiDniWDubwM+vWIt
nVr04pWXqbXnVCbuKOznbqgEUqcquvZHak9pfkpYmjh3Xb6VmD5qBggnyPru1fkQ/uoeqp7eqkVB
jCHH8dwDewTOJIxmDdN9ml7dYaGHszBz3j55Tp0gY1I4z1WqRVjbzVBErPHG27DCU5NNQpFwCi2I
tC5nTFtWG7aRW+jgDb8Mz/XtJC1Eu/7JorbWCwM/N5o19BExEjKp8Byqu78hLi9VGqqH/BgL1FME
21jdR/BYJ9W4hoeWiic2z4qVacqWSGOpfxuxLBaBVMWZXVW2Wa9lSTzbVxhH+7N8w7DdcHAAgEd+
yHvK/UPXNlgvdxjkXgLsCAS5Q6Kevam2R5GA+1pIQYW/dRB+xUTd5uh3uaFQHfWGBHqwCDQt6a/d
vnn8HwB/AtUzmL5qzv9Nx2tRVwIrNXXHsWqoCiVJNaS2xpWAyqiA+K624cH3M4gMg0cGX7LWz8ld
688L0dAXlzmFIF2zScr+rjORrSwrdXiNFIQNFnppAKpP9iMHrUDA8y6m+gUaoXiNLPjOZ7ZBO0cG
Nf+g+rfjvKronu77DdMklhA61wNbYmnx8pt/roJtzugzLlyRcyykxfvKahxO9vbaQTb4rEdckHPR
fRSxaUCzOj10kfP9ynT1C4w+vM5LNjcQlwKo0JfhHsYHwJeXyhzCzjaVno08pdLF7uNp/7kYP0ms
XtWnSVSBtyl/uVkI6cqaMglq76OO9Oa+k7YYci9iIuLGjT3g3m0d6+yl1xGKvI4EjfuMmZcCdQLI
XMlSbBGThDd/DoM9iiPfB4UYLZHUdT7kGxBRFPhhPb0ZTI7P1MduL8nwkO57h3D0YhwpK+34vZes
+gxKbYVJMhJU8VS8wBk//4Qj0tH+b67/Hr3UL5+IscNVHSkffdhF70G/jRA7ypkgciTN+UUfCnVu
dY/bpIyLC6J+dTTya51AMa9pOgGK88HA7BWI75bw8tWkyEcop8JoqTnKgAwDbY0U6oCmui7aCrbZ
4/Hn8d8/wh878c4/f/Fj3dH1VCPCXng6KIhpzmppisKgGBWYfVAOFt7inXlptmbyL4zZJ7kTRtLY
+UBveRCttgx72jXL7zpF4bwzA0cIL11j3bUj56ufhnGjTUpNLFgjoDEy/GHdqYVYjPtGTKg6PaqK
1Trs1lqcDw15A1/q01rtI6dsFl1aWd8RB+x4io1q3NCmkEtE0vmv5oqgrNTiQiEpLrF9rQXvwnR7
YS01lPX/QrGUpMOEPx7TEdHdtNQskMiUp13Ja5fOjFh9wNge4oVuSxtqZ+UhjZq8nxVYSu3ZrhBY
k9BG92a8d2engrP8d+71hmyJbzF9P08gpiEnnkaXpkyZvJy3TQA5PYGI/psZ51+A/j1PB76mSBfA
3FrSfu6oq5xuYcHjulpklQWAvxjCLr1N4KtEYYIDNTaXRSyM3/kL07sZI1FgBqSqi4lp7f7gK6nd
1rpZORKeaGtFdeQmBPXjjK7zR6X+abUcKAbEFCtCqAo0b7waxO4nW22TPY7/yhdt9DJ9WN+hYEp9
x517Z2KDetbxBArO8yhR+8BrOep1Shu1zNEiA4gbUasZW5Ye3kGzBAoFR57ioIO2U/ym5S+N130m
ZeQR0zB1g9Wd0oSuzjQeeqSb0Nx5XC/2sKibiUJfQXREcfbRkSKDB471Rwh7ITDNnrTrTp4xE5kU
NWvnrOh62hTOD0hokOmhBM8OZFgVYbY0sx6yHAWldlkYkOTZ83SoRTflYdnNtsx47Ck9KGnyYgL1
EEl9tY4tK/n3FkjCYPEG84hN4g3aQMwKUBPAoyI47Z9iEkDKtBoU9AzttR84OSsZslHsT6ZGsY7x
mJzN9ouB+U53RE/jpk6Bp51LSbzCw/rr5/pfv3573Jp4GDa5p+R4lF0JWSwaTxmQoWwmNCtxgeXZ
zjEZ2SuBsiWOjfTWkMa59YD0cq7DDzSeWpAWQoEI6ZJttln7ao5B24VOZDTfgABKxLuwJOA//rjX
+sMx6YQVjiA/GHRJKLkH4KwfG+gsyh9uwuLh0J1HyPMp3wLNyFTWsSxbIhF+k07nDRYo1Wldeo2K
JeEJQb9NO5nJMEduAgCj/6SgGoJOk1ttf3cr7ns2FmVMxDWNFjxnKY0h5SVV+FHaK38V/algpTLd
eAw5Q/LF8dS8juYE77tli207jKPAZSNRtFAyd5r5wE9OT4hqINdijNXNLVnD5s0U93oyRo3MDQqd
bY/WR5SnqxaUpCM/VXaMyzGBIgwjT5kcDgl9EzQmEa+gr7+0zCXI2B7wDWn0oLYfAK8cbK94A5RJ
WIIRhkbPlTUhJ9HquXwYT4eHjaMWS007dGNYY/bt1ekg3KuT2ta70fcfhMae15lYbLzYfh+x50jz
FufBEbMm8THyKgh+KPqodCuiCDxRg+nfS/lKy3mgIlg3qRpiU50pQXHwguoaDdkevjz/Nn0ophum
2oS4kKySslaePi4Q+Wl4wHj2pXAiVaqwBuydA2dpk67eahttpJ6H8V0snBcLpDcJi5rqt77IVNcn
DBd7WE75Qntg72cTfY/A7VhLr12oA874cYIsYDknhl3ti3qLTNHcP4v96nu3PYT/fpMugZOeiAQF
X7bg08SVoOC/XrqqTd3aDcKzqaqFVvtY0RbWitJtSlliBYaOGHeCCPqC+IvxYUVtQFjhvJ8HZYwJ
WqEmrjzyEnAyxi41ikMAqUJ/8GXXs9RZHPK2ar97TDj1bObuv6VfP91YzXL4/9D75rAIG4IK2eCf
bYI+1LckiCGrL5OTx6CXO/Fq9aoY30zCXYjDpym4NYigEp5uG2Ees3dFyfYImMeVNwiLzY/kZQhT
Q0lXCS4Qag2NXvdbu3HjuqgY6EcECeLOPSRtdOHv8fV4ag7kp1uNuRPTJSqTW7k7vMRCJWiFeOiy
h31JSRUj2gqgl3kQCoFOrfT7J8h2u8gV87MUgKwn1zYwKxV4TqAeE69757DoGo9aDsmcFKlMQWwo
2eCcQQDOZ0XAJAlzPB1kdGX4xYfRmacjFqCth9OGQMKWEOJeqvN6F4A6Xl0o3PXH5mCx2o8SX4oI
bYyEXC3IwzFz/0Wf+gUbfp1hxZD4cMMTcsxkhZC05fOS0t0ztlP3EFuerKMDWH+dBq6cpXGRPFL5
KdUf2/rrmrvtnEbEi7Z7pgu5vYJKJR/bp7Otb2fEmtqOs3hEa7jRaM5Bp6brtvFAP1pGocLSrAfU
Cd53FEp9zgvNlmRfpHo7CmH1dWcrEQ9XJ4sS/z/UieGKPm7uEcZmhUs1KBHmVRz70MYgg0OH7nD/
wYkEyvbGkjeKxnSuSMovSGo2Kdhoukyc4j7SCoie2W/KftoMGAPYFstqTFANwbAlhp7kLu5iVgEd
4p4IjAhfIPPDyErQ8jeuaEuejnTfLIc13Ck8+w7bjTtHH2ZtVZEn79HO7VKDNH3tvgcBkAcp0eQL
pv73ANVAnA9xTTakTEgG8IUgNTZdEa8eOjIaNrpATAeKDBjo8cwwvX35HUkVmg6jzaU1vziGAsKS
2ngSKQYp5j2gkqDzSf0wbS2g7+Qp64LgyZj8YI+Qq3H4nLTBRxtOt7oHlEo6733+zotT8oc4LSIC
AlviLqAMtXKnPTafUuhMfyaskm3Wk7MJe6LOXBPgUtzBj5tSiXsFFD6iQfBxv6GQ0ecSJ/DKGz7P
xhYwAUohOVmeTloFrWDSzlGVB5NyY3TC5U1g297iI24DUXK7o7iNrkvlAp7xOJHT1jLTgADBdFC7
rireo4IGw6hVhisxU0uiBg7rK9Bz7eJ19ngjtAqF5ES+WFR+mSAVB3vwS/SLCacdCqs939jpAls+
kDpQtlcMnsGx85+QXJJnuCbdkAvKGHJ9t4K68XcY11DlRewgeY1Mto9tMmQOve4qZHK46pBPw3ZB
yiw4sDj/OBhlq+bsUy415RwEtWUMMs41V9vxsHEFdqumEFBlyYrXezc4rGaMjT4FKIFt1K6/DXe0
X7vxylv/1SkhpKI7WvOQhndaBEBRsBWT1BTNOsn9C5jFBEvtHNQ07VlVZ6Z9LDz7FcnaIsTMiV9F
tQ+J3KBzI+PTq4UepG5PGAEB18aO9e53vbhUF8HoSZAFeikXaWZgpzleXx0dLhZdNJYS1JTeOZiO
6dslEZqgdIkPWYybWu9WLT/B473Aof9ZpDMBoNWeUQAvj1OW59/lonzou9wIs5xzbeKXGwM1ITfO
sFNBTa8+CamaIExXewbS2KOphKK6H7xnUKNJ+biPqUO0q2654tR7Pa7lbUX4VjJ0PbU+kwRbDDu7
8n5/Iu8BbMbUIt3fFV7hXDb1wTyTJotYpHSrX4x4laOrDpWEblISKXSJi1wrgTCg7E0Gi76v7npn
SCSg7QErbrnev4735wnuf6xzVHrHumCQ9rHTbmUmMLeR4+GLLjerfnxVwDdq7WeA06mtw6Hohe2p
0HzuscJfEKqPUiVROy1HgW9Ab52dIWufgh9tv04fK6CeCgX1EBjgYNZs1/lNOwiFU9cZ++aJc1z9
av5D2KrYrFWa189moVTTPKMIaBMDicfuUJhX2CUV+WP5OABxgAhg1quEEDgTrq0H9eMIHwUN3jBM
1lbxRSMiGfQJGz668x2JxBbesbE0Vgzu59OegjikfMDT3Rl8Jk/RbJHBOwcwYev8cq2MEfeDuDkU
X6jLxenXtmF81GDXsqyhW1GSoJX1GKVTtz5iRZyRGQ0Up0RyphGi0LsQZPGRZls/4Z0HweQKcNp1
GEGxBGiIhklKHlhyYXcLD6/x0ny5GITDv86WB6G1w/SnqpK9Tz+kpTZENsJHmmsD/5vIDKks2vyc
ySmcY34JJCoR5585Bauo0XqpVmXpI95h5WWwUfwr5BkBFzqLYyhP9XFymTiaeShA7SM7GBntiYYH
wbEdjAdnAA3N9qKKxDwA+QZzh6rhCz6fo22OzkopC7HE3CymkOPvrtv36/ooKkamrdlFTbiKpvvs
71gxy4LOWwZOSY0O/6mfcBTwA+2sKPnz3oBE3zfqH61/eFnjLC9oWeqa+u7cEPEGzTZVHaQ8b+Qw
FzXgT11riMcRW2Rt9732CIfeZUzSXuamZ4rA/rElfEGpbKayoZmFiZVo6Wqm2lxVyIkAB7ihz+S9
sK8KcGb8Vce7mr8A81muCmKU0HoOV69ie2nAzG98zNG0oVN+FVkDmgvgAkPv7LoeO2wBTSwl368f
C7OshLcqPHizTe3lSCRfwiWivNezjWohpx1LopBpEPu4eFHdl4WKaKxBchtd7s6KDXvv9M0ZdTaz
vxqOljg0rW5b1md0RPW6qQkEjXw/3fNGkEk6DC2T/v7DK3nzCiDB/T4MuQQG4TYV9ezWOtbgBPsS
tdfiV6YZKEfhon5eXnGiu4ahEz1dQoiStMgOLfFVTRuic/XDG9nUFpWzLJsX+/L8bSToPfjsK++Q
msLtZPaMSmGE6gSd/aIaDxhdLCC3TJhIg6UALhu1AFZXKwFtCXXCWeOiEFkzQkY0qZzKp+SUMcEa
YuzLUrD8A0FJzExoAbnvukWa2huEWw4iM53+/vmlq4QrAC0YwEwGcsFQW1yhwvRCRvmhpHnet5jW
8lv13GN/rw4G5GW/5Cebjy3CCkgkeK3JPhrjDr9ZTnUPPiwAPtGOXJH4NCKC8TCGJfUP4tC+NiUE
9WRrh6bxqDvIG9CK38UFZaS9VeM8j1O/ZtHdbbjROUtxvP9nlxX411pTKMTOI/Xeql1gVu9djpnp
OBAATGyrhNUvsSvqYL8cN5g3k6scXpJW6GgYBcopKKOcsekG+nYZNst8l8Pi0nUQgX4XKGyQ3kWE
eWLCMEtoeA8YKlPtMbq3m7UEBPyg80H+EMPI1JjUXvSqL4GPmqRCkEHd2SDzz65CkVIl5wb810gR
Fc5Ra9TYQ1aVHa7rpUtLmiCFw7oatPf+7OU8P/Y1rrkEnFRxktJwAJKwOVMoerSsvSQqgbb4/izq
bq3P4bAJEEU1MiTB44ePlfVNttu3KY/E/6sYx7YM7fjJH4wyesCn4WPG1KJ5ZlSYD9uVjz+6F9u0
+F51kLLW1qQdShrg0PdVniA4LJ6+4QPEny/TpphNGSIDLRzYWOekDSdhguMVS9DNvj7tzVa5DV6m
XMEvsK/cWu2r+M2Fupblh4FNh4ecoN3VtrS4HxJuFiPQfJ4yAQNLUunJjH1dHYYsbPuJvEjzebWR
tAlg1ENgB/PkjofCW9c/v4i/sCmiP/SIa0PTAU1oLcvvhMcL8HX+vtq4b0cEeX/Gz078k3eVN6SX
WkW65jckdSZtJDOiv2HPHwrIRzhGn8Sw8IxNXCwCtM3aNPUTc0qMzZyHsovcsJoAstnZSTx+veMn
zEGMPH/CsAcKbslwlwu13xh0fmpA6N1aB/fuUCXGsYrRWp/E/+nDi3jMijlHYK/snlPbxlGdG5cf
ou4XDPXpeEkiM37LDSN7bH6atrczdnJzPGYCoSx1fjRl0jZ2cD4rIPDL8lhJSM0m5uOcB5d6qR7I
jdeUDpCb9+zZPne5bmSwxPRlcSzZq7feboc6hjq1z42+7ESmmGxtlBMp49B9fogaAxFuU8Vv0rP/
TbxahVPC8ssGEK3DDoKDrf8HdH1GWJRU+QE+SfZbEdOTJwSWoTvaPkSdpG2gd61ZRerP84vgWQXf
kdbf21Pxt4Bzhodj7j1l+oAeUNaqxRk2l6U66FDvqESs7+5jHwI6ZQ8KCv9XEA/e1e+GM7wdfPde
WiBplL72CvRXfcAwilRrJlRf5kdFR4lOlhmEjy664tfnveyIBO7bW693VGpWkkq6FsS1ZJTNBv54
JSnEuapJHePhJ8JvEAkG1QBMn2CMe3WDoR6lUUUsoCwBf2DGq8HacNSn8aleG6tG2Rgu0dl2OhQl
LyaghImqsK+uPp9IEJWWwggAYJvFy3YhrIokcf1G8suYOaUzUAUB21dVb5NfGh48k6rK/B53b6dV
CJIKnAV+MsXWAd7KO1eMkhAqqAbjLk5IsiButopwDdM1tY/DCFqQBOi2/TDC6xk9/+ZqAi5q+/So
p3R1gc8A5fBdiHeBzbeQnRQtRG+y0Aqg6P3bu+kbiBaOpXLQCS9HRIYV4vhRUSqF6zOBxBmJg1/3
SmaL+8lnWZeTM/UVinnV55GavZ/vaeQHrDVfWmVAuMePyYZ8EG8GPGBKEY7xyfax6OsdNMAu3FzM
ymxFY9u4atSoNs4wq7MvCKL0+Mcdffd7xKbzKIGIm9W26JlurgdVJay4h3xIq8SL+ie+2P7QAOa4
QoAQOCyrAbDdvtPuaU0qhiIyrKh8fabf2RUAxjHSliMyCMP6j5rK80V9242KsMfgfEZb0vh07OOz
3a+SPmCEYUxAiaw6xUmBcr4t/k7sQb82KhTTCaVzYh8prBh0t8oOWEi08DX6xHP+PrMbqVWac96/
GrYWDRzhTVaemlErkoQFfa+8qWyeQ3yTx1ZyontM9Gswsnr7z0pZNUACrOcsyeTsnva0Ogri/dXP
gd4nqsO5XkGTJu9cbm7eetjxMMIZ35VrwQ69ZjBR1fa39EMPuzMz+/0DAJYL+91OLlTqc01Fhc90
RezumUVUw8Cr4xo0bJyPPayEYjx6sPNsqY0SuEdgLXjYpJTaNmOPShyI1TW92sw4KZKgAhtYCBMv
9dLuzV4WkQ2dYkfOmeyYfWlYSVrV5JBjnVWdn4nk88gNY5h53qiEmBU6GxJQXUPF5e0NY+pSxabc
Fzj8JpWYcUHK53dQz03UJgDre8jIiimFH3sU1fVlai1UEQ6Q3rgI7rRN4BWeWnU9OOU+a20vPdrf
BV8ptZ1sUKfraEI/lXzKtM7e52qziSsCyZyRJ39H2f15rvXCwS89YvdWjHgQnGY/v7gV06RuVkUN
8hIhnK34ptv6UtB1to7fQZoy1YpRLMWeAgotlmv/wTFGq0mZi+Vtpq34C31eMpJS/OPpSBJr5als
i6s0xBg/fRNYz8MP0xayzO25RWQdBzAx0DQ4dmKL4a3eJMMSTMIjjoCRYQw9lexHeDq41rZWVqiT
3+WIloqDTqW7HoRGvu3Q0eY49K8xM5MiOJ1s5FcUUF9Gyr3yALJNazvM2/QaJ4K9hMD69+iyKF+0
gRB1WuHJJSp2KwcPO0QyYDYjG44FEPN4FjFOAAzcTUPg891H+x2n25DtU2CUmrTsQU8ne/EAQNSx
jYD7nuoya2Ap/7oOq2gyO61ZOei9DExjZcghD7Edw0G5pzkH1AKc8BBy7L0ScicvimRDvIKSwFN7
/UQPd7JvJj70oxmHcyRQMPP2o8LxMvFsst2GWY2z7iaKVqH3S3QJfkAIWJo86bjokKmc6US4QBu9
L7ftuw8Ol5pEKH6Qy5U3zRMvwV6oFNwDYs+O5BKOXcoQOA52Nq5R9k+sx821rKah5I2mKm7RkQk+
jUddXST0w2tClVeAvOdPAsgnVYy5iLzJq7nI86BQDVoeoOAsJGjqcUHP+HdsDQYPQpvKuvh+wjEZ
+2U1OMeLo/ij55vWjmzTWABCxDFHyEV3TDe31FqbIaFGkWuDuJ0CjHUXmisVymUBF8im4j1qpaTT
P62thOXZ3DsJFWLbc7CNo+CztdbH9G98/FnMO41raJmPkfl5gcTGtwDAIsthL6YY5g/jdWMTp1ZQ
3nAOq0nCiPEdQQnx0b8r37ZKslG5qeCn6yfJKFYt0e01zLayazJmMHmCs14UpxqAePz9MMz6gmLG
mEEMgj6Utde0JVZcIk5WeZmknOkljTr0cct1swc82qgs0gCg2d4L/fJHRKqWJiIAW0gHst1KNPtB
9UPMYCy+r3GCsA3J4nbV+iVHStSdyZ77N6owF1xgbBTCSEH3B/sa/s2z0ks6q2mZZ8kf2R0PkH2Q
g5VHonX4CRDCGPFQYpyBCQ/Kp+QRHLTYoRLeUwBGCfHhAQwaA4SLczWZrkCgjYSud5K+ANSC1SyE
G++LuMVO5NpYvAXN9R2i4+FUh6K4hFn8TkP2+JADA1zlpjdB5tY8cPbk6flZszAfGOhf4zZPz9tG
hl7+Wo56dG5FkVWHlIV3o41XZJvmI2rG5C3UmuWBqnUjybJiJQeNU0eT05OMjP8DCxwVcbextJN+
ZHDVKipcWH8NnT/x/GKeqlADn4jJLbugFMDVorcnD2HcXy+R+8zUIfr9AqxqnZmlBB4ffEndQgDG
4kQ9YXaT5QHPv5G4U157FGvCoeKfiv7zDljUulKqldoFtHfIm0wpHTZa8pxxxw7knNozEGCKpnip
6zCiq/Ynw16zz0nQHb5SW2fmCnwNN9+j+FklWhXo/PyrhkP9mYVYSphCWEw3AxhEf7A0GWDIDrQs
o86AbM+KgKL3NLr8XP7Hbtg7sob38VZF7Q8U/W7DvG5APyS3sx+s6qKtkiO1Cd6vNpHt9F3z4+2k
ND36bUEXFf8Ix3c+Dp4DgRkPOcfLZubofNsCsqLnOrjjVSK5WigkwR7T5MB+M+5JP8fcYa+7u91D
VBKxKyYGCYhRf9CaPRNFpgmmjwTLkzygBnh7U2ueUYFehICZ8Uggka50kG8fY6FVbrT6czlk2yTZ
ncNjtvJtzvsh8TcYZE9Rhi5jf7kkzX0FDiCXPLGudSll7NrO+JEJ0iO+c+CgwhIY9nZANJwGwVg9
qk+aoNXNWExDX34XraiwUmD6LZVEXU0RNtoDZFUkLydqE9WV9Fr3/1oDzg8K+w8eGl0eSoC2L6fw
5U6N0Wwm6m/+Milz/wrkNoh8MngfHaSGMCEDdWRCTs697jeNyav39YTT1ZnohFEQ/aqYU2AQVStE
LYVZ4Yl3bNrQZkdQYGtEX2retAwF11CwCjdVwubozkzOhmmRa6YCOU456cDfRuwzXaVMVHRw8ANu
JUTk3q/54HGiBetj+xwZzxQdhHZ6T3nvsalv4zFpwZtDTZACUnj56r1RSzt0Pd581JEuOO5PJ7UX
E12iV5bpb66jhd5m00b5tx0nfJDLGOVUPZcY9QjCeoKWIfNMaJg0mBkCfHX6fyI2bq7ZNVG8FHog
EBV8xTHIF/kM/babWEW7Z4T4AwCA8WY8bvy46y9ALyzR3EYAL3wvkGRTMCzZd/yxGxkEkTYKUzOG
fMA/q3XCBmDsfF3bhWNAS2YBg4qulMzCHZnvYqPEYe1NF++IGC9rCsESApyK7OuFRc012KM83ysX
2QWQhkaSDv38pC6SgGbouz/9rpgoqSk2yZUCjat2C/2ssFpwrR/gcVusesiqdRHepG3ZSWujWF5T
GfCuuJRtBzCYFHDBmFlA1GmtRfyc6ma0j6GlxwUtbFylafEpzZE/yLIqWeR3zIag5JZ84Jy6n+Uw
WZ423Vzv5R0K4zJl35q54UCIyJyw2+FpeSL/rUcwDQqFnZQIqHmfzZMw7CGfDrER+2K8CUv6yKvz
TDKWRigLlrGiEHC8UBr7TUqy7tQTN669uTrcCNoe9+2edL0grrTDiQpVv2nmZsk+znsVkuvOipYY
zvZzjaofVXGzP6BKsA+abFbHq9ZgQhj7sXJ8Gt1fy5195bHCmJUcMNhCjhhc+1RdbrdLXlso4Zo0
tEZPuC1ZlGXKnS2UGCIHG3NzQ/HaHwJX3nVsOTfz1wXO/P+WF3hf4Evl8D9TxxE9n3z3OeQLWnAN
miS3nAA4h74Zvg/Lbv9kvh8K5HNPeUo8WByvQP2OcoM9rEzl7Xu6IpEIWHRvh9lA99GH5Bbr0n5c
WaC4qYhE5ealGO1AHpHFgI7oVzdmPF+M+f6i9izVdbkqU8ilsJ63FHxgQ4iPA5mod+6ZbqBNsAYC
eyE60v5v5Ux27EH1JMge4lUZM2AGmxfkfzMYWuu5QBEtZ0pDWWO2bf1Me6wkC+GKGBzSwIm6c37Z
tlngF5g2xB4JmnEjlOn8e2ZgDNapKC2OHqLtZIeflrAIn0BKMnYsONkmlU6UuuqBBen0KVRjVKTv
2fOVdxplK095SjDbAycjIpJnd4sRPOreihCVL8Yp6KkQXjXZ9IlxqLHbNendQFp81FhvaFuPl2Xu
BfbbsZ7kDwCMnHTMQEJSpRQfx6a4OWnGlvZYe2DDkiilJf9SzkTbYQkHKooL2nq7zM7dXd3Eh4JU
qvko4QHVOE2fk0i2k2rzqI6uc7v7mhoBDbPcqKNeBmTM7o7t0fj+wqi3QgqRYLp/wQ1OCW/M6eBh
NkQuF4FXGS7jDeZAo9Koco5JXx+DOs8BRR+Z3Kui9xj0d370oGbJf6e1qD+PqWU95IuGxRua0v7A
IAJh8PITyOf9Y8Uxmbtmm2hEnnGpjeVDUSWHQ84R8+Pfn9gSqWeweqxeFE4aPTp10JN4jIfHDaoL
adRmgeK/QxgHZh9BlKc1lXNs6P0PwEwqRKqi05N7bsOTV45YBmm8CDGfFBikL0trvjoI0DNwl+KW
3bcPbNTjGjw4PML15Ejjc33xYIMUtn1jhhq2fNOS/+qVq1b08Kph4ESjdFQlcINENZKsRLzsrsCX
wunl8ghq4Lahrc/oQbGB9+7Pw+yaLB/AiDHSGE0hln8daLZZYimFB7ULCivYpyY2AhGPde1Bi1C/
5YdryAcvFfUqDoz0i9yJSInAGUcKPKBjUg2FNIQY6hBhwzMt67YPrirYDQS1vXiEPG9nAqNh9dc4
mHkWTOV8bdEyRVDRUdwCkkFemUiTPmYKJKZXn52nC1hBeLMBaunGMTap/8oGMXKTdOteLtcCURIb
KF6XhmA9wbjOTZ4APSve190g4Nq9w6Pgux229cR/WAFi49jdu9BiLhZ3yK26SBkfPkJMPcV3BHK1
Rwki7YnOe1E5zF28OXF86vVQ1MibDm5dUwpeS10QcEfr5x4NSafdHwjwawF9tcnU/1Ed0H6eYvfj
c1JfBLWCdE+dRZue5Z8ekiXM87CaCeTOAXV/uvAHc2XOCc0I7xKfh9kbeJCrhH2TVkRPjjnX5RDn
1ro7aU2ynfG883nWlRj61G1A3MVhdFylqQTfo2NFs9W/w1srYJyB4vYsBUrmZe38u7trfwsHGPUs
+1MQY/Ep2lWWGueVmna66iXTv9HX45RWAqvqaSc2Wrp9sSVODyqEZtxSnGzZUIp6bUpOjPq9Uwd+
XjBCerg81yoRbAZ/fj6lfSdL/xr6c7iN4y+pOZpnX4aO+Go+NY/yQCQeoTLOzF0QBj+k0UAeG6MQ
77HyhyLG9svmPJWSD/2CWsobnFNTmU5BZEH3gPqGEK+qOCA/egzVxxzs9Mo7MzB/3HB3sDLdywqD
8E+QXnlKqaD2xjGz6PMm7fFhLiGyri4e8A3o6rUgURelcSkMgKg9XEtjIttPi3ErRMUSHs4/SdLU
IlB1CyHtH3lUZygEoALfi1rkrr9eTlKbdtj3enVP23ONqS2wRtxW/sQUqlCPp3WyVA4kr61ts3fO
9mU1qlD3GehTkoBUdC5TpkrmHI87iCfqqaPrXCwtS34fYS2bmhm3CR9cqEpcsiMHE1+f4Pww9mR2
cLWZLU6m+i9GkC4GYz1rzffnW7f9/d8Wj7eQfPILq8L24qocnSNUcKJrB74N4Bq9HcJS+dQvduFx
6fbsIcwh2Jm3ZqMG8XB3Iut36hlAkrfIMznFWmHTFzXxT8RrVzZJRGo3g4c4XsyADRpUqcHVsVaL
FJCFcz/b5UhX105M6qnEA/DzcGuKjD5Hdx8hOWUT9Syhk4TVpFuq80ZFDfcy1YesJ0LyaUTOubuw
1lvQIJLpxaAZ2IHusSYqJApHplKikHFhOLIFrWCTIXQBygVeG+Cw+RdArdYJfTWiZAzABV368P3y
JytLi2Mu/9MIWOSUE5r7F1i+80Mt+8k7xe1T4BoWZyXP4sWQkIP8hyoPCmZxLbW4qzWUw6vaLUcP
W2aad08W+mKxyaLi6OH0/p0nWb1LFp2Z4q4t56jl14gd4tECYHHYr9rL6Tag6FPOoAFTXfcSUeAl
ABs53DAyKDCjvH8WgHKLELdNunwrDhVDtPX+zHj7EJCcuUhdnF7mnBDOdBobTObiTWSpJD9dz2WX
9VNN5PLY7YjEMu27wzfIm2/W1GoxomgB04cwdrvNMvi5/i93uRgwM8YZOQkaXruzj2DFvoe+wnQ4
GAL8YUNjYKyzp4/fJ3o7hy94TzT76rW9YSUciUTbTzR3PHP5837y8uD4/oULsSCqzzQhTtv+OO+e
8AkJ9yOHZxG/rwEflownoed3wCsX1B5FmVb/iwL69GIlW4OK4lSDBwNiNUfALDbrixmg5m4JvySY
fopaauc5pX50zNKPIF2KzsgJMEU2AlW8bV/wCfo78hwOnkFIm4WYRREt4u2Y3FFYkgKsgNIC5YIN
S5W7Oiy7c20aAosPT31XDRB8Cwz3aGHUNq6heCV5txdJ+VUq7AFhx3dv7zQ90Kqwn3m+QIaC6JfT
GahylvUj73es7DR+vI8/S/1V/wAcxj80XERdcYjVj3Ec3Lx4hJnGEcyybF/vHtPg4T2jG9z7kzET
h0l83N8BTpZr09fX0G5Ktjzrdsyqtxvon9nBiy0YdAPG3EHIsc5NXfAas/vfG6A0LWKdyTkEkXO6
DI+eLJNjDYd9sN2FWmOXMzjhm9cawU/b6cJB0+eyiecCA1JM1ouaGpMoPaeS0pGGk0AbOLFjNQSo
MnZjoWPTnAZKB8X46oLp2bq/iEFPS6t5meknHC5MROk2W5ebzpvXP8NdL0QLJb8KmAagB5GVkdzA
SGTIrdKM5GsXR5Wj52mhVM3c9xCVjgNXQxrW79tV8xh+C8Fq4fMDLAXq3j2mhnA01eCUD4+j6/eu
5TABtpBD+p8ldSzK+oKmFkvv3QslCUfzofC6mlkri6BX1YrT0pUz4Bg5Kxw/6RSK0NxZpE3ffsBj
LtBsJ5rCQUAYqV+qj4u3RRcfG9PWZuDSMU2GmcpG1GTghuknNU2rkc1qyV3NJuenjZIfVJdhYFi3
gHTpSN9FkwIzlZwMy9BYBTQSWXQWHBrK1RW5kgSV58PkfwMsxIJgrOUKKjkIvO7D1QCy1D47xleA
ejErxyrsljbEYwptvOAkGBQbA/tUnKb2QY/kYEk5Z50o5GH46zZSMGlkHb+pvFjsIasD2qzqz1t+
z9Zj5hWocqqmJzSxqRW42u/ytm87YsLM19sGhdvd6IxXI5WreflmTeg1PVdlSrkzz1ndUgAnSSxb
4rAImi7NHdkyLHI1M4OZ/iJwK579jkzzq879pLC3b4soUeXos+Q9JcDYRgymej4YP91cP8iAt5Ss
kfr+GChZBIvYAWMOc6r1GZL1Nv9zFVVKWBPTDcf//iE3L8ZKfPwT4iWi9EXOpBDU5s6YUADzJh21
xeZJY/0j1+uKjQFNRlzX9zH2wPcFL6cy8VaE4vj87w5PqItvdIIL17mejpjJeTx4pE8rVqr3r3vv
NIaU+0juzwk5a8nZO+FHNRw19elV0/mymmet8yRI9zsljam/iYBIMC7P/Te5pDycCjy2xMZ6pcXY
jttG6tRLo1GkTyc9ueAFgb+PwLPidDhG0xZb9oMS4JgPmQZFt0iO6Bx9154qi24JpsNymIcjANMr
Gx2OHEZG2/TozzJ633JDpLVHrS1dwDVlT6QhfW58x1Bt4CKp0x4tH5Wi8v54YNpneuuRSluihgFL
j0XoQpZgYJ8XOiAtn8sx4cYfDLl5gvN6liGrDAV8GwpNEWhbZmDv/LVHMHclhZDo/tUnsmFYzP6z
N8FRK6UH76BqqO2My4VDg9RUGSlMRpyOri1eMN6nl80MpMzv+mZPO0GKiKA4AqYI4z2rNJ7dP1BW
+x5acjIEwMUP2R0j/DfLhKaa5RyAQkMZ2GtqSzX/v9dTvEr55UjYN05SX95U2vmQISBSaXMbVZLs
tQyyv3P2GpEvSztDYXCwz0SXqtBrBQPjSEFXsvUnqECP9No0d2WNrr+S1nPG/yz8+OBh6AZF00KE
INAHSolDniK/LCEcg1eGArASkjr+dMnlCub9xwm3zL6BuXifxzi7YI4kiTjzCvNF3PeDiuMTZgGK
qWFVJ4dZJt8nhbeFzWzh71xs9cd8D0i1ZoPFC+tZ4PHNh4RAWjnwvDxeVRQl0rIULoWPxH2DD8UG
Ww5vvJSOZBU75IrnJ2Fz6Messs01ZnnG67uJyqW0c19DmwOGbyH640DRS0zA1D4xRftb5w5GqthW
bHhq/7H3eNiFmLqV3oqkmrF8HMvu9wrIaQnOotpOu4vM9mzssAIX+7pz0l0DWIlSxe3uZgD841uJ
jZ/X/ZBprflSqSnf9F3uAhtuda8wFEMzmgZoshkzYLv3o0n+4n4bJmBo/WTITXT3I3kYhdJN3vpo
iSKDxrOtT1X9E//aJbR+4kynwP+QbtU4kvjWVYFUBDDUqIDeEr1IMzoE3qtMcaPwQ0iw7LE4RPz8
7n6pGOfepe/dfPhshr52r36NyTm9yW9ofJfMnHBcMQS7fOFAZDtbrmG7w4ABj9LGiUnO1HgSCOtZ
RtwKasYs/9+6JFvp5eDUEPcKcvG6N2ZJONDslGFlGZWAd3ppTQ2mKenK3wdtszd81hp/EBwn+L/i
78zjc3eRaKOrIb03Mj8UbCyn7/0x/KFaw/vxKCz6X8ZVWcmNmwYmRREGJwdkAHVITqdY6HzgohGj
ZvaCOkoZqS61CFoAtJnDv2Ij8U8dW6joiisVDbTTCdB4BXyK8bBhA+qkjT6Z8uBN/HyXOVBpZTm1
pTVikz+iJfQmSiufb0EpXMdODjTEv/pR8sp1V5GwffwWDmcSu9lD/SqVXQPBJ6X4Yd1izllE9TfC
7ld5Jcm9sAjZ1h0RruUL7bzK8AI9Qq2JkVl/VgGZaunb6S0eLZyjrY/nFdgVJiwy0p5SfHoAD5Hp
dxSW3V3HczX5UtWukJRqerd7z6kbvCoOL2IHLYJp3NND/Ki78KSaWr6p41lfhkVEpP3is9fq5KqE
UKTknvhpFoNVitT4HghUv13DXQVgiYZMYkZH0uGQBrtxBnBXKm9qAIarKFRhWm7HzLZgfZq7H80l
/xDZypzIZ1kXtdjx5s8HeqdCR0tu3+9b4D41EkAv1JBZmYDI56sLCTOQRCF8w7C0b1p8ngU6UZ1a
nBj99j3DOOtPNwtGOxk0w9VTFYfl9+d3oD8QecoGUqqUfjZe08/Y3oVcAgD8PpWmmUdmovu83lt2
+iSmwHpqB6HkgRkKoT/PWd+FxwGuC9lkv7AMFM78bsB0NL0P8OK+AGUOn3aEZHvz0LCS84cy26sj
gFiKg690wBQY7URx4g9PvFZYYWuawiPIspH+cSmpXPbrw9F1ckmdb2Cw2HgJgTI+04heb5cJQy0K
6aBhnn/IhzjJ6ArkUTNEmXIChatyQ7bKdHA1LYAN9SoclBlUG2Vw17EWp3bjSTu2Ji0xQzHwPRt8
xWELt6I6YvOswJTj9tZGagZEdXNPWBxguAXsd0ysLVtjTgEt/bB5GvbT2S7iA5bEd+05l16K9uqy
OlL+AwOKgu0O4jScyXLzSSjfkD5q57ps4HtqdLqO+kHxnT4WOK48zFMCJUX+3JthCp4/vqvoXAJj
TmaEmP5WY2RVWdPqWrjRX8fwiNG/ZXDvjLKEOV9FwpnRUKTSLZ6/JkTuEK1iIB6lFsXOENBR79za
+urLiVu11Nzhvu1VYsfcHcnF68hOzOyB1vIaw40QJx2hrL5k3D2qY286nYPQa73C2F5pKjOAXIBk
ZUUqomd/rYN0D9nMPKkHc038n2cNEhUmIdc9gryIo0kFEMKTB1Mww4+48HSjhSUeRhIDCLiduEu6
JESGHQTfu2vIVMYEr/1ZP076Rc145eUpMUnNHFuEEtwFw6Or7Kdxp3Kdn16q0LukmJEWkTMJJVwV
w7ggpVmWw9lcbHcQk4sYbUoPl4iRqHbOFJX12uojclEcitYGcTm0oZcQXmO0MEUpXNKDdj3iIzse
QjO85eNb8ZqinY16nkxwd+8/pnMVWHvPL+kntDQF6LIfxC0V4JaBhbKf9cT45h5SQDKMPLSKi0MJ
tXMu5kz88RFfhqPAzk8DAd7i0BKvGbCYFlAkS7yNetAYnj7ExqQO+HkACCCnXpop7PDusK0Gh2J6
T29BBFOa/z1cDVGkWsCtkx0bA2ioHk4yOml8D3xFdO5ADCUQCJfTYNveRX9mnI7qN+Mmq7QjPxCa
vtRS4YRb9bzJ3MXSTP8WiTpitBGo5mXkqZxvdsnHMt+6ZMrOybZ7WgjhIZOBBvi8zteVHaNWmcql
zYBz1QwEWqqxJHZdU0Ce+2KRcSIXVmlhgd9xpc2cQqlsVP4sI8vkiUrWDva4kmLbiOixkv23fyVM
VzzQs4QMMV1mLxOyI5S90QLeipAkq7UEQDkyrSlpFmre8rkIMvoXx535pLDzzDw5rrDh5eVxOh2J
otdeF/rBjsF697+l2q1hamr07ptstBd+Q2hFMpmcEzC6gZkNGQcZi3hXIx2wr4OwGNhnUJ0G9QyP
L9emoNX7FlyQo0NYKr4YmPNY9ye3RVRhJx6S4CdS8Aqj/V3j7BAOI1OYvtPDPJL4qkdwlEJiAR2j
Iy+0uVOfpFwEYqLkzRcWjN/twgqp1lpNxqLtr9noj34G1iCROoe4n5rsVQ56X6eNWzGli1KrXmm/
VWsVAhKf6tdFvOsp3kxd3F78EsVCP4jH5G5IOO68jtVd/aVg92nwyKvQLmhJpK0swAR2es1u5rOX
9JCjL/UzITdL3gktM5pOTwyflmHN1AOMJLPRzBK6WZDfxu3AZQdvNZzQUhh9NIp7JYlFqhyRFhEE
U/lb1BfsTHaUHRW3zjExjDlA6BpUmkbHV2bwrWm7SD/Z9IrFKK0JgsA61zw8O2E5SvT1I927hCBv
vmIocAjL6keqleW4GtVgKseQbI2h9k8vNjskv1FcMpXCP+vJxpO4DHlwZCfmfqJD9XNhOx+0vhIL
qbeT8KXnFbAKctcdQXCWTgiLxIueVM0pGa8x7kMG/gHY1egTkXMhUANOGUNUWIsxeEgYjhXUUX5J
GHlj0nfae51xacfxISYN/k6H+zQtGjO84nx37AVpfeNStazL7TsDQP4s/qdZEuL2Iq6w2XQmt/1X
f6V4dHROd77zgwJxOwrvULOo2KqN8xVMe0wcwGS+agKt3cKljtJhoNxcLcwGOEKkFhGBdsvcPYiG
wPBW/1oVTOQC95zq5H9vbFrpoMNpPTS9xZOcGbHk2Xyxz2/6StKQGk0GDReSqyeyfVLfFG+CjD25
6MGzhWZmOeuv3IgZMUlj0zO98RDYEcdeU3iedCrOkewO3YWbWiOedgpW6ZW38CfSarn/0tWip6Er
5VvD5sV2b1Ki++IM451StSwe9+JBi9W9NkLWumN8OFb08BcSHEvlw99NrwJcEOJBykW08AIkQ5b5
6D/OycCrsDdlZeVdoQNk1+8tm3NSZ0n+O5KWe8KKc00aQLLZwrGmKli1XkVQC2Br63PGRjo6Q9He
FiOhkzGm0TQotAcFGmyRpl4nMr3EvVLKemESy7bDeJH76vXHRmKOTduDZd4Af0n46rJJipah0FKR
W5w1XI+TZQLUXK04dSjIGS5QK3QPAFcm5AGmHZkK/bSxbx7VJkkKsZk40lGd2DDSWj+8vDkLozS+
UqRgMHx4vNbtIyAb3BQN8avi4YkrmgxWei4bSRrV6iQ4zyWWQso9N+gnZChXJDClKH/oP0T8v9Dw
2O2Srr7p6HR7i1nKD8RMT9sRZYP/r3dth0L5CtnRuubRlNcXayR/1ly9ce53piHGBG5hbenMRCoE
h0NFsdO3IIBcY3K+xzOsv5Gf9rorBsmBIdrMApHjw6jadPfw/stG6kiZxiP5rrjgnXKK/iVi41kD
/APRFkaaRrrhQY3tqHfUp/ehqtdyMtLCebSyur9iqf3BudcOgOvzcQmAp4W24QCySMRgdqtXaiml
7YdwXvQz9udRNYDXwG9+5YILmRm39SgYv3aV2pyvLHcjNj1Ga6/eiQaW0vleB4otlQc/9C05qI1c
p1GKpnyG+rQ+cdEboE7YHHPVAxEX3yxOgYvsSmM8FR/I2ZFKOr3IGdjdTwpqueVW59M/WSloFOak
tWWNzye5rH8/tdOMIuLd7Fsgm9NmQ2q0AjlmC+Zo/6Bf/0bw9jPmlk8PcstwXCscKFWsF2ql25PZ
oWtDDi80JeVGRtX+VJppjfaCB4+vlx0YhqDLbjH6+UUDFZlUBJi9bvCS7BMSZcG3QQb0c4s23TqE
5oLZc+mPjAND7jfaTMevf2buDGPyp88fyCps6W5uFkbL+tBhF1e6SO8uXLKpOpk3zfLP7dlUpVxz
nMvOOpinhfn74ASc0pogYa0Xk+ZxkcW4AgZAjiGJ3AnwD/uvAeeaCXONJ3BF1CrLpzon1/roNv6b
vN2bfu1mrGbm0ibRb/pIGvLs5C7umOQsoEqwHxkCFlsH2kpDWzmk5xGXV2uhwseV9zSZGCueXNlI
AryZbcTht3WiAkr73H6BpZTKBReIs0FtN7qSOclCE5E3EVWFIAqrbiLRgNHSzZMVdIPXwIX8qaTo
+F0W7QMNIo8Lne6S/Kjdo0v/rT8iX9CcwXzYN20aaG6vTKDBaR5FBHiHTDl095zEDFANQdLpyUcf
mCcwD/09yoxAY8rL3RFLfg1Kski9LaCfxhrtQRfTluRobwloLJ7VLYrGwYOClO33k37hN4iml0YE
ohwBTd2uZ5SS0GrP325U2/qqOQboudQXaQawgmYZ4+mFQRBHNVJL8v3Kv46/A/8bl/DTN99qtH4h
ooDs6m7Te43S7AcyQIhNpvQvwOBHLVt4ujDfbwP5v1lHcsVhE+E8Wc8KXmfHoziqjjGY/fQLKY0S
1guWJrP7pQQehgIIqozkxPMEdFB2Lsvy5v46kakakCOsx6C/HEgwGAolfb1SOv7Vll7XPhxurP7U
zkIvSqMzgFjUId4MXqHQbNByBULgmzHGS6x5geUK1tKSGhYnUn1HZXwWjlZysOsjaZkHYyA+DTm6
Qo2VVBvJQLhGXRRI8RnunMWWiD61rAMzei2UrIhAut8DplbaxzuRAK2bB1T4zF+WMnqoZW089/oJ
5wvJnMSH3mKTkAecUwtHv2ZqLgbzcKDKIzvj6lKLgAcPhUpfdGrg8MtMgeR5M9xUcB5Lov3TUyJ8
wRUIZr9zBMSby+SrtwMtg2oqrr4gmM6lMHR1NAVGz5A/MApakgBCyeSyFdQX1Hev7iADzBlFMHk6
q6Fin+qD6Ythl2RvzWSB/aOT+DrAxNQ2jEJ1IRbuX18ukR1PGog+aGUWCMF2yAEOtONvCd2sqzdI
8RvoLjMNn1I/q21i7ROk7piD/NdyG8A2bmuciuEIe2iZCLjl65d9xRP2GhYBCmDMUZvPejwgxmJI
Hftzo50UhpYPQaRnPMjMzqhlCNYsFIIALVIta/kk2N3jUiORgwYnGkZFA76lkXMGyxfID0mvAMBo
VhCxNtwAMlZwHbcuCHrejOuBzmwLVytctgY4qHHE1IoRXlp2qC34p6bXWDD0BFSMS+TJKABYBE8c
5qstRCfcdh5anjCQkLMuTI6VAIFPdGxmgslSGANJX9hsTQmoj2XQvJnucb0THG7g84a9quPy1p2j
pbZu0POYXFTHfBNlB/Y8zOl9WqplM4MF84b8OX6jFhM1bxjENQ2/lhaMRXAODxLdxK2FUuMW03Jw
45WiB9/RcoTV35xKL72W6F/70+JIt8/ko3a7+RL6RXW1bAFrJ9hChZa0vMbvYn1gV5AnwC77RBI/
lHsQcMEKEW4F/ITGikSpg8J43VFNgmgPXKfI+XycJAcxSZIzgEeM8Tp0PWt+c6CrcfrK26rniHug
UMOaSkTr4fzb/gKR/RKe65tEOhfLnGdDwG45x4/97w/NX68E5CsiOpEGrYVHoGzbWj8Umzha9w0q
xgcXOEEDCptGhtd2DkKc3W8cciaxmwb9KMDCQCUHSfLAXGgdKpAgjI9rzTtEJQ8Dew5DFWJcKAyQ
qZ9dpuL9tIIwtbPlQMtxGrPzD2O2CMYbDXlCvqfm+epK+FlAQXFWwL8nfEOR/qRoUws1sv246Zll
VfvEH1eqfmcOVEsMA67dGZKHR9cWz9IPUmrYGoTrqyWMOmpUuNZ5hL9Pec1b79WTH/ljNPaurKBu
hif8rbBQtU9ovQytklTabJE4Oj7/sBbtIEHefcS3s9+LffY5zgUfpFITK4Cd7nqHW+pCgcp/KaK2
e+Ac4kPQpu+o1XNFJA00J41aHCiI/617zrwSMuQEGFwj9qd+hCLcGS4wRayHTnazz9h37ouvp/rM
ON09Y+ZbLsa0ZxCj0azsua2eF77H2QYfZUyoU2JAKVmanXyCpz+Q6hJyY7gr+DWTlGBvPH2maHrV
UoJSPVEVJkWu4Enlp7ISsMpozwohlQgUyMR7g0IH3Pb4Ycjfu9KZ8f0KrflfA4MWGaYRXAqy8lsx
EdO/VEbAD+4eNiKDxLGddKGVqd56JttIQIG81PDKR1cIqVpZelM59l0Xt+5FIby1/v/5rddM8Kz2
bU+FR6l84oCDRjEqLVbawEmtD6lr0nIOKRe/NS/UVD9nEHppAkFRxYIYCnirhVVTPnrIktsFzNhz
M/Ck+YGBfbFp9O17i05T0ug45m0TqKMrxYwamUVhT0nciFjTA4ceLof0kMvtf5uXOt+Pljc6mibE
yFxYW39/vw47A7o3pGtPufFYcZSNO09JPi5j+hpHoJMRFoLzbAyGyBqPCHkgBePpQEVGKPSTaOrT
SB4WC33440XZ5XCC37K1lTEPY1tl6CU9GCuYm79dXj5ofoNRvh23iMGJ7hkniTZIGY+6SDfbb7+L
lxImZIqBIMyYaKqlNtGpr+vlnSUv9bZ71T+fA1N9Mc407E0SrN7h8Ifh8Bq2Cbu5K3HDIpTlhLy3
ksmom5tN6BN69ilOfthKPcyVPIi9MdStYnBogwMOvr3SgZgVokmCpcTR6moBqdNhWS7raex6LXZM
D5de8pS+xijqyVknyuAZYADzn9MgZOfeJdCjfElxq1HtsIWMt2fg+C+ut9WyMLlbPuW5iF58w62C
AxtPqZBcCv+Ey/QgkQGgm63fo4RWVJ2xlhbewUHlwMsRnRcwL89QIqFQ/Ang3tFOvVYEuv5j4ZzH
aKbbksAkJRWSbjjcz7+KXTRPQYGdd5uhcWQi5y1X0nk1pgkWermwoOnqLgqxAALFKa+1h6XLC6op
BDuUJ+2kM/WtF7kLYtb8Ml6WENjIO4rapJYchcECZFuFEYKfGFmgrYZIgHJvS7qLUqRKp5PZjP5V
54NV7jH1fctRBHVb+CqmbAAa/6Pk4QL9biY3oIZ5ZskJXO6khWMsdnWp7wyP390z2gm4mhwpwwMq
tJi6iSbGm5j1UTcHL3U5SKXgzIxGA8Gkg5bPjGnAkws5iaTXvxJlW/H4Sa/Yr1R2TwmqI0x5PWlW
rUaZFxqI+b++wkC5ui2VqRPI/JLYNTv+KNpEDoPx5Be2JOeUZTf4UjFjRLT4eZsID3jR/qFJVH5D
vYZtZq6CypByN6/Iwyx8nQM+XrXUzkcTH5oaeoyRlfjE5Va/HfqAglgEpkVkFCb8+DADfhFDiLRR
tqef1vfI2IK9K2yW/S0WpSKLzv6tMrWrm4Jo50hTALSAp3TSrmYWmwqf9AFpZKNfvcbiZwRZz5JE
LbSsK6OvAox2qAlw1G+ELzB1R3l/z0OltrM7H+ZjXFTDXx7xd3Zvb3M+lTsuB8tRxxBwNOjBtXXe
qUjo9WORnVGEhXrvYFaJKTbkXl+SquAxpcPpiWm9ADcO8GAzMzgJsK4rLtnIAnhvh+T01Pka6ORJ
twDxiOQl/RcXpiHzrBtMT/bmobc4QIj/wsFwrlWNVLN9DJq0HoL6HOBKO+iXCRl7Kk2Ad68Jlolr
AW8ekEvYnKRMTQEyGtTx9+4W8B/2UY46KDTN0V8aCK2po6OCk/kQ4p538t3t1nVWTb99pJD7JdID
VmPsvFpV3Braz1SrJYe8kyfgOAorZ7nHLyygk9grlISkakw9AYAyUYTlnR89tbb9GNscnRz5FEBn
JDeMOR0bemu7sLsRI2Ug2jXQLIwQg6SfwjywD8t2FD4uHpSIUihLVgbBikkxWe4nF3Wchml5tdEi
I+6vLbOpLXBlbJ5Ga9sf7uf/rQ+RJxh7A36VnNkZBzfA7vzCM5k9UTEwkDu2itvBFfCSXXI6kIAa
n3qld+biYR/MZ1nKAEFAcVhVP4LJZiVi7+hJyxNeyRNwQhALRSpQ979zpMyxK0jaUI9GhzclMejB
MHEwlgbBdgHmwVbaOyBk8deJGPASUefvb0TBMxkIqvaGPatZ2NiYOTuruKVnzdXOaOBB2qrqWXPR
+DxdjW8M1oYzw2klIr2JCbJSJvrKPHzkdNANjYrZ9jVY/CP4NMVK8hgp9x0qCgHlrkU1FhM+je0n
+xCPUgbfI4gPES/TIswEvs9wfCbZyge3lj34S+y9uMMV/Q7BeM/YLCaACHRVs2LnNoUcqpxq0WAA
6950zCBdl48ObnQ5d9skYLNVwBrq6HicXlDvw1QV8pCWTUiszj3Om3NGfWwVRBtIJN+uSgSKFUYC
wXb3d37p/heStWs35+0WXeJ4KCGGEnyk9FDRC+fCKXxyplttLWjV3sFkg3lMxyclanCZjhg+G8l+
Orq0Id0hej7OYuQhgtk51Zton9H8DcZi4trutcItyAheReEaSVGYehN3/iGdUtrNOBH8AM+3sQap
BTA/g2VGqQdlO+9pBSiV6mHvdYlx3UbNS2pL5UutMXRLq8MBfXI2x8soyfggPwIAvbkCBM85ohh+
zQzrBRWc+oxfrYuz2eY+nMnsZzdoShiUOhSUJglaRGQNusEuMRY9P3DTWkIUSJoXDTlen9gtnOm8
b1892HdB7PrH0lWtH66fe5I+h5BWI1PSeQdE7Egt570uao1Pz2g2x6SK3DenQce1PU2fparjjVYA
Rfm9gHNytaIM63MeasA9BCAWEPuRv5DeNOX5jpDOQ4MZl2rG7S9c2mSd2YilQws7EStqOvZhJDF8
gmi8T+/+Qb6V6oX+JWrrQcewpqlVaByyxNem5Vh+Yo0pTA53oXlxK/dUVD134VZkwxUuX1iwRcf6
l7X0p/sFZoEL6XOgYb/N5Z+SLQGfbAZ3vZNIO046OrWklng3NRTbJ58AWs+QdXQ7tOtmOV9fTtCb
4AeAEzqKpOeFJ1MjaphY+Nv4O2C6xGc8W999cajFPMm7+3YnVfCYKh5kFFexz4Iti8DHlcQiV36Y
UYvxfRH4eg1QKipmCA0rE6ziSXGBvmpPganGZ1lGg3dWlbUbv7adY1pNS87pmt8uwiXf+BNTyDZG
qQ+3DrHcuD9muR6HT93WfzNx/Qk3kvo9OotdSBvIOpLbIruITS456SZ38uugX76cMJdv2mcXTFZz
s+mz2Yzo8rlpJu6VykcgX1wnehPf+WtFXPybQb3gvsvvl3KLQY3/SQo3gq87EBE/b6le2372/2oI
lbfje180cxzxYRPEiYiWQRfP89rQNtGzH9QeEAFt/OFelzuaSrYCT2ivyh19nf4Nii5Q24mdGMc5
xUqT16szs0QdRVoBByEsGkJeQI5GtL5lARnWOOLmIXi4HVYy+v012NGe3jcR3t3pHNJyr4zDmppm
gBgjcx+MFsJxi9N40utOYUSNgqMz4y4Qgyivjuj0EVh9AFlmv753dbiMirwZxUwjLzYqbyp+bEMP
eavZhSJNU3uBBWh6F5IoR5OPPXUIBpJOA2AXgTpiokGrue//hkqyjUI+4LCoRm/QL0J9SNa790n9
41Fup1odeIUIrsb63UKE17885bntQ6wiWRoJ3xixkl7hwn2jSh53wJxDlz0Px89mQ/lEbkg0jkC/
SzLgALL+U10qbNagGtCRwQFjIoinDnSPBx6WcBtr41iWix4uUVsdZkG/ioRePM3ZaM9lsmJto9H6
1fmL68CoFlPghHj3wLyNfm8hx6/VaCKK+xDM1MAu5AYVeAr2I8OKkAStIz0Y6Ot64plj5sK7sKwc
dk7ZNP4wiQ4+cCnZcGwP69+eNpqMxXeWBqhUBvqbT1tQf9wrHipI5PQUo4V/4BFFbOy1DeQO8CX2
Sqyu0AK4V/An+pcjGUQDG9mnloNuli7q6Tu6Kpe4JVScUNp6pNvbyBC/wnOUg7MKC6D3+4GRHMKS
891fk3KeGWzChIX7dwytQpPzoN8v5RYeuhxOxfDrDzlqdOhqWqTHOPuwg/etCX/j9mWwupWLRVOW
1ndI++TF8oQIDNkffX96vcI79jnPxd3MkFhnYphnwUyYuXiOvi1+GjM78bUbphoUAAjDXaQeC/Z6
96d4sFseTpKXhsJYgJrrHbHTpOCeOnatZXMb9EaF3tXu5/cw+SsF6oL96zup+lWo6bHKWrubaxGZ
eGRl0Vzcu2Gwwpzm01E2wIlJUgQQfMxiRHh32XZsAqQ3RmhcwTTAVqTggPMe3JemEbswtUqpgaAG
3dWpa5SyoWGvSrot7gBIy9QR0rOsF5Is9A7gajhucDwAddO9w9zmMd0tYgxAu+/kZogRerz9qtmG
BKI8JWTdFSDPYEZQv6XhwdN5nkQ65OL4VVDBUE1GDoyw1qYR/VYUDg6grU1lhhe9R3uFRD3DXdq6
G7V19GXXLGM6kgE2dkCFWli/uE9BkcruOrvMlIJlwpxabNuMMi7XwaB4//f32Bob71meoyqfkrxi
xURuNZZJxrAOfkWS1jYqS8Fx9MlngStlvHuXh5GwR5FB49E6BYcHNw4/0zdoukP2cgYNkoGhQm5A
ibtMMRcdjTf9fack34acMsKohaEz2XPdljjBywhXyoqt6DeuOi4mABONkycjITnt0wpf+xRBbRPb
OsWiELedWaAzX98ONa/xixQpOcwxCBFMUZiUkTIqER7b3GENFlA9NmmL3Dk5va/+czZbyNZEl4Qv
ijFkv2Dzpzo3tCTAZ23uwCJ1D4BrqmEY2M3Smeg3Nq3g+Cc8fUjOh3Bh7kuys/y3RlJYfhWXHXW1
18XDgDWJxbtc4DbWooNBWBD8vapYOE3uKAr9J+8FepoZY0j3RLBxWO31eCMS7qS0KebrBLGZOVq8
8PQ5PFVNFQzVpJ9dhvTXN9OQuij1vW7ZOJ+Jvx3MtVrLXfWCRsK4JySu473WU/LZ8rrAucGumJfd
jXta5D/Fsk3TMtRBc1dPnQu5s54j679bzfHg6sw/+7jVMGswh6lqrYLiMXAX7vonTi6epv7S7X3I
7KMpWNv8lfdHP0KqTRtIt2DW/HK3NCY8iFGWpyrWXdpF16M9jhgs8FoEMrC0FfdyK7hy58kTQcVl
+1t0PqFDuD6fap3d2oWsLuvBs8/uNE4gk4/Imh5ZYhbj74C73LOu6FPqShiQeyHEj2Np+9d3t4WJ
OJb55Nu9cR7gd+P3QxEOZhg0ARLYUGYVmhGwjOGVRyWHjcsp++OZeK0dWn+D3PHChhl/B/gSzGpJ
cfOZEJBnWXWxIhPFHeyDs0QJmMaKNn/fasvZdJr8qrGnP52Uquwjz4+OfJDVwHd9x4q/ZypPfgL3
hKT5JqNXfsBIGfbMZCYxhBNQ2XtMReyFyDzu2Ge7Tm+/k5yCTmB8rUDx1qQPRN+dyLcs7VvUnHJu
9y3tA9K+Zo7Vz401C3ZW41+dJgAxPOB3duSeIuJVJMY0za2OFtBZXVg6t28Oi5cWDsG/p6HcF+pg
L/RJtZELs4VYB3QQA+YichfNehcyz0M2AIO3EFZCVyjKye8pWJUCkMnAOGFxk1Ecc/aHw6XtZph0
hI3kTeiahepuf82juhNqlndB1fEioag+HoE8DZne9ADlXmlZSLJMrB7ki5dtPorZI/jAITC80XfK
Svl1wxAYptueOKaUjajihTK1+f5M7l7r3PKPRVsIUvItI7LAyjCS3nYiiYtZW9nCWKC5yIFZRjfG
z7sTHD0PgLxqmUWykswznZF2SVuqK6Gaf/L72CoKPoU7OMBmCPVXoaGwY/NrQIr27iOEHhOZGVu3
NUx441M60/tvP/5JEMDa6QHXJldxQMBPzxiedKXHPMVjCHgZsSiF6gUZGCw2/mmhIIk4y7cFWiZS
rF35LUGNjl9mFjkjYZ5hoZotCC1lyI3fJy6R8FAAhqlSm3VB3989GzB2rIKoZeK9FRbMFWSevJDH
GxUNRoY/vrR6CslVr4cpuZPFFRziwRm3Ga+hLmlbBnbVPf4LBmGNpYCyDWmoRTpqMkqkxry2AhQY
Z9kPJBRle0HJ5IyZAOcXsj0Ef0lwIerR7//PKNC3Vy7mM2NEMehthfAzBMTBfR/ZMrYW1xG458LW
Eo2ceJeE4xPGdcy2tV+PFY2sSYvfX/y3Eb1stRGx1Iz3gbbQl9tjy5D5LZOZbFsyPUP9AWQtkarp
vsOmI2p37uYNuQIHBZD0+xZqSpUYdE6mJyo5khGdLs786ee4jZoPSX7QmOEi+Cpg7XX+ue7/bv4b
V3z8f8sCpGQNqCbnIyrEFHphlWDn+ffDh377ImBXBq0WQVl10X5GQ7MrNl83DPsYB0it2JsjIO3A
uIIBujmpxgDUeszrq8G8MBGCvmbbzlYon8o0zyFdJAF8Ilc517P2MSM1VzkTtCgbOTisNbjznXCf
Cal0uJJboSQ9iWMz364lS3TYqBNC7c3hxAaFK/KLuHFJyDEnspyTiEsYqaXB697fvb5FvnD7fPCF
0FeQmOa3SFmEIAw9JyE2IuySE1ajC3ekMny2GQB/rTTEwwtOy5qm2aqRKVgEN1LAIT4dUv133hyy
tY/1AQdn5ZpbRRr4RtX3wHSoF7/+VN7eSzu2fRJQuoUJ/LNwD0TOQ2o8x7p8Jx9XgWEm7iPF22RU
9MPmhi+KpalSloDLNZolhUEBbxo74769G82JPfPnMIhqv2SNUmnq220RnFZkjZs0v914MxF9DLv4
ZuYRbHDSC5+6j8fAeZYh5RYn1MTAA9aPkpMf6A98fSPHZ8GYrEZd0Q5N/7Et3H92yv2sibUQhC2r
vfOmxqqicvKwD49vgZOhou/VOlc1w3BoXWeN5S/RkHOJ49l4L3U6+sE7KV8qcedGmxETptxfE27B
ytJM1/1ltzW+izgLxdr97EKWyU67x5yLP6OngJeGsWzDcry9srGNXbiqZs/Dg+DWn6gF0JpRXom4
H3bjN5FC2o9pnRBebdEf1WwG6dcslxiXgtoT24kGv36bH8syTsKohbtpt1tgd6/LDpEb/BbkSXmd
6LVOKeGpgupT2pS9jzHAYCy+vlMX/Nf1/UoCClavMT2whxtph0eBpHTh/nJxUmibvjP4lpZKMkDs
i7JcklTIOn+xkd8EpClW2A7HtvGdWhgT474DVPN5hKi8BG5Gmn1o28egq3QrpVZ5hXIORhZb7ce4
F23ZBkdoQ/vecMfvDkwxv1lt/KG/+d65lZ33RdrSQlA5U6ZbQhuj8um3bMmuA9tclKW4hbrAYcMQ
Wyfoel/OymEikaKkvLDqEDWd4UfrpfX9uk7Xfaz3XnRt1gF+ubikIS+3UwBYRm3LdcOYuEvsM5b+
22fXVQfX0UkIhkdowFi7ptKoqymZ+civd0r/uoOVC465m2LLHYH1RxZoIQFTXJnm6JYTtxy+wRDL
P8BxsUwQdg1ZyzaMDcavYgNjB5jLC6w9/TRrWOWUHpg3P5ibLW+qbCisC+BVCGA35h9r7d0a9S2x
T+NWhU9xOYHNgP48J9beCeidDOElkv9kCfLxmYwzxHxUVfWv6GzzpLrGlKBTb9kLRWumqvJxevZR
ULIE63HMs4lIGHgs7vmlA/hFN7oePr++sOD/PFOJf0hnV7O+3UIvS7EvGg3h+pCA3Eix2hQ6CYGY
Sh8p3cI4tH82m6sSh+KQvbSPXxA5CneWYuGfY0nuGAv37Ff9R/Z0YjajS84ebVlfSbYPlgtarq+s
YndVx7BdC4vZGp3/NU7uYJZb0/lQ2WrH9RtX7Cu3v/TKsIeM2jFL28OxbPEs1h9uNpMbAiDPOdSh
Gb/7AdVO0m4dblSbZV+YY6i3OoSar8a7dIcI4044GW6aNtE8Hm4HNv9YJNAxQr8uqtnxeJD0suJW
HbSxdr3n4/p2QRZm0fBykSPzLcM9kJMOGWlOUlhrVUGIXQfC4wXj7m6dKS/ULNFZ8Wzl7KGd7LBY
DjsV4npW34KAtO3nISJ2jN8CXiZvc07r78oAvplG5fWstBeSXLHb2jfUUGMXwkpcewXdTSTUCLes
8bbK/VeOy7bH0gL6Tksl2AfimANW1Ory42GfU05kCQDmeKbs27alz4YMlxwB7bPROSFTIekJWpK1
b+WodTwpHlE5OcNnEE5I7FW3TIZBdDtI+ocKkCqPAuBdmOA5LQvdyhIBuqxFSDXucFiZTVzgOw6n
USgI9prk7WmpyJ9XNjp4ryJ7qIrzJAKUoArcCkBDAO88F4Jl9ejQObfZp6LKC7CB7AsqaSM+OBrq
oI+v2HoyooXWT6VBhRcV1pl2SiMfeA8vpLdiXxNbn+HoG0Wagk6gGQ8OijNMuLOz6z53MiGggB7a
A5RUh8rRGA6mM1YruTpVGdiHqH0JumwZZVm0t7TZnyH3pV8Yj43Oj8I7NwjgCeFx6jHAWJx3ZCbm
juWxxlCar5sKFZjo/SdkTR65usw/CfpYjMLjX+oN2FlxDbovnd3hV4rKrRM2AxQwe5oi4qcedpP2
BCUjDDQwqXX7ihgCI6LdOvfA1oxtOrKfz9+Y+9Da+uExRr5Afi+72FHgn0T+t5YNlc/ppGJ36WwF
L2Cs9Y0Y4cdvfnW1sHROHNPuweT4+GdoRvqRHwKbeNmmfVL2Aw0ItrRbN1cBcw5yh3hOG/FxizvI
MYj9knM69UBv49XfddT/9D9djDyv7eOrAYvkYt9jir2xgXGcCF/En4VQr1Z+hBktTH+cNAcVOHsU
ZrD+vbg7+qSShYHVY6YyMzIIFOy29cwjetuWxJgU9lYwl+8sU8N4gwO72q1VW3Hx53axHzHpRkAb
d8+cDQ379hDCExK5MNMtaX5AkE5vHPWdQ1EjuaXMXBtR/eBPGMC9+zIdONrlduoPt0tW6JZTVG+6
QIxgQZI9v6jB5Un1d3PpVB/gi3iRU0EWarnpHzXUuzzb5fPzAo7qN+kDyBMiMu5UXdKlglG+6PnI
eM+WSRMi0i4h9iakAF5mt9sNM8Dj/fNI1Mx0a1T6LGCatKcdnHoGlOShB83qzhtW/DPIxwB0Ll5k
Di3Qst0ptT8sYhhgajj1BMJdFP/BNO7OuQge+fG/2Ocr+/TQ6v+q4PegPLjTKp/WrphowbVOUdY8
pBZ0oWRZLZvumSed9CS5NB8dBU0Ryw/xDt6nXCZuZBPgy5G8mydU8hy4iSoSYGDgVWWCE1huwRki
s4GTtEU6mgzhk/vG5RSrKy87eyXzoj41Q6/G1IvQ99iQPNmymgemZS9CZ6cQIlpUYCkoqMDbMsr9
EsJwEq9SzGrBGdZZNVGrj2gu2gd+xhNkPuDPxVtSDyadWvCR60r6+rdUC0294ZEgNLC03WuodLbZ
Cvnm0Hk/vJ/yG/ri9XUOkAIsKBJkRol3NIA4qvuBzAk08C7yHFT73qEAbNPeWIlYcsx2jlLUVBjG
oYn/Cl/Jq5I+4J23OD6CB1f91Eqmw1DD0aDGCLmmH531+vZ5XOvFN8DOgQ71DjW1KrCfIzwFDNRx
UNmkYV3M/+2Msu1rOzefe6OxvYhhomdJdnWO3xLTYt7voxvDc9PAI5RGWYaQltfw6Jrzj64+zCxo
/ouQl7uMTETOhjmSOav9UkA0JQ7hzz0ebhrIwayiCiTGTu6ofJLo+l5DfkxShhB4nkEYqDD1Ntmf
mIDwU1UItCMBAfPwwneS0ZkaDJIEAHxtBG7Lnns8tbvereImqN71SSeXsW6/LU0vH3NKqFUh581l
1JLYoblskwIAHoU1qhFx6EL9LP3HJlNLbONPu/zFyDjqwG6/aFftF689m3PqPfAuytinQoqAGNLj
KZrnkKnCb3tlQMiIl4vTle8xcZh03Lz30HvcACVsbVhqwxULbTWSH7aWtNM6bBmRwEOxHlLGgqdv
9W6613AEGTU+KIXEKGH2jwAwkSDWRGWEo5TImeb+5USbqhLpmV06D30scxgAlkjcxpjv47x+Eoqp
aCV6ogdG6QkWnPhd/tGI0EUuDHNx+6GijztbWpAEAlmPEDYcrZAP3EvFjTvqNyn43BRLnXLV2Gvs
PKoZeccaiJsXOnt14K0e4StXpvS88XpmPNSff/Lu93ag6CgZhgRNnZJF8Cp0mhOvcnYFxDDZSTrh
aiOzv7b8MOtky6RDf0n60vyTK2OEY5teW5nFHU0H4goNuSk6C3W5gdQYy1Hz0SfXVdX8zzXBTz1l
x5ayH6HjmfBHddWBX9zm5UfmPR6GKMXbjRX0COzeTVVjsfDiVpncikzuPJkvoHUM4ovAtvhCLmLt
eZwOASzdmyh/ZmxOrbNLeY72zqLC5sko5Ah1IMDVtfqqXklVlwXDrnV0WyouzLyOLeZIrUacwfxy
VN/LnBKbadyM0HmMV7K88VpuCPJPlPFNMpLjq9Pp/IE4qflWzeckFntfA8tCr7uhnc1DykBy0W9g
LOenf66JAeepS5V+NeHeitoUT0dwrXfLsr+qN0t+n/tzNPj3G7BjX3sYpgAXUP/ibLOjTFaEwA/1
gjNXSKZUdcnThcHpyieNE8JclGcjm19xyMkmYaew1KhO5QmO6gB0TSLGDDj2uIR91vaiwO74aX8b
nkslqFu50bvv+PuxPUuyZYMac7PQ/p9NfsJPqELNuJlhHnM8WfzZqxuGOubMV161npjFO1k8Akcd
lue27g4c1SasFiOaJh80XAk9vJ+xuELZ+4W8bWZ+2U3K34Vs5PJAqd3T1VS2MK1Q+9mPNpCsQsQT
13wR+31m2irY9kc7rYMHH6tNF74hfCmuk65VyBB/8Dfid09p27ibevX1ja7Pd7A8tRvCbZVi77a7
4pusG6z9zsl7m+nDBc7HHWzuDDZQ/jqPXYYCirXo9OlZTvIrnjRlTxegf2rmNgE+aQDujUDvUcLP
i2RgjIoYnOXsHMYSuuWUBlamK1c1q+HcGHUoePKy3DEuYMkuoA6iaE19eT4uIUbbN+Xa6JKE7luE
YsH+bmyYu9fTM9ktTMVgX4SrKgsA8GHbYmQZN4UDLby/Yf+7owi/7/UC1TiXPhXhax+V5OgtsUV0
XW46MEsN6HEKEK15bJgXRYV6Bx9ZFQGNU+M+YNOhBmN2tDKVhT+EVa2M/0QoZp2tj18UifVSK+Oc
An6yeSf8cVEM598M4WsfaIPPEvt4il0st3JhsyWnAT/jjJXK41X7u823MwPfCuvj0hN5hpNMOPlF
ivplivTUZSewjoZMn1mhx4B39YHnGFu9dXqmKicQIl3FaMCXomqpwIGlX+Hc9mFIIRGYy2cncQaQ
iZAuvE2gMyFeTZ2cf7X8PDPLF7eqfKWw/+OZ6DKJemBWwWyGR1fEjuhDCIPTd4GcIoa+HISHHBTO
/RkyAExVNLQomxLiA7PW2w+pVvUHF6PEIRqjAvHgRuUEmf9whpNzbPlAG0aRtTYzt4PleRYAzuIA
n7ttCjCYTNsn+3XMjC/e1fMJbgd65yGYLmNlNnX/NQi8kyAtCZNgV+hQIFdgI0Wpx562ha5kENXB
ceTlPRqRIvMdczzT/JeXOrAt8kf/yOoR9sdmygqUAWf6SXztG6N+a6HxwAGKOGYQo4ZFqfeRwym2
s/XwCGYnLhqnngXnLY4JNXc0GzoxFZdKh6X34uQYybomcYFEdbK+i2eXTdUxiaAaiIGH/RdLQkny
z7pPRThMq5DM+tJXyC3iKvwO1++EURFSzGSqEWlaDTeC3cjX0qT85b4URSS+h7FX0xaJq37at+QE
sgKIVTKRzJukEL95WzM9xTIMK7Gr9vfmj82L6qHl3RrFl0o+2TL2a4NS+5wt5GQFzU9pU6JAsbL7
F/O7uTv9sPfLpKQ+6nv2qUuy+Tb+9EkAANU4S7ZzKr2NY+hGbBIjg96BQjVda4Rd/nu5oVspjesQ
tkrr0RH+Ee5vRdPvyfmsUZREwiTHbI23nIbmmCmgm8I9ZFORwA7eHDeKarLY6k3J9ZHbI6RbeFCB
R7yIuGEaLr+ONhWyOh0/5EdpXfBYvCVMNNvk76hcl8nURw9U1reWEenSjXgO6Z/YYIYYgrrv60hZ
i7ogrfHGGxvf9xKyJiE8pAhbopg0TqwzWs6Lb4hwReV60/5DwQvNOHe15jbxP+2mEMwGTpyhAWP0
Q+zDd84KhFRONk3OX2X5UhS/HnCNA+LAKurZdvVSqu+d0JrRo146aP3RcLbEvUO/E8G42k8rSV2W
4fJ/mjwceo0/CP6SJtu8uy3MGpfsMsBvE1o75slUByr0Geegx1dtwPnYO9ms0miFRnJzlqNGffSN
iBXL9QEsiQ70/TdXRyLXpnR/WcMpG5DZ4jP2rvmUODZKBl5H13MaHQypLmEGmxm49MALZK7q/+3L
cBWjY4HF2Hw+6yznsFlSu2FRJn/cBLqCJFGd8ys8SKjlxhF6N/rG7e0kOSAnYAgf6y54eXn0UO8P
v5cz4b8TDL0thv66PUgXnRZYqfVLIx4PKMrBT4btC4ExabXJc5S+zW9SknHMk6RWR+F/LGcy4WLW
4XH+h+a+Ea5JcQhciKcgI5m10OPHDtD0JWh1F+r3YG1XUuoC4ZNqBet/3kXuT6hmO51l7LHcAeJx
HB9InAycn3AECO2oT6AZsXVwySO13tYb1uNjLKAdzpOY6piQHAZNuRybOvNhFoV7uSnOg+lT965o
czMRV7M/B07oWJkg+GBNIHj9ASkU7fle5++id+A4XvLvsIahcjEnv68ULdPnFASEh3jJwmpg+nSb
Tfw1uC3CDQd6ClFyyvn/eJKLTl0HfU3GXt+MaOvH02+iR1MON+U9afAqXrB4VRUAwrTvcUu8ihND
Sbca6BwnuP9ckbbXAfIX3bWS7P++f02VPxdBBsGIWAGfCVmYoz9DhhaKRdfmn1/d1EQlq+5+x1E3
u512hfo3bl8dMGZC874Ewxx5nPawJI3NLo3Ifn+3nErUl14UlWAIf9VfyvTPo1ZR1jGiE5CGe7TI
lOhajVBJLU4G9a1PPyzAOjheQsfF6z8Y/nlcmx6dhVaG4Bz2qiLDYSZXsquE5PJKHf1eUhvKFTfT
2R3R+luey5HfZJYSF+qbifhPjhFhpjIioq7so2a1KqHnDI9CC7OYKCD/1gcfeUfIlEqR+8muwkZR
k/OOOg8b1QB5ZJg9gycOHzj2tfxB45SGQWDxXIJgkZTyCE+amtTMJi6lOSO9OlK9Krr067C8hfNH
gDFGGye/lk2/VAvYvlpW/jDGiXEtMfMsdAg6Z2fdJ03q6c8tWN9wgGJ88oVkpiQiiS/P8M3IB1S1
va1+JERDn2+GC8pK75b2NOOGSACw7EiXs1L/Pp1w2yvSxmgrCRXIPWIoJ4Y5Xr3s0YswMpUD3/o5
A8VKHbZ0uaAfaEsA12gcu6bXpxo9mzzfAUVw1xRKngU7m5ESiM8/H6jhKifCxLruv9Fw5qnnDhmY
7XgZLyD5uM7IoFw7WyH7IHuaSZbn1M4NhkYzV47a1CVkPaoCMp0MOo2IQMV2j3kD0mNq3v291f8J
adSNXPrF9WDRIaXApLtnl4mttc4O+s0dl5X0ztZtHhKJp0ZLclBA5wo5FXAe8iG+iOgrMwtgFyyk
lzmtRgcPalVTqFxNsT+d+ZogpMz+qP4xfzpOlZW45qc6J0nBaSFluUyve3tevyHeWs//ItpBtxcK
BiVvd+CJ28LXJ1fOgVRIjOMKWKbIzUqMnBkrwmFLIqbZGRAKrvlRDOTSppq5Xq6AaFPklk+JgXo1
isr0b6/vndtuDvd/dD5N0StVQSBaz6TAmV44tMGaI8KlVdNvckiPh/Uhdxcq4zDEd2mHyi3Cx/F6
2udUGnJ6MBugF2q5cNOh0f5S4BnrHG7e1nUhZL3aXBaUN6dpv8+zMC17Nka2IG1swC5ZSy5sV8uO
CQFs9giZ/JWlVCJuEXB5/F3BBe4e5Y6gKicSRMx0nRZedaWUlvwdnoQ6qteE80LhUR5GKKkiI9P+
e6HmAgTcTO1R94bVZT41TiBgMwkeJiFQ2PC/cxSCpyVgEQYWa2X877jkx79EbfksvtpVx2/qbVTB
BI+anZj8X175+8I2qXRvYXe93Jik3BL/5FBhN1kK4z92arzg3j29Lq8jaGLv0Jv3bt2ewOhhBIjF
5ZfjhrYyNpKm5y/rOj4dywl1+SwWPjVku8Qm/mqdvIyIdqso/i279QPSiH6emK98Mv4ecBCxQfEQ
YYKCcwEni4/+31+DyLUSbkOslEsOayu0DmEDR3a/rZSuYp0vt9PsslBUFUTERaGESZbLnrKhHeTt
ylzLQY1rQIiW7EINlD/zBleDG439msLpC9r99zczTeO722hJTl+vJBoJ361gu32bMdXl/K6d/2Kd
iQZCXGW0jdHxcm7LnbpuygU4UgfNWvdyKvekKHlQ4v+tMw4ApIig/skG6gdVi0tjlU3l8IBEJxAB
XW3qXJfzEvzcPjZMmoOWdaqWdO6xoPQgY8reWO9sAvNNn2DZ2pdZNdCRlo7TsjkBoNGnA+WIvy7o
0cTESCDYt3NILwuBwLLY9Opy+KebTQsEIJe04webeXxGgvPHtkcDv17zSUQjHbQdDBBzNqcOg0rn
Nx4y81SeNh2k11zgPaa+o39vjF4YSWxk3ziO9WiPeHeeKGagnd52mnBlhhZOlkBYD8DzcBWbt/hT
UdLJNkqdLGuHZBXyjBieywJFky1cLO4zsr0DJQa3JnfUbKOCBmRmdLErA5ohABiWiYNT75bvDjRm
JNL0sRK03ON6gJ9XuxnuUgIJJpLAZYFHu6LawOEh0QIQydo9tyTRiirGSXdtqrlW1AJCf6Dgd8Ls
BldMMtl6+xVM7QLibi5FmAmg+fW3QSHDm1DF+doSBNKTiDzI7bkm8D/QwCG0L0MS2R5LPNijOWwq
kEaqsnHUXQf5vPeoiyhXDpzbhyCEKWjd67Y7JJu+gGpeK0yC0GDTl5S4HV4WoDoo/tzoCfu1Ubh7
ZWiEIfiUdk1EXnaWjQGfQTFwKyMAphun0EHIB7jKO/L4WGA95zOYkIAGKDKD1dvUbEK0Lowdn0QF
i8YTzhslsbaEb1K3/eJm2yPFnE1QYcTd3loHZfCjyj56ShPqyGCRcu4pI7cQRMxVNsLNvFW3dQLh
JWCKfDbeu07JXo5Zhc0SLnHSkSqNkf5mEzOi4MaDCFqu3eJBAKndb+QPenjT751Jj7WPVqVONpMN
t1fjp6Pdn0OFFsKqTib6f8USXb0BLsagAz+OBQ7wWjhlSDleV36fYuZBgVgQ065yXGHR6e/CaeTY
b7iTAsAvjJ1rUkRcnXUcbc0lx9S7LaeCr8MkjSA7OlNL4Wh6PaSmDQUUF952rNgoKHUeqTL1VAXD
cKgKmaxtr3D859syaavi0P11ZDBXRmidsEIuq0672n1pnDymVyV3Euo554QuUoxsUr/5tSKx+k8z
RUjk5ZfZBrVokWgEE498p+u28yUz4s9FR3RbYukjOs31cFfSgle+a9slNEemNxlO1AAkdw9SSTBk
Roz3kKGF4i82Cp1Ci4wTiwjjomX4CzbsGHvQwwEchcZ/SGvTJPvX7R1QIOq9ceP9glL+u70OiQNp
+G+FEfDrnBqhggNc89ABTS/0nbxjFr9EGmwegE8ykdUZ1Huh6FCflFWr6Ri+HuCkVH86L7sNbhBq
hq8a6R7KbQuixN0sE0/koYNl0/cCVPmWlYe/iHFwRKLXGhmp5NFTq7tM3pCQIbrtsA6/SX00JFAr
o9XsqJvPDyo+wBZYNYl9uZlaOsoXDqsO+pmXOWWWcBPq8cF7fjyYO4f73Jus+bwC2fhFMwMWXAEt
P1DMx9joBLGmJMQt49xWvuDbJ2rQfxR22uUdqlu03DjjqCaHLf75ShCa7z8GT4fur61xbIIEuXDA
Si6fHgY1/V/FvMa+Hy582UjnUZy56joR4Vas8pE7/Np3Szq6ytvnXtdz5y/4SnoNoKLVIQpIL/zG
nvCIMKdDVUXTnnDbecCwf6uTHiX/MKpo6oVUfnRUMJz11bp9XbTKFhHqG8PtDrkszYc2TxiLQ2mf
UebCrm8IlhyOjAlHEuh0+AQuYkucUVJgZJS+pbNBsOqgL8r+RbxvlcpHb9CQebuCNbs7XeJJ6qme
M/UztNRoxTgnNrq6OCHhPJmqswvfYNw43/ddRGcdDzUyBrgwsVUNQE4nQrgQd0c9f92VeHDDtcu0
hAKl9MD9zSXKCXnKkuyQv+UFiZLAD6P/VRTxyE6i364airBmhgqSEsc6PROXzhSCelZrOPZxgRoi
zJCr3ahFk685tI+rau2hE/kXEvm7LcizgNkNDZ/blZvJqpSt/kEsAJapTOkskFZqNmi/WPELKuwT
PaPxsFdbkj3yJh5ygd/JL9rKmsVR9CsG7kUiC4gfiN3Yzx2YBkuPTXRu/ehxNl7q+ZCu3/CLegyY
fzcBd+PQyANxiwf1t61Vv2cKZBJg90475yRKdAtmsu/mkmR/ulIt9xo+9ljz+3cqmQ7mnJw6GyIm
1DXpv5rlMhkENPc5qKdIM7/kyFwGwg5xVc9JG7cvWZ+Vr0mjSv9KEch5M7hEuaRsKEc5DjXFkUfU
4VZA/MTRpG2m0Utawm/ffJMp7S2vOEThLf75xQn3sWNrYbQAPwyTfF/5R8tqHteP92O7asfHxZej
P/kC1G25oDk6wBqDfADsvVKnwVycmGY6VNVSdPx0olRvePVywbJwldmeAhOTYtWZRD/r6N/VzMFV
O5kSuIZO18WwgW6cLXYyh/1O3NNWLO3cYJC+G6/H+CzFU+5Tgwz9N3isPbX5uaILubNLmZez4po7
eSuOH4ohwdlnifyMauG3cETscPQGPADWF+F2QNOmJBQvc521sA5QoxytOiJlbpBNJPJMiyM9xeTh
8wroBbUdJKsJsGkkgdLjkqHZGvgOKv338MKSSqDilS3I88xJcNQtqr1yhdwg/GsgEGFzQ1tYtVB9
W3uXG0x0MK9GbCvBU2yWg3U5GH/3nh+x0BVwdJBqxKWkCmsXafEU/AsE3RJWVDhLjtT66vHjGoDI
KgYiiq5fhbniR03GEPZgzDpC7QNhVCyNa0VrYwgGMYJH06SiELFzp2Gtg3qTxhVril3x+ZSnZERR
o6yVOzZbrAJV7VcLGbXauZHsS18WQWhtXx33/yvFXTFP1Q/c84BU+fMc8xzAwZ3mzfCpzegTviwL
zhjTtn9nl6MJT+2tzCMC6l3uD6bxtfRgCJtAv+yH3O+Qh0SkeWJfces6RLGdzNVtIGp7mE1+d3lQ
J5xXLU8SD2eYMhLmXOvnL10QFgFEAZ8P43CKjtjedr8tJSlY0ja0r/khWTnvzGYYT+L+ugj0uiE7
WeShVxLJpCTSIHwRnnuS6XIxunGkcUH4NaCiZBZ7e5sls6ObW57qbTbFVDrQ1nf7pyc5jOIiASVa
snShsSeZJA2lvZ+Pu+zhn64Kxk2hve/1tWdWGBIJzwEY7/IXAXvB7r2FSu7tltCChl8P/FIh+DT2
W9yCaf6Hu92/PDHnfCsKjSdcbhxXYg/yNKXcV2tw0ya7jiwRGUBMnJc7mNLLZBk1oz/achS58t6C
wP7OtJQaxYO7H0cOUMulKmUx6WjZwWz03XNGGFIZATyjF8iWWY/hJagRVSj5QbnBRqJCbVivz3i9
YsX0Jv3FH/TOAg0UlzaGRH5E5uLNgfmnkvuVlCu3YHn0qzTuapsk3yIgxzFbVLaqJe6B0g81AwO9
hyVsnySIEUJoPgw+lFnp8QVVNUMRTBfjcYorF7R5j4m9YsFrtvdCp74JCejo1CguwMbmKILV9zFl
He4mafk7IGyfArbtYAPHyJIWWSY05C/KlgLnfnAYkw2G5/N1XhMdJ8v8JtjAI7MSvbN5LwoyWvDt
LlIfu1DoEk/QJGCbLR7PIA9YZzJ5ohAneHxxTsn3AzaPhYq7rpwUy2o3RM8wigrtVHg94H5O5yw2
CsbgraUCmmGsx+0FwtPs0V7XCU9IuP6N01GlVj2e3tMXp6qTi6Jq9342WEl8xnSIpP9oqNJQoivX
5D4O6ZxkgXQAghl32NoB70UGOwQVqQpJ9pqeGVxmy8eZXc6huESssAYATmjNHYmSHYirhqTh7kBv
PEQlqq4Lk7+8WbQZjRNJ7MzyZEyNmYscYwjCTlRrLN9sV7GVV/S1VcpGQ/5n6iXDw5Qhxx52lLPs
iIafn1wWVD4kmGHhY7TmWeCpu2U2c8JeAPhPjFGMyHZdWACCQ6AuQYpKhp76u7VoMV9Y8f4mLdS/
V4fLhTZUB118qUgm2l5zspHPnhvmLZa8O4BvXJiCoGs4hxlxfljJoZW1IwQmZpOhJ1QCj86m4Cnw
11gfHebtYExAxCHkJxV+jHgXFUzm752+Rf7lmm0cdy2rNRk56dkgFKSsJWPp79Kz6JiEeVuoaeIB
3FipJ7DeYPedmbZTT9RGPJhvv4KcRRoDIncGTtEVH1qn+AI0AtlWjgFD/I4YtBVpvfHMkFo65A15
N32Qbo1SoXgfpigzhADat/g6DTki+R9UsZ34IEd2PKihBtuhPmZyq7gavM+psusuN+as4nJ8dSmd
zQPWfN3VWT83LwFBRC1OUkG86mLc4it6VQAnXqU/ohkxdYK1yB1l4l2fucv725yDnSA2wYVW2kUm
+m9/7f7aU3ii6CvefTjFSsIJVIiHhlSivIF8nbMzpkfw+DF5WzAjt3BDgSpxI4onNWOT0mxrHuLZ
Ue2RgCjnSFcOKefmo/Fno9lJBoMy2sDO0PW9QzsEjS1/AKWMuuwsImjRbAEO1eSgdNmy5KDtcYE4
7BIpYMJh5v2foNQhnmeovAN0ou48sIcuTraqjrswphGQNs0bcVDwiHRctZA8EzUVAg5zuPSiUFM7
7ljGIH2xCUasVmd5McNqMpV9IskRC2VwAxaFBQOgwQuwe7tcdO1ePatgVatxeosEu1VYCuHCgJey
Vkzg3qu9dwY0Gs+RqmqPxxT77Xowq9A6JxFN4O//Z/b5kci7MO+QO3GB05GmLhJO/Bt9AhYFIzJC
tkB/39442nYoSgVAKGX4u9fFW01Me3kd/81Nw3xnYU5Cq89BEH3adAeBL2AoDQbU0NUHg1tDM6xQ
zUncz08ZBzqZDJPeNOXcnRJZKFkLVuSrAj2X42umQlfnoCEpzdQgecbPeAPeFopqqJqsxn09J3/c
QWgH7wBb6O90w2P3qRWUwXwEyc+3JIx4D2Q4PNt6g+tr38kNL7W+W+48kHpZtLeko03gtnYI6J6b
8ewoC09FqQaeXBNAQOrfvlkT7fBtYyYg+SCjlVx6EoEehYRKzHSJT1bPX6bQxnxW9ktMsyRYyi4W
kKOanAOuPu72e1uMYaAo+0UlpeMf8t924FKxS59jgak0yJIb5e01ZiE049UJ9JcaWFTy+1VLRr12
GlouF33Wr9vJyGvFr4Y9FdFgTVj6z6kuESmqsSI5M485WkvdZtuiKMt3YJ0jrdlTwnLdZeL6B0g6
LI85MDRoFgtOEISvZDG3VdjW1R5NMuggq/yWkio05WW0r7RXo6pG2E78FRDIyeRLbRB7ew36luTo
jM5iFu/NyvQ7+5Zjt3vAuoiT0Fp7Du7nsi5wg9Ps6Uc21WVzFdv+0lKCqD6V+yJ6iGGxga0vsJsS
dXCZB1HgtsfdSrmto7R/UpFy8pykHlBYzurOyCmZEofqy04fppAvJzbvUBh1CwBY4+fArEoA7rxe
XrxqtyfIH50aLnIG65TrZaplQfCxgeEJ1Ao5xzSGyRpk9RjNKUzYJmGStygzPh1395IcIcOUktVM
Egz10JSXxMGxfAxG5G3ua8p7IFEUYr+xHQ3G/dsZlw3njnOh6b5SV2Wk69I/hDVqjAh/4SCDPfVo
5yU3n3bBFagRWImlY7VnHUwnbcsqRK812bO+AupKN9xNNhossJTyVJy5YDvGUR3SabEMSCXgNteX
Viyx9Ber7UHUPk+GwQX/HDCXUEDz7Z9sf24lWchOkS1ECX0hdUeD4xgpd/7p/ZXB4aVO3IChPbjn
OdVSn5QDf3tc4G3P8mzoqNAM/6aQxXE7HAqPi3Dptl4KufJjnhtkD7JHZGajkhk1z4xmX0tHPZJv
UL6aGVQsHyp++k+8XqSFWCcG9yYri/T8q5Fj/CpMdfng56JsAmVrHDZK+gTeoYpV22Rf3pX8QZA0
D06hj312wv2ypG0rEB2PPwGacoUsFlZa9OMsLnInlPhd580t8aVdjsj7S5O/s8NT+QNaexf3NgvP
FKyR1ppjF4MAZlpivQGg99jDDB7/gt9Et2ewfLLFjfPzSps+rijsC3FM8z1OVFA+30pil6duse3T
8ZaUMD8QAceB5PBueEfAhwt4m4X6J64OmNFJ9Z0PPZsdGzbV6FPIVksbG4U4qR+04buCavOjMbw2
nikub73p7vp9uVh4pPWHi6kg7qU0xWWQEVXPl5TWF+E7FTtl5+vt8upCJ3RcnXeIGaYdP4AM6T/U
rW6tKkhPOefmBc/0Ww14UIlrI2qO2eACwm/tHyS0FtzhI542Gz2PDSqtjFnHZz7f6kST8Fes5vha
KF3gW4xDHH0+WkkCX4WlwDXAw2SQnIsgcTQcLnoViVg1yFtHbWERp7nFynnB9/dM022igQW7aEIA
KY9BiDd51NxTmTZYYR0YgJuUIlZrrUwJSy5lb46E8Rc6gneqbJnnCySvEcc/Q+c9uap/tO/xKpwp
nexuTHZ+9U9fPL5kMWo3OaDGSysoum4rhFC81O8yJORgn+SG84iFYvybg6QO5i6qPwbSNcDNm6+b
AuuGlE33tzO+W78r+mA3Vf/x5wjyeERF3NecP6EFK1EspSuUgRaT61t4wc4kZqNyWmDucNKp8tLX
YP9ovJXwhmohAjn2k7w+/LKe7ZU25QO9wIr5+O3/XewL9R24cZKzg2ee2maO6rhsNHrdAvqd9BuX
sprgwFOoeLuU2Qf7/KpGLmf7pDN+LyAea78otZeGGgDUyyLjjzMjJHWU0A9GjXsXLRurxQZafSPf
nonh1d5iD9puv0Bze1eJ2EeuvJTD0csGxSExuvpZMnkp5n9Fq9v7EQTDP8CHFHbNAjfpOHhdfrWK
IPP28CY0oISbg7j9Cl61W9R2hii76Y7Nd8Y4fFZLX8H98//lVfEYVWB330pIVEoC8CY0nFUTYPpJ
YoPtaueH3uKHfFhw0iFiyaBbSHE6GNrQS9G73pBovUlId12kaExAnPh86O0V8otVwbKkQ0F7qT+B
ZVpC0VfShAcnrZJLYJc9tkV2s8PwGTgPVu7cJUYD/Unbkg1DZr1OmwGiRmgAOHdlMy/WljPgyVrl
Pkam/G5zP/LPoNMw5WPin/U3ZsqV2Hbg5011EBPBh3J/WVxyeqj6jwgLRMac8qa/nU3gRzKMMnYW
z9XQh53hVn/PD8jPGNBGJudUReU8UAnHn+viuyeywtkWz8lipAIXNn4a2rvLjnRRKA2dqsNJ2FFh
pl/nHvgvmgqLZnjd2rjtJ+siZYg2s+EGm1Gpvd2sz4EoQuKEQ+zHHBAcPMHGoVBtOPOzVNJ+2Xnh
5uT1+DS97t9QeBQ1cj1XsGhUVUf6uIfng6ZRyUjZFJwHuFPG1zdAfE2uES7V14hqRArAw/LS53cc
znFsEZH632gBMa9fKW4wlkYjbrn3TFjoCS/3J+gsLEG8vRROFcqimEicEEtxSQnz4U3lvFpHURoi
6/mVLEeheJqnMYw9Atk+GZH73pBztlNtEGNc6NQlIIkL+DoyeXOuD+UdYMKTBzOz7Yhyc4/nTplS
HbaIrME7c5cySvUrEaufz0Y0K36JKldkxnX1CeJe2GDAQ2+FpjS7OQoF09mOvt8yEeUBvmD6Ew/3
cfGBN/ickaKBXVzoB/hymjxYdh6pxL6ZQGGIs4sPRGZ1GQeymEUQRNZySn8sVwJ1PGKqITrp2glp
wafc22k8Q/ZR5cqtUfq6+Fv8vf8BIiP8bTYmnHgnPPQB7uCvd+pf6eiURHq3jdkIeTb6guE1JQrD
+Sb5oM7YzOT/2jT1fASakfpsxVLXAVIJJRg2IqMNfMnZIvd8uPlGd4CmC5VzmRk34R8DJZD9BmG/
H32NgWlA5U6iA+l/WbBhw+uWJ7ft+rLxlAzTaz/Yrc3FQ/DKULHCodrNTNBnkkyOegetuYt4ThhT
oSpBoTlXulz2yMfhHUjymZ6lOFfeV3ySwNmdG7WLvvY/OHsDoC1JC1fAa1Pvo1ccq5gJ3EkxPxdp
yRrHilqh3UlbvoBmEvrZeb74N2ivSBUcGGCd+y510Lmmzi+zDEhdGLb5zRDvrlov7qpLhP6JUfLD
TzFoFaFYd6n7HbqTxMj1jENHE4qxrrb6IW2UJAPo+ArRXqwkyfo2GpQRP0P1CXlOdbLhqjOnnT28
hTl0Yx8nl25D90X+UU0WKm4M+y6LEoY9dyVEoTpl520+hhQ/v9aBoKy1T4uksUkTcgvEIJHOuWZJ
OQyBmq6RFLcjMlH9t1DIi8bwkRMTQlhngYLGwnXKPO/ksRhW/ogc5gOv2p4VOygj4seLS+eohETR
ZZh6uXExK3jF3hmVpxNVYvL31ZHadmWXxmIw1E2YIPTs0xONVqmlPY48/gs/VFJNPZN6hJt07khz
ZUebAnJ02T2xHwRUtGdfFqqs+A1Rfe3o5kds9N0rLVPW+xkNHIfakGHitvclmLCDSIg/pREf03fX
SrdKLp6ZOm0yT+j01d6F/VkuJN/V9O8dvyO/ajxFytdE8Wbl9DMltxctIf+W4FSuB+IidC6WuB43
ZisphRItTq2FSoZS9K5TZ+pP6oSaJ+XLj/9p2vLfJbD2KTmeNDdC3KoAZIHe9rWp0+wkj+rhUODW
szZ6qskatqo0OFrr58mJHqsxNWaEjg3MX4osvFOfiCnko4Ja89Hq59g4K97e6NDzTqtfsy61X7nT
yI1WHlp5YwZ0hleHxEeZixVB7ZjyXPK5lzN3eWcfIW0XsdYCP2i3XG2Wq0iuBByJujWzB8toCV+B
5v0PEUm3GT1Y9vhrubC7F83MKorNDtZRgz7Lnio9dJsXoa2j8P2nN/5S8YpN4Lz1X9r5S8Kjg1yo
hrD9VnwQYevVhd1BTCTybvohHmD0tphOg6G6b+xKQ3TN+jNzWw/8YaBsmz8rtGVdxRUR32R2kwvG
OnHyfL2In/OJIyyyH1gYUvQiAQGqVJAAT3X+vZgxDFTdEI575EX4XGTySACdgpiM+uoe8U8W43qZ
4cGa2akuJjpVaTO669tWlKb6ThAXxQCuuqBLMDfbaFZRULBPyPBuhIPvLORw/BUP9bRhgk6kSn6G
FTNa3KXWiV/D2mwnx8jEYM9kKtcfQD178nu1MIXwg7utdIET+fs/iHBJMCvP0R18Z4dwgF1lvzE2
ptHRyqXcpYRstlw2Yz6VESQcxeI2zynJYt7tFtQkRmYk0N1Wp0OuBDBeVA6SGvXOOc5dHPkirDs6
EZ/GsAwWrsnFCSbPlZXk6zARVhrSHzytPvewaG6jpdc5Q5uADFIwPwYOeAQJ/PHcFiSdsqnY6Lnx
GtAzmzVLEv67qESlM2meKUGZcrZlaVFIiV6l72ah5M67791jeqi5VL3WeXeERkkYzoTs8TYakc6b
n6Vhcd9UE7vi0iZr/G8aDBW7xR1GWam06Zjjia+pBjFYkTcZeIIiSY4ZongiqheOwO+Hp5Tm5B+b
RIb4QpE08fV/W5LH3SC4OTEyvBIdcaUe3Fxq0MFObxtVaWbNkbyw2dbMW7nXy48He1zPdVTbL53c
J/NRvgxoYVtlChSXG1xbVlh/7xepFYaaWL5UvnLG8YldgIMj3uW+3oIrQis8G76sNaV0MzUP69AV
Hf5bcRGdkeoYad8mYx8pqg9v/mGcKQwcZ6ESUakr2sCUNWXegwFlG+zR7kn6oGbiXjX+GnVDjhan
AJzQuO1nk0eN1z/PmFoYqewdWemXr0J8uFXSOLwZFsonAeQ8aAwCogBx1hmZTUE+/aQIirFMWLFA
KR2FStqCq3XOsdZ8dPG0hZH/Z+v7XLvnx+LAPlYB8kMCXAyNUCCXTmFAtMQnhPcuJwJZS8aRmtm/
gKU56rpDscHzZjUeYMI01IHpnL6E/8x44ROt8lWDaowMemBTLFux46Gwq9GOAjnqYAf6tiLJt0p+
8O1fqiyoFgwT8CRFsciclsG6Z5l51F++hom/oHEWyoW7cdxVf/kS6xVX2GgdM3uqn+y100KEaXA1
YBM1nAWIIZD/M5g6SILsdV8tAOOrXqqKh7g/URHJl2MHLiI7b9VFXmPyJSOGvd5GCNnYGxrlOeac
IpDcc5hU8pDi8nitfPZK8dSSlCNFUNSDXjdv15IRfNIUi+uWAMnQWSXQ3s7iQblkJrLP0/ueJzq6
Ya6FhQDTbzoWn9N0J8PGjhsL0hQHOPBdWDiR2w4tNZZY+PiMOGEX5GvfUsaeOU37z7yt2KDmgz3T
MYsc3P+illaUtgx3qYYH4CTTOtk0iobDdofzkqMuoYPzhmJpRPHuTSJWnIiJZez+xFGprOd90J7E
4tW8w0YGSGa+/FYvnVdKvIhUkzwmsfwZqzdTlhtgnIsty4wV27wjRXJn9qOcyOnV5Vuteg3YSy5Y
Jjd1QNWiktjvdnupqYekRvWnG9DMGfsEbjl42W/oyd8getVpTA6BcEmy58tLdMt5iGYwYrSnAOut
7WFw1AQpGFP7kE3+1iA6Ow4asyLVJhvv0t5XuGno1mHx4Qc04nvq4/gkihgk50KBm8fKUGze+Oo9
xjOsXiLZmZ6Yo1LyAAmFLsKtiN57RvYdyocYGvcnOl8D2sDLjUmZWmNZWxnjhrGViui/wjMYw1VO
IkUdyMliMMfaTdobK4LzZLWWaCZOHPITf76ssSyLVfibvoLEEMTiy04jcUT8pFXkc7tWDYXREMjw
MEHW1W2ZBailuC2qV4yaxwhxP03bnriw6zRASfEkpAVtTbudbADF/+3hFfJr7Kgyho4ctMuqhbCs
FLPrFuVwGV8oTCV2jpSgHOfE4XC6lKDUbcW6viPrHETagBSaEgzuGllH4ztaVUw7uyY7RRalSs28
slLdulLZ8a5IQQ8krMsd50WKCdyVHQXAMtB28fKwqxrk+QtJqiRChzQ40iT9fD7XDR9Q9AXhnXKu
tw0uucFyo+Iw4l1FtbYj8DVRdSnvOQ3uaa4EhAA76ByXmzYGOAmDjEtLzmiW/NIdButN3qZN5zbf
NHD4ayunihGCjlgyWUmoHDKhduo9MDUz6jo4nyugKclnnYE35M4+jZl2D8MUvfN3Sw/9pEXfP9nF
OfnQ/i8nfN1XKU4LBYaQDOjAf2R48ojENd7UYqunavQRvoWhe6LoUTGGIQ3SKMtxuWoI7Ph2M1oB
Apg9UtWEuD0Jzp6lRG7DgzXuo9TbYvEREq7BQWDSNEcnXT4SA1hiwZgUfau9wzFuNGlqVB/jROj5
73hgUgyFLMZTaUH/7VPrPGaldYmfTXZ4C8qYfLj1vjCCxQb4WQFLsTuLcip7W1mu0Hu9FoK8Z34o
UosISonlL7RcPzJa1hVOGZkeN6D8azP1RQwrm+O0tKTXxdXjgii6PM6YboVz5rc/MMh6bsF2n3kZ
SdrjxfKV1QsHf/Gbtgy7xswCAP1XLdKKQ3Jmpxh6o6CTaeRfQEu9TIYaHtL0yU7dK6mZJKTvc02s
Tu8yyuUWAmdCGpgy3Z1TTd1EOhVL+h5melhaLfAG4XM1yT0x44BSis0JMlHk6EZhmzYCcJ6mAq8D
x2AQOqH7ff519bEFSpjoZtD7dFL4Ve0gS2ra1m2QyiTySJxtQrz2+Ay1QYDOHhKOHsLdkZgwxlpI
UsrKNGN3vQCuFFgo5G9TYdvYCmwwnCsVVZukdOQF1H0524yhjyVjxv0thmEjdkrmkINl8dknGJEf
aJ+YIP2yiWjnpD54gXOzFHwEsNMjURHtB+yxypN7ST6BBAGuZZCsAspDCBxgV0oiNx6lL6+LLH/I
zj2DmPthbNPrQYJgW9shMA0jng6l0Bb7WwKHARkzRRYHbC6ZwSdSynhIcpcT2J/3gjkiWUQs/JIz
lGzFASDXJUbwc5k/r40n/mixXN2+M27ThXgeXaH5LBXN7fHhMe7kZuCuoEyngXM7dhHoVnqEjn4F
+++z0j4fgTwRF8tcNDfM7Od2PX8c2NAA7OW9M0Dohv5FKQ0QjcQmwbTaAmOGKm+JFfamsF2owT2y
OMMz4xhgu/fK2Ll7U4eYjYMFHHq50v2n4DPgw+XQu3N5m+lo6VkWCJCKmd12DQPvggC+1YIxMzUw
L4kLnVoW81v7Mc3vIa3S1RfY/w4/Zh/ZA5UGwqnKu2zN5MBEjvkaMRK7eKP2lvuXlNg9y08s6xX/
ns2k17owxe4FysScTC/QzCBHFw4Zfz3HbbFslgduCLcrvQb4Z2tJhRP6RaawCN9UfASKEh2mO77n
cVNkHppXz8TOgLOWlPSEThPfeqBnnwARuJu28dinE4v8Jb0UVRIBWyyBpSXTWoievS18rSPlJWev
m1ocjnprN31SZIosVoIi24Nk6VpKq3ehRdF8vUQC29Ib6TnxGxr/E3iClhtdwtSUiUOA6OJpRG5U
4FKRTu37YfRmCf2Q304IeLrbG2damxckWb98wQavBCp81cWD9LjWHICam5SKpUOoBvMDGRBxxrhs
NHOs2+i7xkBl2g+/YqP0RD3vFhVbbdoJRUfeq4mRVBti751FmgLS8NO836ex0A7FLc/lsVKz77aA
cBdJcH2Ncgl4m31Fq0Lr+/HLqqDu0h3MdvwoSgzPDO51TwIUtyZSyXShUQ5CeZz4YE04IzetP4Wd
EdqJTx1MYJxODW619jzGuEPBaFQsRD6/YMa4PWNoqfe5MyXM6vZjjwd2Ksa/5Yq+d/K8wjOj8Ll1
ACstGhHh1KrrX5bNCAr6ST8zn/qHa+oG9LQN9s/Y3+KifMDOlGxDHlEswd0pZHwoVcmB+X1YoH/+
oaRSAlLKLU04PWWwW1m4kt0IAR0nC3aKtBAzr4QHdKK0qHdcp0aS0wPpis7R8LeuL3o+3BxQqhnO
Z5Tg4xCRTgdo/P6O4Q8vpbuPcSo00N8HN3vRVUpPYpOFGcaUceY8BDfQ09u7MLIXi69r83i/l19f
96Tue7V/SbjVvy/EtXUpqkKBARcpY1dov4PA5ENtlgd+aZX+Zy8N2sFK46oFevURAwAJDHgr8rF8
WfHZPUyKuSkBQHncndSjqo90dYiTPL7tamB9yjLSZ4i4Hh6Fm3qvlEAwRelkVmwyU8mwfoFn4bdE
9pI1jGhlfvADE+++/5cnpWUpHyCMXB/RDR/A/lBNEKrwQb+8sBVs4DZ0LqJciGoMWDept0Wqn02h
3xLABy0viBMqcfQlMyxYQKKlheIv2ETNI3/hk0sFpPxUvDEWy8Eo1RxCvR6kibBI8AOBNC/5W8wt
na+My0AMx99IFitFzrEhaY7Xcd+iRpnxhfP+/6RBF4/hFiRTInxNvD1+NWBP+PKfmTTozjx9+jCB
Su9Wj5Utz63gIZ1bbyzdMcf1Ta/r/hE65sq/4O4BCOv9KtWT16tg8mdUHkVsaLjYygJiyL3XCbBz
2x/O/OhpXWad8V6klNBOin4dpqoMNO1Y50xCRtRX6YKHXy91zQJaf3/i/nrO64x9G+BXMGvtm4Pg
+2KV2T+cqjDCbzUqS+JcfcYyPeSEQ/FrwpbCuzXfy0wjz+qqZ+Ggt91LOjwScktRp153NYDwtFDF
i+27oqKRrWMsNADl5/SADh8lPMItKIyVAnh5CGJQ488muriTQVoFgEf0i6mQkb5TIoq0O+WyxncE
b/0wP9YoHU+d2KbFnanilSfDTIgEQD/bsOXhpBPAiRPXS0zj8vgGrNOy/BtXZaU5xCO94aomVyOV
m1RZliMUOSr4AroJACB65Lwxhpj+1H/agnkT3x5PLLJnagBrbmYWoD79qvphZQoLPFHx877OOmy6
mWoZZI1def1rYs/HXIQGztjDYDaRe3K+ExSZ6RgtBYoJX895PFBh5jN7zr1qeX2Az9STHr/9MSn7
aytbkY99YNNo9VeRdIP/9f0z8UZAN17fHm4rYQXlc43KGHip4vXQ+cABZMo5K75DHc9GttBvt4X9
EArEAOcvFSsRuYlQqi4sLJU9k99fKlJZZ55EmMw2M9OwGwZBrY56NQ9Rx1WHHYe77YeJZbuxNgFK
fJqYED0SsMPrtzw/+/JFtUkdv86rdzen1/kVeVdolNdfPQkEdMfaAoBCn3T3L7etxPymzWdlZ0xS
vB9P5MS25UjNdQIvTdTtFLQD2oVQlSa+iaZn9tB8GtMd3fCeqheiNEajt5r3H1nu+u65iPhQb+QP
1JDzwUHtefQ8n1eNDzq7wnPSA5Imm9qSDHbF0t6TZPe0uy/rv3oLq+ywcBYtQfHQT/TACG2RgqG+
Nhdk/Y07MJiVlyVDMhXDQ7WCSOg6SteLuJUbdEAjsLL3qMhQbHgTd1824x/gQTS+GTwwHbf022o4
aVDWBkGAovpIYDsZLDhP2+00SkiIYXLe2XNzddXgMEQ4v4AlDJCDLl3c1fRwUlm30VWxAokgv/kj
Nc+t44RjbHceXSP0LL96qIaNSaImXU/up0myFQihchP6WOvnPwqPXcy6ZjAulIgcJMLIBJP6P+bz
OeM2ahJq9UhQLV3E1lfBUdyU4912pwS8BMizVAy0It1eYXaDTSRsHtVc7P9Eni0Ac01nMBxefz9t
xyrtE1mHxWtsT3gUQ6/0bmqF9hW5Hu7SrifUR6d8y6mF4fZ71UwgLPbqtcbekLNSrtn+SWtJgZ71
BKJt0h1P6ETS4c5RKRhCesLuO1OXkmGCa54bhjPoPe8jByRCYXvCHZOjxMYNsnMvA0JsqhthdZwk
hJVZ99mf/droEed7ljsX405DC8FQpw6CbVmvbKNlrB9T2iTx9d0MXcSf27k3ixI5ExELlGWLLyk1
dM8c3BXA/rZRqu6k5yipC0DTHS7POveARJER5jd2hj8zZ0T+tvd2H1Pr5K+hr8PJ82AH05JJDqCp
vzFxr4uO0sPC2NFvRfDeIBNzFhiuW8ON38NBVcSY+HQJe/ge+jBVoLlXA0XtMsi2LbmHfBSeVcgu
+P2GPIvZkpZSMM9+8vN2ax34CiugjY7wIQn14Dck9OFYuuyNuNjMuPWNkevJ1I86M2F0N7CqD7+c
fJRJq7RniXlypJ4nGqgs6a0ay69IPeBJcFxsA70vkVd10Swxf1mMw4mE6vsYyAnzsMWxHrf7cqIP
/99ScQX1RuOkMgLg9yj4F+8qCXd1Ig/s9yPMUKzogv6fbBjlZ4+VRev4I7OmVwg1oD3omLPW9we4
b2cTVcJk/s0+uyp+5utPpmb+CsS3d2aOoV+lN/XtllyuOImx2DJSHdUfMB4hCQDPbA6qDyUeuZfE
zlhg1EGuXgi4wtkvT/cWijCqGNDURp9yW9vnaFZAIlucFb/EgOvLwczBq3PpiiyZRRz32+KYJ+OZ
SUcrqzpKM9UunNrDnGXYZJtuOXhFq5VFYK9LahfKG5fE8akmQvWmRbwYU9Cp26reElDuntXxJHZx
Yb3rBt7tGAMgTY4hRsOipX/pr3zBfqOxSJT8rdCGoOJZJfJCAJBvKDRwMOur3CnZ7TbT/zA10jr+
sEl+afKwoNB0kNXui4nfuYFULfMpGCwzq8qrD3BeXQiOQy8acVQaPkIKaZoHfKXLkV4OXVtI5GIP
3YgcNs+S98IE8pCaMa/jKTn9zTKRLrhoJKhsve81jyuGcUAd1PQrV+leiy4aNRRnArsUZyQIBanJ
YzzRC9Q1VOOHM0uMBc5tdS3pOogjWs2QzzRP0lIHv06ILRGuvxhmowkojdURVm8BZlbQSfzD/mqn
9opbJnhAt5tkH5uG+K3o+2nAQBQyb8O8ygL1UZKwGx13z+tMvfpxvxw4HO3RpmiCF2DMhwjlsyTp
1OKnQWhttwhiG/fvC/U5FrQ2XYP71GxXuM6cJH2jOQnjG/FbWbfwDcEVolZnMhgDc7aTguE1W8+N
j/2A3+7R3E59F1IZ36+FKaGVd/7itxp4AysNCFuZMSZJIV9tUsuT0Q7s3kYYvMtvPdJXq58lYgcC
zhqm1jiT5T/eOpRIg/1WI/wBgEWQxcggpvhdrNvElCtvdbUfP6wAV5h1X8H6HOdA/gcTYwvS03V9
12+cp38tw8YZE5ngXC/U+f0u+4Q9YLVEGuKCOJsjeYCFHs+Pds6w5FEDl5b6dZsTIyTP71BfSJVj
+DyDW7LjKKHaDZ0SHb0xks+aWBiupycfdp3Bki4Fv53au1SF90cIkYD+n52vSnhUbqyaQhS/Vc9P
MNcc5E7ugHdPiZLNeN52sMlXN1/P56u+kq9fcDLO7EdM+Yrcyi4aRKUuhGyessMnwHcEu6XlYNv+
Ls3H5PDWUJN9VS6CY35eX+VvzlY/NdBN88PDDXVaZ/w4xbNUEVK5R11x3AN0M6v5OIyrgf9TiR8z
Rg31xUbjUhGJ8xkcHz4yHZ32zwvCX4QMvUBQjI0ifG4AWcgQJpcaCUvmGilN25XmybSkhvtZpMOt
QuqAofZr8cfS4AfVpWMlKBvJ3bXnHv/YMxDLZP9tYEomM/DKKzUuubBeQ1iQK1gmTzRWQVQp5DEC
/WXpLl3aKFbRHmOPtBe/uWnZL8l9NBLE2+dEKxzMCX2R2Kls9OFVjLWsuf5/ypx/gDwFUEx9R5XD
N1lxhw+NYogWs+GD30GRas8VzA5xSBzzwR73as5Tin51/zbTK+oSqc/NfLPKSZCM98DuJGaV+Vo3
w0GzNawJ68wgPu2ZszOT2JeAnh0GTtn955/Gs026zkn0wiHe4nGYOJqoI4BmXDG0oZvszqS0lfN6
i8tGhhwf9iXLBxqr/lyKDGXPg5uqJbJxeniDMapBgobeG4dULVAns5OWw0ItYNEBYg0S9qXi42pz
WPdjeQcIxsK/R6U1c3nn4lm0azQnLDLz8yV/mbNU00iiaB7I8VByQOut1cgF0cbVofyK91Evx3S6
gQSLbmCbfYR1npvs9kpToeLAShb9pgjc6LOXXcUkhw7yt9KcIx51gdcRRpYFQm7q5ZguAszyXHQT
7ervmZkUdsoeIJqBggdSDbIMwtFo0wWgd7OiezgnJ3a+6OkiTXo75CzhVD3W3vUvl7aVKc2+5Y2Z
WdtZ5V+zyCRQbxbSS6Gtvo9bvmwbItv6RrU8QlwBGDDwa48crcq3QsY5+ddMjTvBJCoHfCTT2eoQ
sKkIvfR++9nPLNs3/C9Yg1yM4AOCJPtF2FC2ty+brTHdjOVcFgMvqT2X3M8Tq8u+8XTPtg5PB/kn
KN1u49Jn24//JRVWKA76oAXt+uX9LmU2uRbYgnqsryh+sQjox/YgW6GbXiXaVhpsGLkfKXJ40C2H
TcFOmuM9NM59QjNoVCUtFqd7MW6Oi0kBX8xJK9O5eRhIojRYx6uKB/vPRUIXS57p9LI13IZh26oF
O6bLhfYCG2xwlYzRyB444N8z4yc51EdjmSqznkHlVVJk65udKAiVFTe7Mr099vKuUnNypZUqGXvt
67PSF49JxKPa1dTN0jmSx0V6qxcYck0tIVJSXIR1Ati8fGU6bbkz2gpfJe1hSUcAVtAjvWPutRR5
DK+Fl4EzxhkjzvyPYfDc8ZyZELDbSbhhrOz59Ha5ZqOyjEAXP0IrrF8gTfM08mmtyvg8evam25xz
Gt2ek//D5srdlFv7gP9q7NpBjGZue95lhOaCyLQWmkRk4Wk85Xxuod+zDO2Wi2UsORrbd3QdwMGL
kHKcMVfbIxh9hBcNU09YLR4UwB+XGGbxrZmsGqCpylSF1D6bqkJ8ak0j89lFp2zq4YIowdNajp/q
n1cxJddGaD4JGFsCStBbmB81QvZlGRJCSOZw56SdEhplBeWYEdeTB851RHHr1dHJj4b7o5Eb/GdF
2S11zJSqyaFH9kPhGWADrinZFggnotdB997m2GBguT/OMHUEGb2UwmD8aL1CLANeHI+9AVOlR0cR
gQWTjPk5wAliSGkP6+ZGSuTy6qfEGG/zMv0g0DmkkrB+3+3+1mbwwZ0uRnc/moNS1xtBCHYlsZBb
9raes11H0nZzQJMPZkfOtMMCeiiYgvzzcxGc0Hz1CSkPHfwmp+3wHmvxlQD51nqxphbBe5Bop+h+
hkUsFZhn2tbmtovPkOdnEFWE1KACTqJygEQ99Thuo4u45Wbs573ArtcXs3rEEzNd32OjJazdAJWR
Hf889YH/FhvtGrHTjRTJW4bKvDo0me3gRm0ogwdKibYyejrA+WqiaqwKpK89F8v+aNFJyX7d3GI+
oRDJNczQq9Jyu2CjMkvgL85IMHGGf1r1tNnXYFH0xr1xDMnbQDLye8IMJAmZp0UAC9+mwoTzowNr
t4uaUibAMfai3kGIwK62ij2a6nNAE7K5tn36C46Mb+B2QNzDlRIoOPzCGw2chzER9FHB9aIjVxpV
eN8BB822e719loahxHMgN71iDPk7meDz4a036JoFV4HXsJd2O0nXQA0Q/GksPRb2zYKVzYPZdLTT
YFEs1GvBbwosZ6P3r6yOW1DjlvmTMkYLlW8uorOnckpqNdKqQMvQaTbeuSC3D2xYA9LNvbBLiJVI
dOZ/Ky9VVmKsWpcewzuPqR59uCC2/44vudFm0C+4RkxO49bAb0eAZJn9+VhofSQQMYq/eDdwIExf
jSzYV8FIXiZQHLYpm9ykvleyHD/QaBVGg7J0bR5SYXlH2p7k0/h2xqNvdVNl1QzX8VYsD14QDTn+
8FY89soz/K3PiTMD3r5rIQxqJ4jeo7nU1TyrXxGafg4eWIODyH/J+9OlfiKV1p20Uw6vlF41enum
S0q6CcpMeHBSg5IBbgHmPny0k2DI2ehtAXvmwYuRYneTLxtebYGn/yKL+06ZFEFqZpjFnrhgJ7I3
Bui4NqEKgIInXznIba1HdGKdEFjc3EWrKXW/zjFfOBO5SGLc8uCwmfwKUK5XT1tLNA1+iTHPY3jR
P8beIvh/XJbJ/9h5Xn2Quv6iMPZW5hOig5Ytn2U+TfLvUpFj+smfZJ7FSSfM+E1b98Fb8LuI2qjj
HwPHH0lL3jS9vsnz1K7Bbe930H5Xcdu2WEp3hIgxSuafx46HrZhCDYkQm+8hDeGCBJ9F40QXV+Fh
qd8ep0G9XObpP++c5IAb77VktSgvJiLWBA7g1fEXobYWGzBN3jE4VcbpJSNDUjxDujmgY2NyYjuU
HRAo9caYwX4sFqzDb4YxAUdcYf7zsSW3lZxjRSBh3/C0ZcEZEtjxkb2TGZa9nQ48v4A5NszM9ZeT
qobxuRV4+njazfUZSUBerT264k8/2t6JkvrwA5CrbYsVZlct32Mzp4rl562GRY/snNCi8kvJfW44
FMPioccg/nzh25CeYi6+YGexMtMbcMnbVLEDpZAXwU8shSUBdlcoG/cFZO2bzxGWNYoFJ36YeMLA
v7K0gHVncYij/EKu9HKYknrnrf06klsvVTquogUATfYGxgJjS9WzwfFofeyidu4IGGWht7TLI3vb
JBdKQ8iYG3uCM993/S/A3LbTQl8hirpO304zMY1q1zUkllmvm8M67AMScbxo0zDIcKXoLOOkvsO5
DtnbUiweoQyov/XTRPkjv5ZJUN5zjAb6Ocxqx5bsvfgTNzHyRgVLYMk51nnEc9HQWosZA+GSdQ2W
CILZQE0wtQG8d8HBAjMzsyphd+/SqoqRjpHHkFvAWXQPjij6IyB7ZFO3P/w/+C/yGwu9iZ624l9E
Ehx5a17Jj1t9+I8QCQMey5Z1dF8/nndJC80GgrM884vNa/AxcoR5uAjROsQjA4xq1wLRIVPj5M1+
JgNZE5DRmT3ofMKAFJSyT+83KsqOYaRxfLE/m0qoFhGxMIiy1lKZPOyq7b6qgVzJJXPGdo0FU0I/
0zeMm9XK5Uy7XAvuuLY2zC192NE8RCpk99MaghGugow8H8Lhmq491KBtOaMDlv6S8GGN8s7R6WEq
UHEwjZ4m/+BoZ6ns46tDxg7B4iRLF2TPCZ2lldEiKQcdfeW21CUuCUCkR5RvloZPRdzA4qktRVUa
xdiyEJyB6bBNG0mIddAw2QiqePG0Kaw4UcjRRsksBYL5A8ZiAm4O/59sL6er1GNvTJLXBhOWKm5Q
RGGacORynXzk2DJakm47JiPIXan3CMVEOLxIESqhf525cYSmT/MmOcFxCFYt5EVvEDH/uutYHbEX
QE5F0aTc262/+c0xXw7en0vLbJ5EVCQ00J4+fyYX4DAfshzcLTnT4KklgTRZuUdzI7sSV44FJMVg
I3yMSJVYkDwnAwpGMjxXtQxPUZyvJj1XLYQgkGMCPGbW03qNeKhAderbbnI1OCRqAoRYCG9nS4J+
iTVNfsNVJBXIKM4dmJkdnp5iEm1jCJEFXqCFrF9r4p7iORNOX9TXz4UiOM/+MQwX+uczLAZydkxg
ZkwfAzwpFZ9zxlQHpbU/KDbx20mqzb47Hq5jXtwGoZNT7xffXLWL/G927gTFzoerPQjC80J4nxNQ
k93Jn3lTNY6iiH4VPVz4DPEhEYa3XREq8D8pAPr400L8jh5TajugfmlFaStWmMiVYF9b067Tt2w3
npkZ8YTTsTqfrK1gTYx5ALb2jVaq1NclwUNswx25K1gbp2+ZUPbeGeNw8XKwqf+ak5lKPP9LBKbZ
eIYh8Ttle7SJCdTghrZyVo3Qt5mnhNawB2IgrjTGjT/EtRvv+1hvgZVRuw1mzRBtyj+j10cDin1j
uKT9TQXeoA14ZikwWWe7b/4pt1uvsWoFTsCDQZjMGs5YYaEpyJ6qzdFgbVBTrIBSw0bFLKFgyvuG
4pLaHw2K73DK11RN/wRTUd/e7YJOHy3LVlUAoirHtDruUgVi17v1IFge9D4WLytSzliWC2GjqoC5
xg+lFn0RRGykaPIrGHBg3UR+Nr+cLx4AxInxunMyaEFpT33apyVP/q/Bh6RhXTuUNt6uEkztu30H
9yC4NwfNSWGCz+Tmjzphub/rss3QTZYxvy7+Yr3fmCnRrkC7CFS0fzZSH3uh75hdHnwthr+VY8r3
+QfAvydXSSYPdtUnpunvHDDbpWK7maoBxFO4I1CAvpV3ezSdB8tlYISkFpXWkNYmW60tpc5ipv81
Tjt7DFXC5CSwkAiXF2blDgD0Z6Qgik5RwSNLgA5KghsjuDAOx1IbSOhsOYmrubXhC/ZwaJvgF0yZ
WgaY743cY1cWU8Qcog96m/h+MhcJb4rkntdzrRjEVmH6OgYTKkP7509wDmV/vVz1681gB6LSa0yb
hsQBuDqOBdopqwdE0g2e997djXlMXhdWbEgKBqwpnR+dIYaMNiRVGG0s+BLmV7QtuPYghnNSaIwI
u+LGbEXnR713LoZExnmAc+UYi20K5+2jrXdLJE7TXvMDOlrWgjs4Owrj5GqiDWHl3Ko6bBUXgc7q
i9xkIUz6RDmUGMfPGc++xU/GqEnPOnxHWL55C6EfFf7ZnqVzR4gSBXk1Da9rqZR/SjyetqZF4SgS
YNH4Iuu6sK20LUT0nk/TY2fXG+O3pQ7H2POtWnXQRr11irVFZEpFp+/XxsO3HRIRwh/PfL1sxtg/
Vw95zXLLL52++xZfzsHxVKO1wDCt/DaYUBElWEClohpU9CMO5SsBqCdtqk0sVaPeKvVJNngJD/qy
MkP3w1Biyz8CP1xEICB6jWtpEK6GLi78n14H+w6VhXFWde2aj9vDjSAlUYT+lAxPaBckpNkLWBCr
iTSqldm3jgIY5MjGDTSZeJ6C5FfoyfLQbQMM79W8EiECXzCKs+nhA+vTbbQx4CpG+7BYCwOB5ksL
NWvu2yOd5UMWFlMeggV3KIOfi6urhHgQGJuvoekHoB8SIi3OZMYJLP38qICxN86IoQlBU36uRqgl
77fOm5DCOUwOOQ/82f7djbNezp5lTX8HcfWipvJnBsGzA5orYqW15P6TFEm6gk4WRH4oLh3F5QF5
0Z5kdlZAjdEwQvdHHJYb2VPuqg5+Ad8Q39P1lmevdOahi3wP9XdZGuPSgfGrgE9hShhKSxC2rsyu
GMkSJcYHWCnobZmXwSpBSFmXaqU9lQ05ZLgCFSdUUjM8tcTe7vAqX/9xfQ3+a4zQ14z2riGMK0Wa
C5gwGwn4cluDL4iXGoei2RPl605sqYOKpVdzFTlFht7qJkommhS7JErGOvDzorcoI2RDoqmgWjvr
caunPuTiEUnrE9sxguhJu+j1RtUv78R/lzRzFJhMfonyjqW/YUUBLbzeWgbpdRmTR5nZQ22ZG9vF
1FCnoQVajCZvLpt5FPR87E5auUluL3sCNYJ5qW1j21UOcs2wcGrIq5NBfIPfBqvI+u+JZ4OUJTe7
oQIJoYSQBxTJZ5MROvW++pBVLVliOo31MvgRDzBF7bKjt5r7jsGKxdorw/TpxIQIAVABnqJ4mu0L
vtr5x1Hc4l0jOlNtL6Ihgu8EIFHB41e42MoG7l7sqWVnvhSsxeSOJ9cGj/swPQqLnSl+YeV5sHKU
basjsJowzRY3yuWRPrjxVZNxve2PgMm3QMnhldpU5+/+KohM1UDog6nAIk61+yy/QWm0eqpoYFpi
1A6U9e1GxHXPjIT12tw2J5LcmOILCNRr/7i/Xkyi94u7bWovRS4lCAbElPj5B4zaY2JgE2iSj06v
YHe6mbq6bcNpyz4gK7HIFmh9cZt/7mTONBirXQcLDN6DbAYSo8OJWm320V2J0EBXlqqUJADU4n0u
uFVLWOXGdQj5CY0chdse4dSN6S8ZLyDB3WhbxEKb4W9qq2u/dRqcOyFlge+Fmx8tcBrt8cBOIGcC
iEF/yujKXUjV4Oyszvy7Pm8Huw72hVm5RYt9BXOrawzGSkFkdW2Qpzyc07X4ttvlnriAHS+Q9Irb
uaOh7dwkdazAwiwd40qT3G5P28zZBr1ScdffV4/DnipN9dA3gv4LX6K/DSqHXVRgozu9p961ok+e
ka1sTs/MUWqYkIZWSSlMphjPBS7Ofaz0PLdMFxEF60x7JBv8A/x6Sw6+1ya2sgIhDdYTnDUBF2j6
qFNVLnbfbrrkdh5mYcMGg4trc4Hg0G7QBwEIKFIE961PVpH4k8lF6s9FYZP13reAvH3x0fMdoKcV
XB4oLa2uinaanUBotjJnHU5W+BB8cTJA5rPWIJ2n5/ci/SFfzcono6fvqf9VgL8iRksmg5MYP704
iRsehuot4R99XFwGNXPnCFsY+yddrOJ4bDZMZko2QCMKgjBO3E2YGZ2yei3oq2rdPCauLL7v97ZL
OfmIEMbukZXpWu9QPF9pAnatiyI0QB1sLVWCwrUWbNR61rh2SXq7lxbqPtrk0SNdAXNMy7WAVZMs
UmJwItVMdominyoMAeTHswKQZPsw/wNpO/fVTkp5b7ur566uwKJ7t+Ku9oxASSmlbhVXMZF5xJyT
2ocwndkNly4kqcXITBcmmommHTuzezfUpDXbnRIZfToPWjFJfYHCHWQXBOb9yCWXkAEW8ANv7lPp
YXr/8yaCri5ERFXcoaoPRVlg9SPu+tw2JjX+gk+kFXRYYaNAQOV5n6eKwnjKu/wN/YAwr5bLZdRL
gYxXZVg/XK6OyztC20jrAIw2D3S5f9IHL9/q2M9JQnvplkEWsMcqqWfMCbgeBTLYnV8iWuP1qhr5
t1EZRblUQTGGZQe1iGWuLnIlV/Hca71MkcRGM20ZlCI3WQtNtoEy5uuaN6Y9M9hYr56eqIJWwQHa
8EghAjjyiCU909NxsD4wzhdssxvF96uzjUukw3gwJ3SJv+S7H2FSV7wsSYbTTfXhNIQxWIivaVs7
poKaj747DK0tba5rnsTORsBptoLeTw+WZbPq9nYAPPG5GAPBXuWC518PcLCo2nGcxBNOSAZIJ0DD
W95RMMaCDnTOk6qFQtpoc6cwGXJb5ABpyMJUVrxu7rs4BrsL4mQ1Up2JDLvhjJqGXYVpULAsMrot
N2LnOaz5NAB50LrV4FzV6zMuUoGqV2oT6zdDNBtWzw2ovh7wM40aF4+kfu9xG9mdYJM3QiYL+iGL
S+/1iryvLqGauKBph1fGwqAz8XItmWOXEG03oZdrAYoXrH7NfYCB90+eC3kdRq8+OVleD5SZl71X
Wn2cjOpyEw4GtReo9s/aKGrbEOOviM2sp/aGkOfut5S6i9/ZWyDyKfDAxGl8uaJOOeRKcScM6Flr
kjLe/RNhlMIJPByjw7iO/hDs5kjaREFM/4FupHY+UvnPiiIVyo+HicD8qzT1UpN+ekG0sQbCqVDf
nKZdXM6t9iEZhdPwnotbfvNpGwPLZf6AFAvff00woZSw8ryIXZ56PEWg8PVQCU7u27Kv4t9bnKua
KuVK5k25MrfZ4g51q0GRV9/aZfty5pjkQGck3D3L4vfY7sx/3+yJPk0iA4x/M8cU27+jcylRbPh4
GzULZINN8QSHOuI2NNvXzpKQVh6JeuNCtJLjix0BapmSKpP3ChK96AeFYuzgiORtrEQ5gIuJGC49
BVN3seET+2W0Z6l8z39pSu2MbzOS+69ZJEsMJu8+Zsx52WCjPWVVe4xDhNFYXvFaA6NqEZV2olDj
VLHfhRi95j64SKDBWICqtfqoeTHzqfysQnH4BEfz2ZK7CbEusDqCrGZVcOVS620+InUXhYLUiCiC
OcJ6Gy6Jc7i1bQmtm+aEWTFIzFoaQ1uSmohIFusVGpFh3LtP8wA6QqBdWs1HMW3loUh1TmzAXaS0
OCfdpscGG4uyyUXK4eGfz2XpWRMUB+5gOZl1z9Tc/6KG6VUvpptP6v2R+iJyqlPx8wYjGN57udEy
EbWpXqSokhQW2B2rRGwedsKPTp/G68fj42DR4L1cE8Cdbz5EjtKbRiTncqIS3f57qcf81N/GtJon
Cjyy9JQXJcXhjbg+mV8oAuyzKy4wdm2rjHCGiNVvdr0imzhlQk58nFtXWyu12X4ThN5fsjXqGzqY
nMxeAPX95vHT7FT7g7FV9WwjNklJBgaYHTR9vn8V67eIhc/uXqirDZdls61CAp9eh5JJ3LI/UNlX
BjBKzLzY4v7XAMcvrKAftDoYVCMYtpgUgNAIX+qRDbDMr+z7C9QOnvtR3Ml0TnV2PZyau6C4FXdf
lwpeeH+ZUod6Z7gi71kEvIeLG4QXiWlvfxPcEd45V2qGtEnNbSfb903EnAis4/1paU4TL5YkvZL3
LVB+qZUxPQSXZzE+xJcAbRYXWzJoxHd0GbxwsOvpq3VrBd9WPjx1Y1ul7wKOZvD1dIFhmmTmEgAe
7echsu52Ouii8Wa+zpukRQLUOJtVBXYjURPoBQlgvM/hyqv5+HZhD9i7MIkxSLoI+bc3B0hXnrDB
ipxiIagGEEyELh8NwreL2DrAtxAxTXyeEtFH77E8IvERR0nyJS3w9o14/maUy4x2eJXy1klREXke
z1mnezoAxi3oR2/X2Sij6DqsXWYuOqlqfP/0vautys+m6fy9I9MblPjyevtBgjkp5K7frJ982Gg6
CPsDEK9p78il9N7C6ipCp1b9+MsieiUXogcWqRYq7QPK9td5kCM5Lvf7W5FPWDeLqiVjpdtbxYXj
42BSpiOHpKvizOkUwB6tdX+QUMPyyJOTftfYl0wGwBD1Sb62iRY9TvX2HR/HNR6/4/urQhgbFkXv
xLcpPpcGfD7N4k4EcE0otpD4sWxIRtBvCpBguSmL3ylG762dZqpVEdV8Jxw/xAtQFp3XPhS7DD1e
S1HhwyK2t5dW/SB81b/RTwfWYwskCxqqsajHFm1hvJYQVUJVWBdPcbhbEx/KlftVRgMq6WO9rFno
ppv78Oek0f1u8Nc7dOCxYQVUUOOxlDsBPLMvLWidakPsDjSIzyo4fAgHco7Th5/aDGU7bbE0rGJh
I7hxGT7UbWuZumNY9SqGpuNEKTVh869Su18kh6d0a+nluEc0mPNNnXAOVBqUPq6ShR74joXMlewS
K//oPVyDGK6TXyPwB3UBdfC+4+38TZlMyDn7lDdBb57j4yEs/qAJ3VdYG8ymJISb1dgQiZxMLjJ+
4yOeIhu3fVI8U/ef1LU99JmQOIBPJnsgvsA/hBYGZj4fDNzVwy/t7OLySLUeXXDiRjxTYxSps18R
+iBHB0rWsYNfhiwEB4i95XuTu+4SzvFdZmm97/E50YXVUUbHHYn5jPdutK9hzF0GwSmqbRCanE4x
Mn1tep5D85Pop92/Vy1WxjMV+79pFxlny3/nSCFWoNQU7AMDQG6JN+YC3looNuhjylTnqWQaSmyg
OXrkb1buQGpSAG9GtlRVifNMT+5Bi50zMsxHy9ZV1Ok85ldCZeA9ltOwWY8rqlYKVrEcY9inrhHh
x6pKq1EF6lrLbE+rM5xM1YPF61rhN5zx7AULCBAHyTayzA4QhZST+9gWnFym7bb5MQe/HHWIRomG
UEOCMQff/xoQdyNqzK4uF2n3M9ETqx4mRCRBI4AzZl4pNyJ5ohocJPRsoJAgPUDnXtWDApKl7YXv
RF0Js9lDje+jQmQqO9iaLnXSffrKB4x3WLsti6yQ4Qt/RbkmfC0J+5WuBUgiBXD2FrSu01Vvw3mB
HTWPgy6VVcqDa9qQ63t6X4DypCT2b72hB7A1wNH55AztneWLSunRnizkWybYUBDGL4wRh2ux7OxO
Lh0pxVyq9MkH8sMfjQzmLwPhdlyLi1cIYn+MCMHWaKOODvmZ77/jXjlr2sKMvDNBLFhGJxCCHJul
6z5S45daF+kEjv98QkRG8Qpmr1uGV6tsSpsSmVt8Nu0zk3CD90npIINKUBt1XE2d69v/PhkhPPsc
lLxzW9cbV1z60Q0dqjpcZmhnVXq1cGeWu2IdYBVs2P3KmsOgortr5Dxur3jKMVxhm18gBriswqkR
049hlXAyfF0UxqH8ic+pwEC9g9LMldO21X/IZA8BIBZKmQwXj2rCc/tqiTgmsgMyan5f/fOu3WbU
Ly7Ilm3KPZzKRit4CKICAJkuIQHNAb3xSvJ7QuO+8bnpXVS1QD+7mUAMcRpsqibRtRjwzDUpcrCJ
Mh03LRhwsSWKrFR/cAIAqKtnLN+bJwjENZeYfpUrQRQvghXcmrApxM9GalnR9nREc2l5p6F9vYKu
h0YgaJTH2OUZt6CSPLITroinR4e+qSvClvL1QRFyGHdOs5mVCJVkvMV2RiysKaauo9TU48cs0cwd
5s7UMMFYgkCnb3csbcMCsNhUHq/z6z+qi2MES4nXXMpYaFRp8QBSekgFXS+GzF7zqr738oKQ3NJw
A1ziaYvZF9lZdVO69xfjZ70W71E3FoD/j6RozVjlMdWdS/+5pyeeP7XPRwyQWm4VB32Wz14WdT+l
CF0CuXxxYmr072c22YGWn41LSSg33IgOtTON2uwazLBpLjmdRp0hHHO93TFw6W8gAm3839vPzK6D
1rqUnMgb/Yi80SpsJ/cpUloB6pnD8FeUtZIf7vRDsH8ANVdb0l9YzMpVsrpJsDg7h+AfMIoJeqFi
p3MkzVwEJrNFC51pt5Nvf2hn89IyB5G7Dt40S6fDeYHEf42WVGznwJuNVFQjnf39yiLmFfO7nUj4
2h1aloX68bVX+MT9xyDoxTxPppFKjLf6kP2w42sg25LyrEW9nOFwY5uiZSBWNgtWBviAgi0bQ6Kq
6SD2yLNrK1OsfMK0MU9SF2KOJGYSrzIMkEAi3Ca+mRcbsEIVayP/zXZdga3gobrlwt0xULHjGZlB
gQANPBT+2RG7A3Tv5zfUYpNVCO+65ivKKVjo+1sngEcHearDalNMGOWoUt2wu9f55ZaTNrymDPyS
rOuInx13jtmPhxmg3Ht3DgeY109GG7aGxe7NmUzab28WNKhILYDiP3BpR4/xE0sB0yH/ppKTIKuK
YYMBKTXQz9KkJZh5lZdVpayErC+VFlIQ8/MLUll1coSnwtLZYKilHP/2xvc/XwLnL3jGYS1doC63
2FSMxzmg/zeJso2XSgs8Bo/zCWxqw5rObZpmBenyxHj/ODh4s0AI8bGB7TmW/5oSZVzfckOrP4WN
jXLwAV4id4J0I6KpdOEmUscZ5DMZR0BHY1cUOfjeF338BYbw6rV/WyN13WfdMbd9cl31OXQV96LH
654BjWEhRwUcD5K9U8kwlrb7gE3zR4k4pY2NHYwqSyy3eOK6G1oJoxcQdpVJITHVGDQ641S8JPP2
/bNartHtPrrT9cSSTSUj+74dZAbRv5qq5NYMju5TYgWJnE3nJA3PEiRxnR0K2lIeqhIQGK8RLsXT
VSLDXBHIuFWO9Jvg5MR+kPEYqzRQIwep44ngE9Q5jSpa7rMt+DWXhH8aN4/OdNzwEZQZxtZXQCKj
p46RcHV73yNKcUnMFmr2OrHkGdbbTRfCUnU55fARciJv8bZHlMx+wyo73lDSn5i0QwLg1Szq3fS6
VQHyRr0Mku+jG+9GHpLIxKpEnz2NR7gpVBNwp2byvdddvRU/jcNuwRwOokb+4szFP/T9T61O5ktn
5hhs0vXrVPUXmXMJKhIj6VzrED1u7xlY1kp/tJy2auy9G2oxUahx2c+7NSVRw21KDzJ2zk0+l53z
JxYfqDsxyOMmq2a79eRkIUAjOiiT6v/dEUUeklaxg9ugD9BKVS/jpYK/ZrP7bX7OQjHiw9U0DM9y
dbKC2DRbtVP3TFxURx7t3b4tOljw6gOwloIzft9j8xb2sNnJsC+Xwi/7NdYUuA+uAf/nWIbVD2Ly
GXh1PUrgxnmYFgAKTw+4PF1IEPQ0CZRGwPDgYO0dzadskLC5EWjodELCGUhBCA5UD58pEzk75SjM
A5uujVOPUlZ63pNb5cuRm08HHb2LClKz63PKQxINaX62rImdw4Ajsgdhk3qY9hiI9SziWELcfxnv
Pda/zaKOiyGTtMuNerZBpHsO90gaZTz0m2sR6qcgtYQqe6yMDC9cxLHBqU2aeB91yKfjCgBWS2v5
xg0LKXuW6x0BdeF1H9RzcL0nl773RmFtr4gAklxJNGjO5XYXSZnwMvFu5KxjsduApENKnBB1kSvW
YAsm5KXo4JCYE4grKbqHSK0yTPwON6M7YeC+MEKePdhlNNi0+6IzcqNVtHF+9haB44iBtW7fEl7U
E+M6BOhoSKsmY7Ac7EfkPiQeExOLFLiMKqNhPuTvXukUeiq+Jo4jXdI6NKi8j8HIqfUP6sy8S3gG
MJZaXoKwz0TUkPEg4yHxvusjGWlzWBY7g/svJi5QOTgWIJbFbAFvH7t/77yuB2/I/NhVGZ0szOVx
zat4wAsxZ0T2EAdhAu+rQiw2MxLnFSirGNg7YLAkdh40HhGfWt/YN9KzkZufbJXnBdC1pK4lDt3Z
xVzA9U+A7oen66PY4Wac4OM/dntKCRtGCa5IbVnpPFZxZptgL8aHqjEAsLvyLHnFgEPBiCKNnFqo
ZzBdnpimipSL9Rq6cxCxLa8MVQRtaqiskD/mCD4ScsbsaZYReC1pCs3MMXRqFDk6tlDCHcP6jUm6
YBfIT5OjZij7toDocXk7j3NzRuWAhRgLTUtx2tw8Y/UP0ctKzYt0ZSERGjDzKDP+l6UFuO8mdno+
nV8FwZCX+VplIuP3L5pVH10hHJhZHCOFB3x7xjXfW7RnYSuibYiMBjg1CdCnTDoULtdoijoqI5if
FPYcpi5woRDTrVUiYJn7Dzb+TsV8+wv2gVOtQRXhqTj4mUUJEXXw8a1FVD+jKLPQ7cv0U477Xyvh
Q4qwnocHUU0in+mUBTOBLtlwbLJ2t89yXCOvmnz870PfpjPhz0QtSiTatzoUYDI3xh9vuqvYuRV/
f7P0liIRBzPgMgaUVqeNhtB62SXXfrzviYJzvEzCjVNFckjMicQoBsrjUAY/7AhpXWVSmLRnMTx7
evqeDR5Do2AZRXuVZZhnLgEUU+5WCMD2x+XxIFMsySS9z05fMNinGIMXmkjAAgrik8GiwVXr2Ozt
c0e2NRR3kS/cZmndXG+4HuNYW1RAHeLCMu8yZbXtk62w9DW6aB5pDdY5ArtQAQ2zhgDCY0atUFh0
ARyuTypC97rz2R2IoSrVpwuferQjq/bkXQ+BGcb1+sAVx9r5U1d8SEcoGpZLVlMN/s28IJikPbQO
ZisKX/oabZYPffY+wKmOnUekE44k0uNY0msPUwZjZiQRMdXgm0Putm5vtXlDpCGECJMI07GnAT2j
fCj0tEeTIEhGj/v+8qmZScIZ7dcuGT5OKTcDtXNRFUF4+x+sDRyE5AGg4fYDuv9shgDoaa9ig2RW
O4Iu9tXoTzNvRS/+mXgu0nz6y4AP0iHgJkPNIfqvwbgIcr4ZBLqMeYeLJh6ARq4pxOgbSuKkMAx5
/YkRTodQUql2FP2fIX2wVrUGXoBgnIkOL/nEU5jJzLAadLMLJCbIX2b+NccjYNeIXM3926YYPrk5
6HnIDrqeD1oySUZcgjUg6J0fFShIXpv83n01jwgTpVjTGJcWLgcI2JJKogVHJu3mlOue5Et+Ziel
i51ElGc0PAWys2RycR6GbmxzPTQ1Z7kvDAf/bsiNAab5Ew5PUfF2jUEGYFYFBWs+mlM8F7CBioJj
PFScAyDrqYYXSQ9LhmNVk9/x6wNU0bVxEGjc4kEyKEm8dY1IDFaxP8iaUj14zlGX5v/SGC5Hk2tE
mTa9pROWz7fiLK9d1XDDgn++IqT9ou5cwkGP2IAX0WLMIY2Ho3W50a9rfCyB7KIQcz/7x1SI4yJo
kvjf/kWeBjqyG8IHN6Phf4gGntrTzBNeM9lHP+1BssJEZ4sQNXd6EfltGHugeXpescGXjDCIqXE7
PP0TqIhThkbYdlORgl/F9gf7FkUFUOEL4k/+Y62QdfwckVQNw56kXFOaXbEJkMpH6WId8rOa+dky
FbfiKs9UYJVAX702ZG5HPVyyzekIy0dYF5iYBmFqSLoamjctLcfvtiU02cbWA41IEfBaPUA9ggv5
KwfGLyDzY48xTFENONAy2DFKy5AXHKsRVhjXeCp9VETKhSArI/dFvZXjIdde6GDQi2q+/YJ+HGIN
ITu6QZwodcUXI+RVI9lWWLwA6CfyRSUY4yvT1r6ed0nQ1AYw7phl7fxOlbwR3UEjgXFY7UmPip5z
Hmc4YjzroYkAU87wNYL85OVxiYLBdd2JH42QXNOuFZPtlM1XR7OAbaVIbQxlNsRTI4zWgusjVESM
GqW6xCOuQbnQRD0BDWqr2/Uf5qPvkDKCVARDlCyQMcYkDFYv+svmG5IivGrGdwOXbLBa94UE9MEF
mbVPufFQ4dx5GjOjFEPfO4SMTJPfyajPtrae3Sqb9qBZMFNLDsPm4JrZs0n2cp7Iz0vrheaZhSHh
/7lMUbEnsxkoaKJXUOnSxEMfUnLDZ1kVBYKW+ct6p05ep3QDYnv8NlKCSw+l1ukix0tYx15TQ0ok
0dR1HMlpAGQ6XgDBu3EzVT/k7y27u6CWivfhD9Mc8BEWJB6BxAH5eMcE6HxDflRTTCQC4MtqSLcH
N4fwUJH3F3QwTApDE4PKjNwlwY0zsaYCeYhk4wC4vE1g4C8AMwvSYPFhhgBJGcsiWJ3RV4yB6SVw
w9OaHPy2vJOF9Y8UEoPFd2bgmSkG9flIVNIPTzQEKn4mK+FY2Uin6+QWWgSr5PhtQcyJ4gsl5inZ
mWS4TG6UvMlskXpyE/UKc66duPaucdYXozbt5nNkvXyauDicg8G4LNkCLgiZFsgEdo9AsCpjqpQu
6IAtRnoEfg8f24wz/+V/kGDag0h3fQpHRKyz8pssKqx0FDYA5eHXi4TDAxYCFGyRy+TkLw0Prmc1
P/a2Bga5uu1hhzEpzWtd4Q1+8EXla8ky0BIWRHkglj6Tv9kO2UsxeKhOnFv+7TnAIqLI3MJydw0d
oMmTCG2aAS/kTnIZFGvSJ4VlOc/dPzB3IaLDd4PQ6NJk9q07U6XVB9JSUe20yGyAmChBwkaO5vM1
m88nLilj9Jvb17f1p1Q5bTHat1h9Wy94qJLnK5YN9xL3i6++jZH/+3z7s9hXlbpHdlWUV+0G1aZY
CaPGEFkhW7fXRxrktm4/bAkHDzr1vh+OXEVUwbzK0WrHlYdFjNh6OWiya+dIZKG7rrxdmShz7ukh
wcFcKPx/+8It1J8fCQI15LBwX8jLHAR3K5FviGzFTJR7Heyd3mTsiFXe0jekI/ndDfiscOefE1mb
iJ+9BU7ZxbWzg7BlAWkAgTyu2FFkEFh7XkNAxXWas+kN2PF4OrfB7Q+wrdx5UPQOG3t5soEf9xmb
7MOdezRzPV9K2AeJIYd+s3Ko1jsiCl02nrwiSyjGZI73zcXjU+DMGEgjrAEqcKv76CsJnYm5DJ3B
I7wDyhQHuvp+Nf+vMA27Tt3Be89h5mVXpoPvWbMd2MNjC3gZsInDjcRjQasMeR2CWa1rRwyJxlA6
ifgUubNwhQ+5WAlQT8DthcWqRifsoP6NNcbl7FENV8R3me0vcbrCtV2BJStuQLfoIJiJ6bRFkJWk
IJNyet/2sir6Eo/V0ZhyOe2SSk+Q1AKVe5d8Q8mM9ukIwLBf9FnZBqKISjAd3WLB+2YRaZWNFQL0
HDbGXIOgJa4ElOLfYJ4hhDC2SXTA4SbmlD2HVOCCKGP7RTgGPnCpylBOXRJ+G06bZ5veayO75ith
RIosivy9uRIMHFSINbr3JVU9M4afPuph3zqHKQAn+m+kHggEF1T4nFp2nL+CK6JQU0tfOXpqYsg7
FQdqf01Zuq6O3kUB8aErG5drGNMXWXeMoopgCIkotOG85HboQu9QeYNwXIEFbRloMmB5Pe1CAN+A
RM/9sU54sS6PMBAP6OKsbwdTiGGUXVXF6Um3wPM0KKJe6DMeVXuc4NIcFbPGV7p0afcXYtvhYC/4
NGv695eUehmn7XBCHAi+Wmzxx8yDS66aNVZvQN2G3PWc9GEO8sb3MERMJ1fsEUoJWsAlwjNCBby+
8Ip2b4KWFLzEv1hxhxzMKy0hK4fi7zJORxwgqq0PWKOPW/y7gQ18ssA2N8uuWdFfSCzSLNRfQxNQ
pQ3DXJSuJBzrSP9VIy0weQGcFMuwIvz9Aopfxa6Lgl8AldGxfuc16hsFExHEVqbRO6tDazXksV+Q
zbj3OB4orYMVQgh1ReO0zL7Gg6Kid9u3UJGMZYBxzOLfqvpHhMQllj5MGIkc97NIWlGG9AHhfDfn
v6vbIG1Vrah+xdEE7TSJxGFy3pglK3Fj67fMPXS40yH1VUGqJcIxtYoZCY5xqp2oIxH2f/4dVPmN
mErwn1HvnpYDCLGk4mBQRSMXm+NSE8DEExETYMmmJrYMrF+P//2MYnEro2ZsuTVBRcTAUS7oU3Ba
4LB30BjpKCbdN7bcUe+JIIbNZK2H0pp8hs+fODeAWxkbKG0DcGxlOTntzvTBctVy306LZqfYgsot
wXA9GP5OTIa1n/EPkPRf7Oeh4z6uHIeDQskzdTsVl1hAuPgBXJc22hK6lPElKBSwlhhFmIv56hLM
r3IfQguuKYERAncFmJQhhzfZklIjQ2S69ZpIrGsylQYnnP7gqHR1bM9YD4+1/YbSwsvY9PUbmrU3
Ec9xfJQ5KCKj6RYOHLlqOxCcCLTG0pBBVaLZaZIROomz1cXvOF5QjJ0SJaXi+1Mt9LQLSCE9SMO4
oj7Ja3H8T0HIgqhPKLB5bRfkhaXGHEbrdv9noX8IFhN4sP0XQkEdiTjeiWVivlLgsEi9v4Cb3Xz8
KVEDp3ObQA3E3BszramYjvXnhnuoKWwAkmsOSv2FTWLpoTpd47cEM5AS5D9bC1Of2mIhoCu5TKNd
Cr9tjuTL0jGKnxP0vVlIOa3jPAfJEH2dJiRrNfdD36edJC5R+2ZN18JcJJdYXP0iMdDvYlD2xTu1
2P8vGLn/EbdB5C4D7Q9chf2uILCIrRsY3P1xdUAfxrqr9j7diTnLGvOJ1flPomBBPaZkgmwiV09c
fQuU+0vVMKCGJdf2gQxL7nAjel8/nu8A/Ri+W4NlAXBNJXsvE4Fj+WVJYxVqYa8xMShht+dYoAEr
wtnZPpNHQzYTmvjjSXUIEzd8S/2iQoAAoZvfqZthgR0DoxXZlRFtedzA0stEuqoIUzgq1S6OiMLv
0qxW/7XsmTLZA12/DpD0PtKw6mIBJI8CX6cF7KgO6rNwnwAgNQHHllaGQHAr9x8nb4jvy+h+GkA2
PAWBHB7LGpfPiXm4S2araacLAJ103GSJK4XtjwV3jaerWCBrb+4R+Eglr+RVqfg/qLV9/XyZRvrZ
re3YggEp5lOeNJPCNgvEhsmZsZpp+SzD2FI3QTrj76wIEZ2ODP4WhQms6NkN52gafxaJmH797eDi
bWlHKoWEOohEYtzpZWIeDFb+eZsQyxLal7uP10yyk18P0hfmA111Jv6CNzAJsWw/WT0FvwSrPGJ5
56dUL9AOP1R+1R9otiuR4iD29WvFsG/kqhp1EchdjkdjldcWpvylxWa6HB3y7e7VjXrsC2k3ry1l
vEXIKYpd7JinO5M3jou1rrb21gEDmOfRlCfGF9lqKLBWfTKBXlIuTHOPiFRMsPzv4oSznXHO+H+x
YnuUCpw/KDoAthTFkowLEPR0BPpi8wvwfq0A+u6BYlz3XBSBGlxN69RTce1BuuKFGxMFLj/nM9Fz
JkSkWVtvhu2/LW60fO0ENNiBpkk8XUnXcrfgMvhDevPtcBVgDqXkkWmVAhP+CAPUiiuW5zl1RWPw
NoUUJZXSZm91XyV/o+KWTzLApCyRWxWTsCCZjzGgoJGdMSJ9QHl1LXypXb5Yx2RtL6iaAIV+9les
iDEFjy6Ih7RxDYFnpMqKCwamp+VfW9UL9jrSBxZ6b56fkLUb4ljZcy+++BcO9PGNm+1M8+aJhWjL
e64Hc7LFfW2vQ4aDTxjTxZlUsal80i6fD+RmhsXfKrp22PT2edrqGJeG7xLiK+Y7ztL69q+AWCGB
m/SUfzpXse0hJSxhxEU9NLwtKK6sGjpcQNy/2/6mM62O2KfMwCTiSafdSmrGctMBxV5VP++HHQ6O
t5IBUZmEEemxwoLquRmvkiGlU8xe+D+gz6M2TrF/cSRTf0g/mv70AinWanXkoprQ21NzB01auiYJ
YCAvCUT8fJgZzmjSmlrN2zjWwvudUZG2NZtFPLCAYIdZzKwPfjsx98BPv7rJHIvIqL3uj4sFDLFa
fNIVY/eDgy7F1ONm2whsPikc/MG1A8KwfbO7eGW/fTJunMY7rNu7jcfKxNoE/kQirkmw74v7Sax6
mKwfH8nUsUN9EUi2pJ8bu31N9sjYIE9D2TLJLXtvkGDegzj7zausmP/HEOBqQj8TFHTXMAwUHpkg
C3XM+K+7ihk/AJQv7gaoNx1NS6lHob1MTcJuST5vfB7SUN0qSSDFnwezoySyHniyDnAkHc03oO87
pvPqn1A5HVsHyeHeKVmHleyLoTfPOFe3MjoA9KZLdOh8FYm6H+b64vJ2HGCwPs6bUgTkrZYg/IOj
bCveJEfW60uCBDjA68jw0w9TgtWt0paglsaxHEmfNfkh0gJNfiuLlCxv90NKyz0zzmS+ZZvuWm/a
uVIlxNb3VefF27i4k3Jo8ur45eTS7ClZw6ubqPMRTFzjpal0/eFQ9YeKMUpIr4qUWhhRolhLQz5Z
AOgzb5jcaeXZys0AMIhZkNvbuCj/t6L3kokhc6LA7Ii2rlQAJ4t/q2O4dHbKWX/jOLTRPPBdQ6RM
dLWJzlXD0ro4t6Z3q2IFwdJvXx2S5LVM+ziEHWKCsVxxtvSbkAaMPbVEELKEGRTRkWOzBgrT0B54
O/9xRYcL4/76ygM45nzJv3R1U1qBaNg+Q1LJp6Ew4CN91MESTKI+7yeZOOgJFDI9DARH26IMvGl+
Fa/Zgz8wQBioTCNxgEbfqXw+c3amFADO0BQ85Yqmhi5/2ooVGskEdlwA9f/4NpLr/96mGB2hm45/
ggPvwUGfeF8uPQPmf9N2XHkbAlAKjLiVFACvn/cIG4AgNVq1el8jKWyzkqJc487lU/c7Yy88/YJm
E9Ld5Pj4S2QRmtwdXWPEqfDM8YgFAihfdvr/g3Q/EKRINtdQJXCh0i2r7yA7rgANr1D11inxyCPW
ittL46r2iCQF9MSmS2rdpURiwUzsvGxF3qF/D4hCLEDtoSrdJkTl0bQITMYH8D7Rt2sTKR2S42W1
ZM798j1Q/zUtS95OfS0rNybKJqajchvwTmA6hFh9PzbT/VBYFp9coiRxkDLtzvTF16q/B0tIWemg
2ahHgmcZzHk55FspHk1qfAClmmbAVhk8lILG1qiuHW65IhG3wjIgbj+lgpwA683NPXcmLBFpwDVF
KQU1LNcJzdHtaBzFGjrua2PBXeiywbK7VuyAJbmm22zemBSQQLWt3gEvb4Spg12XbeRQSnoclFmW
mO+zO1QNGgCNZIiGMQzL4Z/2zBvx5ty2wxDcoaZN2GDe0IGLNwfnpk+vqU9pHY3Y46Etx4Xys/MA
jGdUE3GNd4DVZK/2KC6WtmPkDbs7mhD14olte0ujllKQGcOSJFHj0L3EpMGWxdH4KM94fncQZLYk
AYp5kb4INS8SJIdPi6BUEgK0ECcjlUBbHVPo9hwsPGdBFhDGnO7tsPC1VjRHQdu4hc7QP16yhT3S
I5PYEFpaqecdoeRVV6oBzW1QBJd16QTVqZcF5MfyXZhdndi/8Ariyjk8tmxmYLbKfbYjV7q0/Sv3
jEVvLpab+XZ9wFW2GRJhscPsq6jw8e7LmdgVancUg3b5663Yu7sT+PbAnQOF4PCMiiTuruVcR8pN
Q7jtTe0FeNc803hFSfrtK4/ny2XSRtvqPEZlodXxW9Zey58F1660635BHGBlTl0kfLjwalM666O5
o2BfBVLp9mxh5ud50KudU9bt09bJ91CF7n5dQAkR3roIqpkRgD5cpahndRBaJaHvd+L2jB4p0Qjc
8wEF3OtDV4gO14K6Opw0ke2xB12+GVpmGdn06JiMp/1oymaAceB9CPJ05kG6DeiaEQTRlotGFySb
0HQ/E02aT4LHLxdLw64lh2Mld8w1ryxivaNGNX6sHhTAP5SY/9ogLFK3YT/TqGo1JPbRhERgnMmo
l0nmiqd+Loaqwy6tuvYF5p4buOHAGb7WNLGqux3b+H++7x0vc3QmeArVV+JGRhFDWsZBEUvFduIS
fSBxA4vnsh6NmpDZR0QjojwW/IskGOtbNW1zxIafzXNnKVpTbHPuQsjIcyQJfMc6rhIpiMITGn7Q
htRyfNkEGyI2fzP7j+1mG4enVxDbkCnVfB7wnaAJQJqXGQz97uNYME+mPpb1M3OedP7lJ0Hz5Qyd
D5NK1zqZdjXE1UulrqNNAM6bXAuw/0HNl4ba6ajeqZm5ciLzAeXE6FGC1v5PkwLHNsfyjjxfAg5Y
qSRsXzA5Evff9DjtXG4pJtAPtsMQvFhI6D1HIIqv0394cHfENTyiZwFBAfoIQBdin1y/rrVqf9uN
oS9ZO8fByUDoOcNejFXTEpmOH2jC71wvInbPeDTtC+JaoSC97HbHyfWfdHOZa7RfwUvxyRVwlq3x
uOG1ptmm+s3vnFHpWJkBoo2whRtxxKoS19bili3kyh7dP+rridwmTUd43v3rXsc8d0tdjztaAIf2
A3Yuu+F5GTI++AtfEDAGnOOVbA96fE8P8A4DfnrerydMdoJUSpDkm0vMaEGeFGAKS8MCZhCND/c5
3TSW9Q4hobqB7EMeLMmHN1IA174dVSMF4YxU6+ZJOcMAKSke8aGjj+fWMQmSBspLK+bxAWAi9WbZ
sssh2pNW96oaPygqbPzXNIPmxZ1bPchAFhjcky042/UkQjwnfx77TtuYHLOCOEHw8+QYhN/I0fjb
UyYOVCsac2G47RQoE0vhFdIABEpV7VJU9gPJ7Ojhr73WH/jkyfKm5+GfvzA4gIkhSQDXBKrOuXOo
z/lD79/jOO90l+4l0wfehxIYDTf28xGtnqCSKjk5zkyyNcn/eZo/aAK7VOrRDBpD3jrvZwrY87M2
0zACAGiWoaAxjWtiiVQnDqN3cWROLy79Y5Wpx1Dj157AL1foJPoVr+JxD/1mDB7mdZDpQd1g/MuD
9PMO4H3cCLNL7mDzrW0cn7vNMJ+W6pe6SxJDb4qi7c61pWJeDhWgOqtui0BetO3Rt7NGH/NcLiz5
6uXZGJK/MgYVSOh0H4rgnU1X9BdmYRcWXsQC+WpffnTzAWq9NF/l3rU4q4XrXom67rHsP6HiIPA5
TtE5qEslcOO6Vc2DTxP3kbLmxMXxjMa4rO3ymf1xZX56LmH9ZN9RsJ+jYNf0Zsp6x0a+pQ9O2xhA
VebQlsMlZF3yj0YxFrCnesM9Yse1iVJaX3jSyQSiQYs4PgpigE4l/XD0kPJpqVA7OhMFXgut3oKN
2VdJ/eFIK8c7DHEv5PkKrM7GJvlOuYBwGx/DiUbED/TvP3SYqx5ghsIQF6sJgsTMvw+4A0VjAwtu
y2cDr2XnNGbgaqZMDXUBkjZ3GAMmTnvGPEu1ql9RhKS3MpbassrpSFkgiQEzM51tVVBbrnMvrMBI
E9CW1PRkqoQWBRQkzm0nZt+4Y8WCjm+Eb3j5B6BLDavqv+hoXseRB/JNfWND7po/0xc2KEH9tXtQ
AfaWuaNgfj4fktL99juOWhBP3N6k3ps5aU0tzRTI1IzzyyB8elS6kvuScUZxbgNYYKoitQWGH9Jd
fkkUdekL7+o/+1NzedykuE7VyGFOIEoUdr3ZyUas6s+gdBry/Q+NMzJSAAI6FApiovAR28h1JevZ
zRJQ1d9w/TJ97G1lVTljFlXUTjbgXkgusinzwgHX85ixFo1/yOqhjtPVqR6xlQO1oEpt4E+uPCmj
El8cnQGi6IhfbLk7iNymhtyXw9jJCvN+YMzWYfhppiAzctgnP1bGg0n2wv/nyuylFclcDflPbTSY
7vCqTLhDvWTzI+azttaZeoFgmxL6KcH+Fk+u1UrwX6HLIHaLnPJVhpjTaJlhpzz6uNsG0qpUqxFv
Xi9KGoOhJ67onLDk8/P4hAE+k+1nFJyIxIx67KzdqAhi+YiiCtdskrhpKReqvOgOsoRHj9nC3vXb
Qef279iYUg+bJrHh73gi3QeCP8+ZRiIW+udAdSBOQajo2fuZntV0Jd7/bNYr2k9XwwJy7kN9GWj5
8xHuk85RMkRrvhLqEd7YkkSB0QO0oK/TagkfDHTLgSmIHnDEru9giutlsxpDGcz0hRqw9lXjKdEa
1aEvsPOXEpjFczZRWgm4Dx1vR5dcSL3llrqDgLLmrc3nnKiKdryQxpmZFaRv1hcl5Gz+Kt+sxYAA
8Bs0ptTXbQVk0XKG20IFlBfMPBeY8MVEjmkcLF33ZimJuyNSQWQClTonRJjLP0qckQtTQGi4dMEe
DgNJYn43y+Ijb5CjkqiJfsTWUI5idqkidvoUpcMRVoe5Ckh3ZIDREWwv+5GDM3L/k/U7jb1xxWhY
AOpZ4HMNAn0cZvNRTkBWlpFQounpXRB89jgPQrYPtLw1afZ47f8Pi0sHlX+1O6Hy4vd2TwxeMNsp
8l0RJtaiSqiy437JkAhJVtjkcO8rbikDhaVgTNQ/ju++wosi5VUVnmR8n5fALiowRhYO4VYW1VfH
3aJBguwPZnDspv0UFX3vtqegEnhchoyb0gj9P6xC8iYXVTIKI9pATHqbAW9PyJKP9wUsvxpmXQxF
W6yzm/f18Upn9k4YJbuhzrNEOYs+2c2EgZLabVQs/eHeXAKLzaYjSPYgeeUXu4HvA9pk2Q6U2snd
UMY33HtBi8bvb5VY8E6NdayVOpD9xjkaO/lMMoyyHMnDye/0xMMregSyp+GE6weygLxZtXVlXma9
HEP+BohUJL+HbvO4O43x2ggj+OKGNSSAuQAXA8iLK9qgFZwDV+XFcYLMELbEJ1yFyC6e7+4EzlOY
IZDHHWIHIZ5SAuXZcf2Ziy6PLsK7KUuWx3SZDeY9Tyx99T5SHgZmRorc8UiM1Yu6xivtlQRt73yu
+dfCJ6QthW3Y9Hv4Fstey3aZKY7w1s4t4DJWnw4vzOenWOwFOHjfF9BznOZN+52RSBhAbRLz6dWb
+CZEaM0tOsKb2m4klRStxUwuCK2lD2KnhqaJ7onyGZoV5tnj3sXwzLf41noMDdrppvBDVcJvDiYY
ea3o2iGL3RoZAqruWwZ6ZNe7RFx647GkZ/s4/VCR57RP0v+hZ2n/Eks6QxDxh40Tnh0ZvTdnbfh+
4q9ywvpcjsETUWZ6Je6FsW7vd6ovo1xKGb45GWW89Kl6SfxWLjXHLngQys86XUIyE5c3cOiiUh4Y
yzd0sCJlDRCeUGyjG5+IR5MJQCF1AYl2Wyr8vibks6fyCYMtuVfA7hQ0+7/kEne1asplwQ2vwn7e
qLzhaARmqgkwyN845kGEinXpOcL8sJ3tvXLb5f94/DJW5SZhVCu9Ap2qaXS+puhlSzB9IK50I4WH
2/IL5qOTMcDxlNgOguOmQmktddp1JeTDqyssqbriI6OtcX0cCBzpk18KflLKoGsfN8Kayv+wpRrH
01e8g9ECLb6Ie471ihnm+Cn4IbvxXlGudHC1GpKFT8mInubq2dWmGdDznsjXnCEp5G74M3jJNrGw
gmKgT2i+xGLWLWWSWGo1CYQX91gSrF2dv6JXw6ZDoT4xarGLi+5hngYxlGhoIFxdrLoLLr2RvaVw
CiNLlk319C+tSalaOPBIfP/eqEDbM3X067lo8a6wryAC2pa4RfzBBSIMYcne6O6ey2a6mJf7jsZV
QmE92/ZpUOazqY7a4HrGfUN9wHnH9r1GzYQuUEXsEnznvjrpMIkoDWEKNLA1VSw0SKknGFuyIIfh
5y9WdP5MHQFwAVasXmipsXVl4857Pg/TGxCFjnxU2utHBkbadmw7Dg/YeF2kYt45MVbtwePUwsb1
LZN5+8HgBwomKGOV/6nK0/ozp54/MjjFzAO99iQbmvAmtfV5kxt8K/UHuIZyu88/eWxAAnxWheqq
fxzysaEpH79snWTvjb1/3ehUne9p5QpzDiWwrjPG74zPZEsrspnCp6WWcu5KrhUgw8QIedNZ2SYA
HShSw6rTHuTNATr0VWsymeKi/vR1JJbjCgg81UtH0c4jZKQiJ6/wg9oNtrsUuNizOp6d/SY86znD
Ggqgi9f/kMuxnrW24K/wHPlMOlyJip0zLU9Ck0W3g+TWuQn7zXTyAFM+KM6HyLlDX2DcQNyPyy0Q
DsWmEjXZRqT4PiG6Bs0oWU+m73tJcUVWYdNW+7D9xIIGYDF/u8Biy1+rpDdt1e8wh8FzcTSP89WN
JVVIM9IiX7MTtzuGvOVGqqWgYY3h+YNNkyaANq6y9+vjuBUzuDagz2e+nnYsfSfdaci63JwglPh8
pACDcDee9yfQ2UrH/cdzPtM8YgCgyVu+bNNBVEMpiMCZWVL63IumbbJIV6fFWuAAHK8Gp9QX8OkM
XK9tyPjwzq2/Du8hqEl8XQBxxLmWWKOub/tDYqgailGNuhJOfijuXFEkAhcrJqMD72urNTzJuqHB
vagp2tmoIB8Y3DxdoqLm3dF+QrOLCtbbeo4bWuWlJcmPz0uWJ+KazYaLqME8x5ibSkIlfQkE22m1
OjpRixWlYEfacmqofy/acfB0vJc/8HLyKu3inX9LLX1agbBo89YCwzm6eC1wG9I587tMEvwMlywe
pEH2e71jXL8tzpK+Ntr31muRGrDss6J3I9JrQyZdudwjjnPiwgpNsvPmk/jXtc+Teoc/RMq4jZZM
rCB/R9m/zys434oCFns7+kLX3fY4BvdR0euj1GFcWFZ3xsRouIW6aeFTzsmuIGalKvnhvcCiB3pc
/8qX/7PHtgmL1taaWyC8N9vAhrSBUMAWhXhKVQFwzNa/dDGgAKgUG3PxmPUx9rHprcFfk6I4y7bF
S67q0bgHQ4bhHahfZDcpWLk2qjQmGNKXuOdgnvfuOFqnZ16mR0oOX5KqFlZVrXuLEnJnVAW52u+k
/G74NL1SSul5R9N87r4lfuYrdjpn46t96ojidwlNSea8kb/VxxDUzpMWaQXq+HuA575M3Q2r9PaV
eTyutsDMn6kXgcA22pysoV9dLejSKQiUw87slaXC1CJvu26kM9xEOLuFIBZ/szyL5WBUzJIy9qI2
bqrwwzQEpoyxSj7i61zse23nLqykegn9d/U1PvMgtOQvSo6ZrVs3AnQp6HrbAyRanUsBKZ2nhdr+
IQm+SnDZNVSt9kLuM1RoJPfsqJh3VBxDzt+zVv4d4+BQaO6tGb5P9PIZ735uonMxlL8P3RsiPtxA
hFWEGbmLODfk6GrA1xOs6ef5OSy2z5/aZ8tzm+ClFtujp/bvfND/VaWvdxONF6p0lQURNgds7qRF
VcaBc74BPoV3Pmuds2FfIChjldZQDpmXdj1UOYd7C0xOFQOvKhCiFcbiqn3RtWEVJ18j6pabkKGH
wFfaKRlS+0SRpbWKtZWS74P7k9bn3411zMM9uDcL/AYkVXacGo6K4vdZKkyEwxn7kUtVKokEtYET
BV91WJ7xJHKDzQbTAterj95YOKzAaMLnfksaFpAFkY5UgBdP6+1B81KpxqkvJi9MXYJ29vDiovRu
cD6bVoYlvoKh3xHcePROtbvum18shKeMCzSeKsG0kLVTHS2fz4oKoMqN2yEvq6uXuUf4s7qMhurb
EjqSdvImWwn1gWFc59Rgv0Zk71RbvIoxGhugYfPfHt7ETehnT2Pd2RbeyvvFiZF+lWdOfRrF7V4c
sKhKQGCw9e3Idj/UvzGQu07+m6oK//DVr2gTXDKIz3ZfMvAncPtWj9zmLIcPQq1KdOjOpA+93CSb
vYEtOVkBRuBqs0AFZmpIgQrK5uZTiCYS/AqXMqUgpxbbio7KsCtpupanbHZTrzB5x3DPRsz3IjRK
5E3t079mEOigfza/y+9+78+2yG6C0tdalVlZ4y+AEza2N8gDdlF1rUGj2AYJGcNOAr750s8JxAJJ
uOkGW0yCl7zyfvOyDhLRZOH8Th4YMeWv3GmYMIqCslz++CtTQ6zLxV3JSfBW/FAU44tUQ9Hmj89o
Z53Ahgg1UxNAwQGbsdpJ3GypabR+R+tlp3WQcj8Eao+4vqd5EY0Vp3FOsqy4uuu9Lb7IUjAbzQN9
L7DHDCXPFco4Hdp1imA7tBIfnmPX7OQzwxtYpDV02ZZU+K+UBehFP0EZyNMfvvcTWMMYFjzTVKEP
jzu1GfzWonjGeTdonn7n8gfx7Rhk6Pak6J59kAEW1mY5vY+4/bMguGHsFd3962fAR0O0k43Xt9zf
9erKKuvY73JOLmN5alhNP6dhpOOF40YuOTmxj6VobAGQPpI67ij91GgLmmidHFE2Hyn4azEyzvPF
8dAVUb+L0oOEqq7tMjVAxly+paoEKBnatz/RxpU0dyiTLEKjZRBv2+0uvUueN/PlLvLVVCqKAwm1
NvkWSeO0weTjxK/QS4UVpEgT7cS9IKX4rNx2HaD3LSvahHT/LhMpsSjfcqUBm6N3MzpkFzcFB3Z+
ZzWnSrLm4Cwj8sV9pyhIVogIborFze7gUSRzMmSOktEYofI/MJo847qCcFX9GACvHrmcaux4lvdZ
SwlE767mWlQ46YNPEt6jHg5a1nuUinEy0hLjqBh9KzeuiQROk46+CF43tytExDFkFgs5CyY3YqBa
96pHM/jxcMYldX6xgyyc3/69HpErismNmJ80vAkngr88YsuRIqHPV/VwQb8Pspmfde+NdfQRaxyr
zdOVwVzPQpT6SA573G6YU94k4jkvQrKhKugYYyLyvbCdwNlg7d+4op/e5gHCRbl7gSxAmG065QTl
wH+felXSGDFJFOTAJHlXi8EZT5XlurOseSp/iHOPrecqTSdgzACI/XUr8yivaFhnmshNfNBftfq4
31FHA30rQPX+pQqdRwAKs/YNcFvKbYYVyBuUXv4kbyX6hEqOiqwhNshFbhSPKcSHUwRmO4SXr0RP
l2V8GS8kDnOyJJKD2jWNdQthVpaBTdvmn/CJJZHTNesy69RXU0xw48zzMN3D8aFLVYFbtUTTVUr2
/Xk1AJ9YdFLEC/uUgrR83zjRZUGcdyjU0AcIDgS7WaF2i5UOpUGi0gI0RCo/Pza/KAliKmJTHHfU
pTppThvU3cFWc1zK0rmAIUbVwkr2NXXOGKVMQcNksznXKWJz6xqe1iPA54JB/eusTo86dLk3MSHj
7kBbq0XOc/2+NGW4+ZvEYM5z0loe5InpOqZUbRI6oM0fEfF2Dvrml9q89CIjr9NNealNtjUwSKaU
JDLmGLrDKQB0T6Or5uMJoV7WHz8cDs8qLrmC3cLY2/8UV9X3EyA/9cEYOP/JeCS9oukZG7VHzm5R
7eIJtQO+ig+IeHuU5WZejmofoENvQt0lMpoK+O53zw3CFLY5jBZ9iw1hO2LceKVCS5FwoTqwBMGY
WSfjJ9Okt2ZUQcnfaY+FQnL7ogq3Tr8mUUxMWphrSpoOs7xq8zuCddpHUjLmMqeALQHuqMUgM0sc
O2fQUcntDKDDjuGkIxuzzT/w2otBtRX4GxFGNWEg+FPmR11xjxZoLSLHEfiN3Qd78wTdDvTtnBnY
pFlw3sstnNuEcaPojn2rqkFigA5dYL25oYhsSCvrqx3SRVII3pdfnX4g7aYzY937dX4xPApFiC1B
wxcj4pdVnZs82AdPcRlRKZT2WacuDNE15xBz/bToU/fFLaTksFPZBwD0Q42VZHQzrAZAv71UAMoL
MKZsExyRxA8h0ij/C5gG618UFjR6Nxd8/UEDBARBEJteNwu0hlkrZ+cly4F4X8oPtlekR3E+VMQh
IlVC0JDguq8HU0MiAavsMP/43IjkW1P/4iHAYG9v1V3HgJfAfyam5Mgww8dW+FYQaZx5wVcfnmtX
gaPv9nFV18RBzrdDNvbp5jNDQs0337L2BqxW0p19xuksImp0XuL11UmuMisf4jMJ6Ry0RI1GCjkG
8Ky+dRczRo1A7kWjxJ6o3aRsPw9b8/E4kDOhZMcPJKq3v0ulxLdUAXHNpnU7esflrCSsTrIVlU4n
llNXpM1URrYFvuVgmz84lcJzr7+KEcdK/LLHisQv9GtLeklFPyajQl890OcCpEsFbrYSYpDXxR4W
NTFfLVY0FpG9zvAwiMlyes2Gugc+vMt0qWL4oMxNUydNcwNgyEe3tCzr1qMy/zjAkb8/LlYFEpat
Vn1nhVONZy1yYIa9Yg1YDRQ3pmGrbhncQUAFED+vVzHSPxULrm8bEMHnvr+M2NAzjmZcN76qV2iM
s92xPmIFQdtwRQb2lXODMHdI2aIvdYm5K17Fg2wJlR8EwQLWop+eTQapdkBuqBPCrziS9OaGxZwV
k3e1nDFHoMzneJrBhAF7lGmU6ZSWsTTnwzKJl6Au7toE+G3kfHpOCvQTXJn3BJ1Gwffr/O/iegQT
omg6GiEimXg99mmDDKsx+J2IPAr6qNEdNAn/kgAsmjZ98hndOJtemla55m94CqnDOdkqEDhcj061
8mHbR6FYmm3auRKfbG0VwLNkuiyXLfEl1/epf1PnlQ4ipmGwm9ZBvv89Fdn6FI1E+Bazzumsb7jp
VMl9o9LSnTzLsw+VPANgE4yUfMOoMGcA/TJcQQhBweO7lB//P4ScdgNYJEUGrwBxLkbyxZxu/6EV
f4L1ubWBEtUopAdNE6Pi72S65wjJKzeSGGJJP2Z7uHricVOTflyBE8PR5QeGzQ66TBWt4FOmdWlk
qCH3LvEhtuDSIdRAQPhuowwJ7rT0R17fXZgtreJu+HPi1xwufZOHIG5ntnz/Km3x7rkZwGRN55Xj
dC2WnV2M4MB4yi/AEpFXxVfMAmLjd8Q0gBix1leqej3Ov5w0tgFlE1kRnhfHSzxIWDSf8kTTwb5+
uiGQXJeilDFsVpf6qFWGv9VJzj52w/vhPQGXzxyInT5BdrPA//DJ/IjSEMlKREztoGTz08QOdagx
+WY52D6Ifz+rtDuGYZXIkp3h/4Fm29710p44YhXHYa4bwHSh/IAqPqo79ACLPi2LVxLrWp2GZSeV
AL5mhiEsJ1R0d7Ngy6r4SWJ8hjEdF6JrcCHQW268vF/oNBhjFVVxE0ATcfgLlsnMvPQzxxwdjA2A
H6kFSPgbyxqmdfR9qCRsUbStXsbPqB0mnEo74RyVyLilxSb2mpCMQXsDApz3GELBKOLd+v2iR4rz
h6T8Bvp3u/N8Bv8zyoRpGJGh6fOZhiQWI+i2vWGHx71Mtf7gmCSemWcrlGIgxtRXp3J0Tx8L4/8d
vdp9fGoGUmdkQ15E/hGihBUAcTb217kcZK0WN7i/O5wQ6NxpFKH879gWMgJVXVomhCRb+jbhTYYH
1r1l0jTROuPQ8GJQ2WyB3pJ4lwqFphj2bDnM963t333kVq0Y1e0cpSHAVpAwi7rt7Yad3+W+M5lw
skQDMHBvR1fcsFxTjpAVefPfQMwY62FNnUDb7kWIMPs6B5P1uJZNbnqCFPDXVI2UEAImUKupvVJS
RDSRkPW+ZFK4YH2hh12bRk4oc/W+djrtGoGge83o10kdXuQJ1IEOSD1UMd0UmGtKjcciIRSCCUsW
mocMyH3tvSQnmZ9Kndrd31sw+HelpCypCsF1C/mqsLBsFp8O+ZVGPcL1sEw8kHCX0l7TCQ7cTH4g
DKv6PW92Ujg1hQAEhgc5++Ex9LgJKGngfUmwI2IKHPgqAhhakYUhvdomkTWqmwOuQwEIP8oy3nUm
z4RMlfnOVPgsiLuj20AgxU4+bWWXuQAErjYn2JmLAFZVba4b5l8cxR7bXxpyCMIAjM8JpHxJca9X
f+D+8UJIIV6zfPOmIVvV0GqAhGbYKSPA+m1woXKBUUDR/WYennOqgmcu2Ins9MDYARyM7y0yDZz5
lpOUw88E2HrJ+2AHHaVhdN0p+HQ/0oQCLAtFy6qqG0w1r8K1bNxt4r44JCTiRyIEnnN0sjFNq+0g
51wf5UBukqNN1gqwEv6Lz5095RGUD3gal4t0RCmX94LaVdiyhx3NxPHjinOH8mwtq/h5E0vzcOrg
lXuXbBuNiaQE55hKPJu0hMdEgoaJR/PtCkV6OFZ0di1N/PqYHO5pf/wSihADwbhH+x2iu8cU4Ce7
og0UXvT4Mpkh1zS7R12WVZAs0iZbCJ1/tSBbWOcabmnYkAYnVos7KyN5zjqzcPcnwMTqYkCayvJ2
Z3IWytycdIVXQv57+C05CG1+TIJ+EeFfh1bdX7PxIcfzqq7TmeKAj67ELdpZziEHuTgbgeOds2jy
El0yAhWoFfavfbIjr4at3Jr6jp25rMVrl54aUs+7k8CkDUgFvYzWwOYqFASFm0Ri2M8odxnmsP7F
iMezHS43Q2QGFFhSFdDvOvikDpKbV/U0DfJl2zfRqb82eVxaNDLR6nc5sJgkaU+cJVQyuKPG3d3l
IZN8ltzHuEAVcWSRI1fkEhp/MtB8PBaO5zL/T784FlW9RPnC0+3fBgLbwlvLkp/hjiSuDrnJHMqH
Ob6c0gYG6e7lTlJhvt0L3fiqdHAekZBmz10QPVrKeoKwZP9Hz9afQ7Mptt+2/nx7TXxWTayL51C+
9zc9GTGAHnebJKdAZ5VM3+UQqojV3lkaTO78HzKzq3ZXN5BsPSm511VzN7mEQzD/XT0VHErPIXpM
vK20IZbQhBmlE2KvJaa1/shs2BSA5svxtQPhp1laufnOHHA8SUu3LpTCmD4fGcZFkM1j/civ2qHd
auSCN0JkByJiKLU809iVJO5xCgbXqJVDpMw25iUqG6RFPX94UJPMebBzdJCUdgPLItwyNzt6TzKm
kpk7tIncIue00LCdP3nzMFzPqxAQ8arPHLpaP9LGXF5S8G8gkVQ70Na0JxMsMrlh98dQCxhXz3tc
pb9jgH4z1iOBdjB4wZJRdQf1jpyWXLMZk9+g+/6h5UClIUeusaLoKJjzt1esJb+FyNNOzALrBPmF
tn8sbqlmjPaQRXaQ5yKLiA3f8gPB2LJk0ud8WXxpp2dgwkh6WW6OXpOAxvLgDoB+DDTCTJcgJ67Q
IrRzQBhuJHJxxinqUm++7ezssUZFvOmqzKZnwYNQ5dpszXiA8sEsV74J+KtMc/os52qqffFBeSQs
AWalnorU5vcAynVlrQr+YcMhe/6eIJrWIcHCOwz1Hde57bqdG4aGzMQW9n7OpKpUXvaYRisHv2hj
Bz/b1yMNW5txKmlxCUNNKPkgXLhIeGZS6eP993RzAfTr/HK8uXpsmxmpWRFfoWHRSl0N6kzCYt9i
ZD4oYTprmPizTognrrWHSapSMfu2WRR2HqdF4GpXW2bYrk/P/y7tKNHFh3q79V8GPArvFOqW01zn
aTFmQZQaXFZpBuFxKO+XS2LhY/dE0rTW3cFIgSjfwQx6yabsj4It8jNUpIsb569nA/haTj7txKR8
bOpMxG9NDnQ/l38RduhgwSGmP7B3jcbFoPHvdv45FzS92mhgfKlTX52wfdTzBlC8M948P1VTaCNu
iYLsDaF6XZJN8YCtZjaYEi4jtCuln3whxZXs+WiNt9n3G2gCYAagDVWyUWFDDo67TAmq/0wSWTdH
zGRw0XX7c/DeNocCP/TL1uK4gXX9xRleDf9GpBLaLDq72yGXtEWMErqwagkc3mHJNMngQEtyKRQG
R5NVS8h9vAsqVTJGpTycXLtRWzYChlVyq8qFNGTbLnzjrnNE4WKMtbSdOwizvLzmWXialRmntLE/
Ee+o0mxeFsYMKwIJK3GNtUCNZtJnE8KbqztNAWJAZJtctg1tfxoVDSCgvFJS29yvmdkPSJmZ5kuS
OfVB8jP5aZEMw6Qp+gqUUM3OegQtTrBoDHyr9RIyyGq0n23jq7BRZ9JNnWdOgKWCdIb3xBPlS8tT
YgQaMcrfYcD/b6zQP0FHUaFKJRzRFwksMyxXHB1/VNf9Lpb/E44Twrg/hhThP/cDkRh09Xq45Lj0
IIb/QIYhw5UaRtF2qk7m0c4YvFSwHLy5AS2V2lZkCx0v8UbAdywLPkHthdUUYsvsqPJkcg1724hT
vX53lysF0oAfc9pZBr+ixUuCg8AwmRZcjX/Pt9dAkauun2rXFaB9Hq7e2tP9LSPH7glrsen1BDGe
rU764dNF22xLXF/UI5o+Iu8BRvSzQfSegEbNx7Zh2PtXMlI5vE1bXrCMMZSVPS8sVkkinscDKsHI
dUoomsjDcknn2GPfiE+cDdUOCn5hHjx8ILW6bkAm8I+3ROkOWSiFmx2kB/3iJZwLqcfN9LVP535Y
lw4dkDMFw1aSBEcAwovqhAWZtkxbIabOwnhD+5yvoHGCX2njx0J6jN3nSJw2YIaha/n20v/Tmr3z
M/MurrmnIJ0d4AUbD+UWVhI8hK5OM3bPiBNvUXSIErlZYdExcwc1Jmwk/upYmDtzHqqAov7T/TLz
jF2T6fTJ2YOkXv4oE6xfV++kF2vlqZiN0B3UJy8teYLE5mF0/W5XRsqlfVbLT/2P75WdW208Mxq9
YVKopq68CknBD0/m9d9B/+SmNRnYrpmSoaUBT+dyLoG5ic2OXl9MEIzq6jg6plES9fjdMjkHerR+
04uX8zCzQdd+7VovtgQJB0vFteCWewu2JNZWlnRpWVeCWN3AvsxEe/7BT2vHeiZ4DXFf1947+8+5
REKeK7ZXcYlQNZGkOmmYNWILLOi6nhyeXvZQX8e1adCyj2ao/gC2dzgT7pPpS1X21mi20OvVRFAe
wVh45gP0JkTGhVYFXOl+6czyFwRIkWJP8GNFzvPk8ay4803oui9hh384Qr06fWCFe+0sBoCtsk/4
CuSSkzKqkwVaaW68qPiwixu+MOzxacrieKt2eAXNF3zmSLwJzRErMfDI8SJlte92NeKOQtAIBexI
6hU/q3hQ3Is4p74pxGmHdd+8C4RViFsgaAHexi80cPfKeqcJKDOH0soWUacf63uzVvI8xtqpFneg
RMjAK4H+nfz5/IJ1FXJ0D+jnVOL+mY2JWcPYYA8yf3X/sai8YCNxz467O0f1xeoX/J3kVBalBjKP
KaeoBXZRB70r5cqGaxDPyawi/Vw7x4bUIuI0j5+cRq4e4BlEr6YMjIz9esqZue/tSL7pa/ziozjO
WMhwLCUHSyEM3SnwitkRn5FNpJPVHON3r2CfgpBygKw1pzAdtf5Et8hxuy1lAQLPnpOL/OSf4srH
+HlG6mTmtQiyysNxlt3/GFHDvV9yg/w75rZ7L15uuIkZ2tkfufGJK3vdDXJaFKEkwh/JldeWUHpO
TyhpJW6rIiuXQpA3bTgqiIdGWtEdF3PHqV+qxF/tzzqaXonaj7jSJ7LLWbMb4ubF6yP74iYTx3U7
Fh0QqdIHuqZkLSn7yoZp99x4r3d1NwcJLC3P8JDsj5+v13FWaWZHVkh4LdSd083PgFKKgTsXkzg9
lw1IeCb6GgyQ9nlY/VNoVysIdaaLhPZTGn8UrRDu6fNQ9+AW7ha2qxOmUPKrgUkocUhe91NObSqx
KmUHTiSK1tJ7JL4d5lqPvCqZAWt95/qamJwJSau2m8cs0yUjG/V/emrwZexRdXOnXLvQjSBxZ05+
FhrYn3yNjggDksKXLSKWiFV8YQGduieUiYT7WNt10Cm8pR2GmWJxRWradQlGdBe/wmWA5WRYuR+R
KfPVy6UHRvinPJODWywhgz4GjJjcx5Z2uypzmi5AaCos78/knGW7P2CK0xB2ahF2OZ9SQYB0Mi0v
R3Y8J7k8AZyE7vGh3+gKuPZVT2EIIu9zx0058MKq6SvzaqBzELK3QQqcMo9zFvlv59978b/EyUZb
EGhxtkUXp9nE92YmZzZ9jfTY71g+j8Wz3wtzwFFR//6J2gAneVn4Zkog/vWQfry89GediZQDKC3Y
7Ddg+1lymzBdweIcrQ8nu6CBRJoVGUoFh3BrJpXr4+lSynFkYLXc10z4JV8ZsfmWyUDRRY9bouvl
28Tp097TqX+bYL00wFX0Ph+eFqMURdlKGhQ9HvxRyfpZj3ZgdNAlcAN3eSphwv1fBHom+aK9URlM
/RvG97CXSmBgvDh6gtaPa6EY5I/IyGl08KscNWjkpHT+i4fMC0x6oonlQNcFfEBf6KP+G/eRVcTC
/QyTexqyBs3oNd5oeAbIXl6mjT9sSiABxGqwatTM4C0mt6zId51pmMypQcuZdN8WsmmHiPcDG425
TBJQvthy1mbNNAKBsh0afT869hnXbtSW4zE64ZzszIIlN8o4tFERmAwH3QAHdXw073trzo1jI6fC
u13PMFyh0i9Zd6ixEdAtqTBNuQOBkv8+1sDFPNnwIBgJt3/VPaOWKyiE89/n38SOrZMubrsAPm85
cBN/6scveF11FxlgGyPlWbNDMnYue5XBSIEYFwkWptC45KwugtWDNkBEnzPhYniA4oyi5PM5roKq
FNbKBiJ5+Dx0SfXxw+yXWkBD7plQvTnmfasQorRVYDpL2VDYoXcQ7Mghwi9pkWYnST2CglW9mQ3+
grG+ZwvPJuvXV3/j1RUr+alL1eEVnjzLKeRyvUGRrFWHzmj67P5KgX41Cyheh66YIf9XvTtNhbQJ
w2vHMAGbHaYydoT6y+x1Mp2LyKm0PiJsugn/BrIQzNmPlkM3niRPW6Nu/Vdv/p0v+5kXgTV6GuKV
rsPoz+lIji5nkjJOABBdMtuyrBMeJF99vpnsUgO1q7RyH8ecaZR1PEZ9Qkjp5fVJLwkzfvkYWCZT
N99e5WxPsP+b12ZC+GH15CZQctld3yiA70iFJElREbc4UGK54yhbbBbGyxBi5FZitBl7sfuo0/Ou
ZEIB/OICb7YLYPD/+jDza2DOInKyIQKKPnQLx9N7uF7pnpwshqAQbQ676cgChX2tLBupDNg51hYi
zAsd6Pvk1+tS4C5YvEiXDarz12IeMvFTpVE4xTUUBzReY4zF+Z4FPFzOXNMXzfik2HXO9uWUoc13
GLKq+zqPQzZkj3l26d0sDb/YVEbAjo1i3AXrJT1O39MZaD/vpnqXbO012argIDPEU3hXnDUxwvVY
1CuhshVu6/UF8wPlXpHs5B8ivO+gy/j46yTkQTQiSygYeH0iPTENt8cb1kO5yFOo4jwNiNYzpgzl
5MwNHlrdfiZHUBtwlGzULLUbIb87gAFoc2lgfktswH8EQUppz3b4UMOKjzvlV5h6gRJwOdidgtJI
Fo7BUwoRjWMduu5uETbNeV4Em/AFYyvUaq6UUgHhqSvkABbQTAq7y/qIWixVjJlH7s3tZK2C7K9N
0B2z8kTmJiXBq83XeH2pARiBQ5HeNxvE7BD1Js3PNLG5xsKyMTxphGflzB/HUPO3PuNsZn8ODzNa
5+MV7MNq30+2PiCEnZAY8a8T26iEHMCYnSvp3/S7qoXw6TgZslpmYYQX03jKWt5b4UTce7KXt+90
rse6EWmcHHJ1yeBO6yu3A7adDZJb5Kp2cGm8ZoiW2AosOcXBQHEtZn7pfAhzrw50A0ijDYQO/T+F
ihlDTeSbtm7slP41onJhvOobrwS8N0QmalfXhWIGH/yWbnJ8hpRIRwvjQCSQr2D9faN1p8x4Q2/n
LK72HgqST2txIZQE6ukm+2FnHyahPYP+fXzcUAbcVOdxqPwz4sVRaiDKPTB20fE5t8xoKqSX1wD9
Br0x6tnoowTwW14XdiHqQV05y4meA5SkN83mbuXq9XD7K+DhDOOrjxrWaC1ULy/QThTEZK9h1nM4
1NBwmoZ3iK9/cc6VEfSMQb9EtDo5+QPm0tHYpofuErf0VHW+J54Hxp5xFADg2ldrindUiVtIGmTL
6NOoNkBsvnR0+q2D0zhDMMayKtrrtxvAYeJvW5ABUDFjREIR/VOZYbi+QePos2/zzHdVE9k9b7Vp
hlVA2bFy1N8MPlEejgsAGTAWFwE7dtnH4gURsZu0X8ZUmyssJM/nTAZW1/mGqHmWhiUssUrQ6ItY
S6pDD9BueEItUV/thqj7wwCUGVZM7MDo8n8RzAhOiJDNNhC2f3u4YLNsxw+M0HQzIrTxWyX8VMP8
JRsTPdYYGJdAKRu5KjYFHOVCTxBg1R3KkP5jE3e7ACQ1C8EwspY2F0W4BTB/OoU5PAY2mOT5nNOP
9uHRQvTUjy35GlxhpidIqgaGukzdpRmQfvucx1OfmSIOTVSv34hDdcFLJ5YeFtperxP7p83A/oAU
jgrXO5nJCkgBzit3OGArxbmElsdHlRW/DcecgYji4Aq8So/6avIgyoWoEk4dePU5lm+utc6Y7qPZ
/HNnCMg9dmPCjDCajj1XQTkujdoGkVh/htozthN/X8HHQAawfAIIX6c3tEdmQrP+GUVpEjb6aWjc
v3SAXW/x/3eSRqdVGhOzvp7yylvvYmFhDc9a2dugarQJQw99H/Xcb1kByFaIel1nqKlaOM+/BbBJ
8c67mdlsbcHWSdN/A586VBPOOXeYpJcqoimeXeph0Z7wFOVaIppBVl9YApnJJtWjJFla6umAZQVj
byOeMTkqmKpRAX8DAK7KzqGdOF7sr6tLdeRaIZxx3FwN5211BfV9uFqb6W1qc6okS6ES5cEeXhM9
L901w0dDaSxrjSHidLajUOLbWjzQ3keGncCFcaWV1UCByt6HnfR2pi/y382sZwvBjQ0AAbFxGWEG
xaTU98qmFOVILCePuFIBDEOt1xVZ8yiFabs5tsIxCbWucCxLLNXuePFsCrtqeiplH/tu6kden97Q
G5b/NUqn8XPRUDUu3NUcQoOrxI0+JfRaVLpl+bZSqWQlkewq/QRv6Faxzh5Mi6lhomlTmZucwfDo
gSz7t0LE5FL8LzQI1M088Z6AtpcUqesndn6T4QueCoSsgacsgdhgL5wChWeUdUKUAASWBDivI3cw
p4UT7c4jz6r1HidfJJ1Eiv2/sHo8+Ef9+cdCztczdoOqaSQm6tl06VunKdatLh3Yw52E8hDjHBhN
JOWx0ZYGKpqUmiNju+xU7UEWFl+VvRCRW/Hz69Uef01XhCykbdbTUGtDWTyfTAvml+ocIsb8/kyD
dHJvVGppnLD5Scf5XOyrrxAKwWyV6YK8tBCGPUeuybIFK0NNZ2rAQ8b0wRduXnnd2Sz6dLid5tAM
Rfj+EeHQWJ0vylNYt6F/Q31o4EQPBlegREwAy6LAlIXbJuHl4kREGdkLIHjtp+GBDmptsP6YXrkn
mYe7c9L6it5wNd2HEUZ4RG+mazhLNmmflynR2V+4FEgup+lAUfWz92rxJbfNJVMI8mL6+wKtQNq4
vNRqB0IxaB0B7ea6PjXlrTvzj3EooGCNjxJaxTZD+59XOFcRFz+fYE0tNIjQb5CEWuC0UCVDKbUS
JO6GMFvA6+d0dSWc4itW4pR7bafeERZzO6uEDKOI4dyeZ90CqPjRKQ0W+ZfkjIrUxaE6dw7ut7lf
wEoRXrQW9RDB/1MppTrMtcXZrLSwPtsn/tMYmXeZb5lzYA4WUxtapHM0vK4wXUB6rqwsPMjBSOoM
WWB+OZehKht45LOvUGk/2Wlyt+I6Nyfrcr+Kiw8RHuaOn2BpUoI61cwBCCGN+bf8WiKP8tj8x5OT
6fvmeahMpBvMrJtEuTyALNrVNqfAOmT9YHlQFBGjM459bHmLgkG127yPnYXOaWGyMotLtI+ujB5m
Id9z1IeztUeImrQUZCaAcUDGRBovQ6onUPSAK+e+5aUQ51M7rDEXgJh/eGpfzbqWux8IRZXM4hx5
zac2la1p04qLUVwsfvJKaOHwv+rs/AtIBkSrMDnVvqswXg3iy1vUBmniz8/lLdcJN8dt7GBpI+4U
ws/xJ0dkTfN2CswFFeFpwhzdAXu3d9qMXaxP+1kddeauxQT8bYLLBSj8HQohrDMYBuCZp/knC29u
KFKCJYKo3cncIclhXaCZyn45OHyJzwsifzWb9mcCWBKM65DPGvE3lnbkwQuzQAbsRYVY9VnaGKSi
sI3Hpq3O4BWXtjm8CSCO7HfzFgfz7vKiiEXFoJ3HlCHmkHDbAcKqW/izz5X37Wrp0730ch3eIILa
OYjvJx5VMGR42inKKcyBkkESl4QwYlw9v+p4IHdIscjB1JwAYzmGP7ZKyNuiwsF4QqMpZkbR83JB
NYrS9Yh+BOad6a52yV1Q603Ngd8y+NL7XSaQmYlrpstH/lmWiKMOao7rU74VpmD/C0cGOaKlRmg9
kJA8o5aU5rfBpdAqBckgRHcAeTu7I/4FH5ByGXKz664W56QfV31AOD52x0mYkQvL9+9AMAUjVsjP
TC5jreeV8OMOGWrAMSUohIGjsg2eOkiE75aCxMVDAzNRqWpT4sXXdjSnhyllSGyOUHwFB+CtqilJ
6/LHj2p+HKitQbX1vaTyJ0G5dxQBGGXeB0W3iAd9BQTYhj2NoftnWRMwzxdVsiINUd2Cxbyolz1v
0GU8b/Z/HQ8OlRFEMGAUPI+egv4WT0WuGD+YUum3NEcGnXokTSeDckcrIqrMmqB4S/EWcrP+gkb0
7jQjd2qiDvY4k3mC6LubT3rark9mIcVQ9EbL8Fhk1B75aQtFHQaf3itik+VqOyUdSbu7H+t5h0j4
ZWQHLrj2VIdJosjarUErU9BY9/TmvfsVYWCIVeBhBAMlSpKjA3y61fMDONhx1BsTjlcFIteAynKm
NdAjxsWtS18NpSQtVBhliCLL7QTjEbinFT3MJDvVmOlShDCQPFNNS2znprqaBIFZ2rR0NdaaAlMp
WiLWCJMEoheUT8S2Cd62cRM4xcXuaPHNcvPxwY1vDe6A8AMvlhegS2dFaneU2DGpcrXdH2pd9fR/
3ip+Derw4PF2Ek0A6yFBPFWKcEIosE9LJf+GVrYMXb9rLoZa5LCzfa7mVsIpMkhWgqQecMSpaLY9
W3fDFwrmpl/mxv9KnfSruoBiDhbVGY15dJyU2DTlD965RW1sa7KzvJwAYu+k4i4YmoQQuFw1hypl
Ngm9jrhILSstp4b1iv/WLRXQPG3fD3fSKg8gnaslOt+8NflwdhA5JrHm/gTY5vysA7VUlhEk4HFK
X0EkeZQHLSP+Mq5otczxQ0sS6Z+B67lYG7i5o15f4KWurn+y2HHkD6ugz/n11L8GQsel4F1ynwEE
vXJ2WvMVq2cep+dGniOACG/JFqswShppdvMV2slGCUscUOUPkMXrGGKIRAtOXdddLj1MMdtd3GqW
ASLSLiDqXMU0yEtkUzcFsucz/y3aAUSb16w5rsSyQRQon6Zz5fF2uM/5lXNIy7yXpAXKQysKfbLt
hDr9YcWvcD3mYEFqpMXH8AhrZmh53ZZrhFD80p+93pwe2Iw7b+4BxlV3lXYIOHcojX8rCBJjaNqE
p4tFadoT14Q6y6qHKVoCb5SZLwXlxSwhx61wnygmi10NFEl5F9sIjN7V3T+38ls03XLzt0okCLAI
JZw9flwChoD1s3t7YDeySKzgDXVW63Rhm9pAyTiyqwSolnM2v0Y/FrX89zjNV8ifK0jaqdyl5J6m
lpLx0tPzy1686XxWDrCLfMxtZ29sSPABXxXtUA6AtfSz3iWPb+Gl/uzugIhzE2loP62YYIIOnVJX
I0qzY0XV6+/EFWAtd1rsNt7nE0hxiV1/FpHnRA5xbJOeBGtCm3dsNY9NlM5aq/E7+rWuU/Z1cTR+
7393PHylBYf9pwbtu4EeBEzG7WbQX2QXK6ojmB6myKx5ttOiPBS01n35MlAt8ZmHuDb5yCmN1OcL
qZX7QOS+rUi9KV+Szob22NYgbCqnP8xn/nooeik9O39nfTsCbRDs5eT7QeWV1j43Nm2geEu/inAA
AtUefZiBIyaG03hDkg+VOFY0wz7QBe3bLfw19bb+XYs1NvlJPgd67Qjmq17e0shehD/Y98AQ/bgG
v8BTPufaOkM5HmBhDL+NYdazSz1QbjvhyZZ2wcR8OAeMRrC/2guNmYhdDwX4gNIVQpZ+F/IfNDiQ
k5b0bjRfBq8a+EV+72tA4+z7SwO0gR8kXY9isxG6Kj4LALdJ225/0Cn5htdZ7IWH3g0My6VZDhWF
5dgiZ4bIxivYNENttVxUmCi1pRoYvk2W5TwPO67bQy1Nkfx0PL9zCrVzsCjVmzbxjVsGlPNUio0Y
Slh9EpUcLmVGMW0oAUivy5t6Oar5N24AKVFm/6I8o0ttejve6QBU52uR5AIytIiicceW+kfQ4RX4
8jhcj8uHiTyFI0cgemTcTcC9ibWqUfE5U1YwzEfF65JjZsxxbfItWeDQac93VAvf/KHg5ueePETJ
dcMmAkilm4nKL3jO17V8jv+J1GrL/Fszh84KMyaCjTvqV30JA/nUcuIQGW2sqHfbk75hW1igw6xG
7HpCOmudVMz1U0Qo4gpThGoq7AtJvae9PXq07VkMTONyo/2k2piJpiMMc4Ma+zlOnCJbITMhf07P
pr3uSt2G8oFLPL9t5if4jA0JNepLrcXQPL05BUz0mlR6RypGC9TpCL4KqvuzClGI2z9lrZYWiIZG
/HNVK7bCu/JEbfrRtlLHYVANFiQYva/ML2oqSsDwsGGfHQnU01ruZHvAqA3OmRfKBIi5RnHjlaLG
vYfLyMTd1Dzfo1quByVN3PU2I62Vg48FGH9L+9DD/DnrSzo7mZUgHk6oJreKEAgBS6WCMgInzcom
ox10+ZKn4pLwdJLUrmkm/x3fVO6BWvECWHElxR8OjvMFPlMunuoSBVwopmv/5IC2PxJR+R1Lmld/
vH1cl14WHdonIA1KFX3Rb1YPOLmPYsEuA7IJtMxMTEq8wGfwMj/g5T/ZcDWRAw8ZZ6U28ispyQ71
CtpQJTAGLDOWoHdxRigBKg9mw9ACtWxfMiFZZdWv7R2VWusg/h1iDUdGwDeLWPuMd7kVU7sTAUiQ
L5kyDvZM3A5JfcBWMLxLFwtIajYlWs+SMR8AAMUnWCuGhux1P04ygBJJc6DSPF0yvLWIg1Fn9EX2
bSyJNmhvb85XRN6BcvkFahakq/kj3GY7Ts9CmGnlOqhgvw5wSJA6SOV0m67hiLN/ck2+KvLpdHk7
n2sQpI6fAlny4xyp50Q1XbtE8y7NSq+/ZN+MkYr/WpS+dctYvH72sMAhpJgqpsfn6T3PSqOj54QE
OddhNVss1oqEgKUZRIj+Vs8qFSa0FdM0n7hBLq74Oz2VVRYzMZsQKpY8jXYFzD+bE9nzaedCy88Z
rduCYvYk4o1qN6X7e9OmlqgkHhHMde6iwkujPiDIZ1Z6En1swj2AqLjCUuCszRpuEkNpr6yMAeQK
I21MH0Qh6l9K8i+AAthNzGXBOKvWt3oDalYEsxA+naRe6gDQVgy5PYchbEjT4+az+4L4EZrlA7aK
sWHC5VmfrseFa7dHNzEzGmZcWcAlGUPz/P0T4pxZLCed9vQLEqqSvWbbu6SW5hfOhitZmga82nPn
37c74ZekVCZkao9uT0bQlVHlVoPVVfaJjvlRb3/wWxV2vNl5mI56Nhf+Cv5iXst989+e9Cvw2Bhd
So5OsqeTA4sfgAPDmerc14Xd2gnAS3MKHxo4WvMSNAQzThvzLa6u6LM8D7Ywta1NEV0ql7D20MWr
ByPvckxOuuHSqwCsquuETMRvwGfwquVjAFUcIjCPPYgnTB2crhW6vuh7dMwnWNtB+6MwoRUyApof
9EEFeSmj9/flJQznC7iabxenBQMZmIXI+1ICW63yf9XoweZv2f5U2x/vYOyPQMEfkxyWHmaseiHl
OiihWSOLpiAB8da23QdTG+WVVL15Cwcl4JneCk8M7UxhUnP60asSUvcRukJxPzlRaYSnQ0pk4f3O
sX5lOpEA2DLMynIg5yQLYUFcZlZau7yrg7Be+bqIlGaeptr8oDzaoDpoG2DlB8xng37wt1Ok1b1T
sB3FB3fb121XfzmeIDyItDOh8fxlwpXDDzcnxFmXIip/a5H4UAAhXz1KGid8CSjSh/QNrZisNvfO
FTXid3oqtXK/ZWYdp6OadM+KAhufuAZ9OBd9vGFTEfNmhYFDdqJFf9wud05DrT8MZuQTLb8OSYd6
gFzsb6jOvo3wJlQ3g2rLkHfWvnjq211E4lFygpETlfj8WM67RMFqNX5Jcf5goHnUppj4ovODnxNM
wDIEh1vpIjvzBZukDPDFR/OIPE6MN8/wNclrKDRrLVEQrWKPbr1FUNW+7y8b+lC3yLcXKKJQQ/4Y
j4SMtRlyNvO6OTCcEyOCkyQyQnzWnzuu1TZvm4NGOqyUAE/Cai7JtuZL0Lp9r2XZ86i3ONz01KYV
oU0IU57joYC4sFjIQLXksYdHpk2+IsnSMuLLh1BcwRXQlWqj42CXwOOqVByX+z39p/rLFR3fBuxR
126mNOsQ5RzcEbi/TXZMd/YIZ0MUCad0eT6j/kGmNwxdG4npPX3bzu/hCKUYmPJauzkV0CmiuOZm
1nPcWu0EcOAXkIyGgF397kFcTbCWVoekmXQm6U99YQLqmMT9vC+3aKhbNx9yw91VNUzf8XE4ogs+
AqCdc7tCJhDkPJMU3GhqeUbe4j7Hi3K6vJUdQKO4IYSxpybLFgAfHr1dbY5cj9w3e5ypbwuTHvZ4
2nc91FlxrE0PWWTHEEjrcYZzGlU1Iu4WHo+zZArAIGB94p9Daek+3gyuRezGk3y+qfKRABxHwe/g
Cc5SOIp5S4mN69MF4nz4qkArDfXNx1qfvFzEyQ0ehBTCsbQ4dPDDdI6Tke4TX+RxlOYyIgW2NteS
r7gM6d8AxcFZcDGrbe4pRl2XbAgFlwkngk/Mz1JTIyv6Qvu+7rRPRj0h7oVNYW7qe+jkFzPXJKFk
0he1gH7dEvnxCY2FLJeU3MdFfhq5KD0JATnr6sw11hZR7J7N47b7dk0Zdl93yTOaU0vu95OkPOsI
/5R4DJ/sj9QsgkzLOxorB8kz2r2VxR+zDuw/sj5DtYoXC5yXuVN9hTGgmp5x6SjUf9Ngoz+LD7RJ
7E+Pb5WZfjoNilLXHkwImWHEZASHo8uAYVP+Gzndz+FFsNxcpuNyErW2joSyr3bR/Ug4Gzd7NibW
Qf2ZpsUiaxiXeWF+hkyoBqgSk3poT6PJBTUHjHNA8bRqTleRDJOoptm/QmZWDR6Jg9n4XYuXZKMw
HJ6NXkX1WOiYTR1KQEXLSCApO43h6b2n8T9fQt7v24Q8B2FMw7Mu3BpQnxegZAB6HkSVlwqRnff3
PbRqJ7q8rV5NPqQuZkEV9K0pcmFiOjNz4rQU5vx37tzJWhVVPQWJ6F9pLwHyTWGiety0OoGqLxCL
ByqAWrI130NRd5zEtqTpaE40agTUnB/Rnr4UY1Q8n16eq338on6b72wnlu2W8nDOXkvaxOXJx3Wk
pL8MRAFuMPgFLQl+T+RHF485GhFg4AILIzKnT3g466kzYbRqE52I/qYrq5gHfUFEw6QIOkCn6LWq
76gliVjGmGHvFsDaQq+8XxRB38M734+H9xXQK81K1GiSuWbVNeu/Tzv7FEg52gW3LOfS+QBnRgTz
timQ/Pa8DnGTR8S5yAY8BcBg/8bW8lbFGSiE/7UirdpoZsNa4ktOl3k1NCD0vs3JlPCRYpYohjUL
cV4PJTSmh5XkqgRKd1/fR4VHFVoQ/t0oc6m4sttPdV+kw8/MmIGoXan74P6b/wqEpm7pml1bbZ4K
eV/wo0lqIj/4xzO20rwufOycSNFDMKpcaG+lUuBvTi0lwsNdIsnikJDiGiqABpOXSJ2IuS4CkA7M
pvrO9WfAg7Ti69YpBdR/cmSTg01lIalPXOM1W8Hk4Jo5osBIWwGobaKT6/uxTPd8GSLAYQTblYtI
Z7eHOcVDgk5VZaRWsl9oPvDz9vAcnBodOBbgnAbL9lCU9i0BDvphq0Y91raihg3LEX63IPOcwFkp
VbxW/Up07aFYGZsQmHqOudpV8ca+sBGt1ax86aGCSGrNwIMy2Zx7/hnFs9f/nL2qgsHfQejlw8y8
1lCeEBT+o6iENVBDYdWD6eHTo7Tdu1Y/U2guMC07c1QbNPqQNaWaed7qtTg1ze1QKgyvv4TUpETM
K+l0+SbsJuuUlEdKG5ra6+5UlH1pfxUxgtCKavgxeemmo5iUoeL/rEQaZAJ/xQZHpnmuNNZ1LvgB
TovUROJX45Cn3dakHMLgIEoIQqa5oElTpa5vLj74UfLhxfUHXF+sRtj4QST0NfMwrOtn66sip15o
yXWipQUeZR5WPqZGuYV7PziAzaL+AB4J0UIqrpdS6J5fMnf5DsYNCnz9My30OLsE7AKT8g03epOM
FlCfFQcPGdisSeEajVWdSfAR1r8S0Nu2MclGbGe/mMAr0gARPNfkZL7Yy/L70oiabywJVF20y9Lz
d7pS2X+FPeJW9BtO9qoqLt+/5nRoFzVhkuf2CUkWvdhsS6FX7vMiFeWNIoBdukBstjohSkNvFUGU
zSO/YsOGgbQIvZ08Y+dqLIx5GWD7AGTz4dJL6j2sk7SU21oQCX9SSLp6TqYitKvPEd/7RF/g+ijs
FDcShPpNdsBvlEvOXVnYdC4Wk6BNRJpI8+oFMewE3/ZgU3SncLFVEWFks+hzg3Ok8SqW0VmN/dhi
4k75fCW+qOnqzQ26YSy5ECkiXcVYkVH/OiHJp303f5lQcAEZt2mqBccd9cpzCUlBtbicl9FNTl90
BV3GRNcjhOChK38nSmxSWqvpqNxxTCqXJALjvyErwY3/fsYO7CVsvYfqiysL00nnt1cjGUnsUgjT
iFUVD+Sbhokw86dsemCMw4qAES5pJ2amQ689DDop3OQbyYzkTYHezxin8QbR09/do3u9rrk9IosE
mN7Tn3ZXgGgXrfpUxY4hCULnP5WI3TOqUJP8ixJQ+jR01ME3fJg38R/um5F1aLXq6UdRJ0+/BS5q
NDpgoyBMHQ8Lw/q/kY7HJPfkIr3FCgBQPWqF1cYxo+ZZRp7+VSQKnX1qdNUKKg6CPwvDx7xWhNsm
eLAV6fyVEkhvn4sn68+2XebN2JiPcfCIozR7BgpANySomfGH2npKoa/ImjvUpaublV5p2fiklTWS
klCNSBeZzIW6JVVIhA6KYy/vCResKBrKHZcPe7isNDmZQPT+EtTJ5KOeWSSmlSUT9VmYCv8en1Yo
XEpt76ZIinbK6cFbeJVP+HoZmIUnnjyo1soegb4/+K1LV/gU/e5OdIAPaNxw8KEzDKxIhjZX3jo5
ospbEn+u4la5BfPtzmFn01gDslwarOT1etA+XlHHBSxAsTCaOMavSr3CE6VGtzBfRemXtfTXcPQh
EEMADG9two9F0nlZj2q8jL8QEm+NEWWojtJQ+lJO5GnMkkvlObVwyyhAYmnEEy4YwFJ+0tFn6u2f
hBefOOludktCZ980OyLkgdEKNc0Vo3bxymatykAp5Rtm1s5JhSWQqYBYBF6UuMdBeWF4SA2yqO0k
s4MagHUybswi1SRoudcYFsfYDccI5R0vK2Ozj1T0WbkS5NY3PY/DthTLP0mchlDGHajFsB1WhYol
X0+N1EmHVob+JXNoeqEP5P9jR0qHFTFOiZuSSEq+UkQfzvzb0YphIjVvplYWiJfyDAeUqgX0kGku
472t9E9916AYxl4elUbcQ1Wkt01/p9rSUFDTn3iLeYCQigYtoI5w1joRDeLOwMckzEFwtW1pn7Hx
IfqHdfO5vRPVvHlccIXenlaZJr3+WITDFWh5acTz0fSDzejpZsc/LDhkigI5rqNv9pOAsaTeP0YL
Ku/8ep70Tnf3Wps/EEZ2EoJfsGRrjjluNfdWaHaenWTQ8PoZ+J3PSynkwt/G0LiHzQl/QqoLiX4w
J57NxxhAFUErqP9rQ2CldJFZUR134X9NiW0VnIR5RTxVOJeDQE7nzd5PE+rWnTS5EMyDl3Sp3Ygn
7J0kXOvuC7zv+uWZ/Pe0f6GWtgVWyPJYz6Te5OgfgPOMpP22+C3tt2Uf0X6vEWxx4NDGaiDfHBxG
F3bS0zxPVE6xqOrm+eqj9pfcz7CrwZWI54dOsfLNMVZLPjAZAk9MbcIe1D4kfAUwi6JEpfw3LgqZ
HCckgrfwowdW/3889+7EirnTFD6JKAaYTk0BL2h9nSbRSvZbMv56tUm69iZrc1/nGAlayarBvJKO
YYSiVC++YKelGf2cnze/zaNYFWy4JsaNFpwGQkofEoViFsUstElUhXJJut4DnF/mRu5sqECVrE2h
Es0MgwlYP8l5dCFI9ap/xvlkSh8GdYWxVVFW5PXSgW+bKSE53fbys7qD/65JWXWJrKDqkw8yZ1mn
X+eQT+Bf8Oiky6FT+DU80yya57rjKXKNpv97Vkwj6yJ5gYm3dozMWV4V0lZv8tb3R9rUutcz8E2M
3D1kkYrwPwQFa+HiBkvF2kClZUV6+ehhYXiiUJgdK+9hMql/YAwVjjCyGANkMh+x0thfFPShCyu2
kpEsNHzCG2bP8EuHAV2gn06oczbTgdopZbWw/5R7XkEUyrZ2ZKXM2hruSgU/OMaYdF6MfcQsSY1G
0hDEw3V5gId7Ijur4gaLDiPX+4UsPi0EbAKEYL1cTOpku2l71T+MDY98BGOX2kZJx12Wk6/wSHK+
XY4OJ/skLG6I7mkDDWALxFSVUUXS8rpOq1bveFZZ3uO6kX/ZIAfWvXiaHhaAyvftMIapXTbsAK6X
vrOTAWuFFdWYeOoi4hZHEFL3JKbpLD3XLzfAmBnHO1L+b9d25dgmpRK1Cnp1Qzg6u+MYlxe0l5SI
upDPXeOQG6ugmIKIybHi9/uzogYi1igiWcpBQ94KIKJ+3BEW1Py2sORmBmrMHkav7ioqWGRlYDMr
Oubo+QCeQfQ7jO8DdN44hFBoHcXko2oZ42khKoRWOEdytIQ5MmFruxfSqHHIwvs5ALra0uFI2p8V
GlzliC6ZUSX1ky2hGdJ4Ryg8rc9H8mVg2G89eDkvH3y0ChwMeAYcGhGU7UuFLT+4XEL+qIHTPlj7
95hY1lSeXSh4v1eTM4f3VsMV0Kv/lFk/KhBE2GlpGhIP4/3IL9lbAeMBwNuucqOQlpQln74Onbs9
SI7SruUg5gJ4uDdbChJliMDI2MAn3ygY6aD10NIs95plNwC6D1iJfIogvSG/GHG3xGMqnow0kwh+
E2WpVLhjt9QLGWV5DVap9Pumh27YpZvwl86n8LsofyfMUmuUdGQLdU+/VxxI2ykDuxwIWHJOFCfM
ILp4GXVPE6ad3i2bO9j8sKf8ujH3KlRwMZqsi1RPf4GCvVMJ2B0NgX0gFIiSAF2lj6D/MeIzUKLC
UMZ2j/E+vuFqohQLmcLctLefqkY1vzmB/7G3cD0k1oPTDR8g/CUrhobP8Ad118mkvdbjgSvbAybR
pKH6M0s9tsTsHz+xa5fu1A/Fb1WuFCsPJeRdXTW9alY/Jd/0EVV96fsNgeVCWKAERnj+iN0QsasH
klW8yGHOKfQtdGNvstbg36zozMamE/IMW1MakpEjDAA94JMq4nA646waIpdfzGELalXPMr7w113y
l2r6yFtjXvYTXYFaJWDSDq/OvddIJ5HBHo8AaSpkxfYvStN5ySbEIIo4DKu5ec9MNYf/w9zaNJXO
5QCvDQJaBhQZC1kac0vi4+PSsx4u+TX6JOV+8fMVTPGQ4S8Ekbu/udB13TZg4JUSvDhbtmmdcNqy
haxWMozdi8EbGkY/xY8Pgk6nCMaL+j/PnSyTIf8OcKJUg+zs5rsStv9XlUwL6q+ZnnhkTSQ3Jlwy
ClCn+jZiXdBJ0as4oL2XluMZjTU1gekVB9iF7HALKp8VjJBpo+GfXwkgvwsKZwUTm4RtypS4qy6a
IAQEqP7REGKPqXep49O9bJVE3k5+MfXWRzKUJOVzVmsbNRUFchwrJcFwLyCxK5DIryaEXwFnfrpI
kO8aMJE4bmSTlLVSrlyO0EfbfR/6SewKVMcLbew80WXGfFESy/EolkrlUWfKkqsu8ukJ5DtYpcxJ
eM2i4mJ3ZA706eEf9HWZGWzAS7773UYI487pnSaGh0SphRxjOTF4SBNY74nzWKK3QwZLWPngjPmY
Xm0VshHHJW+qsF3Gd1g5p+l5p8I2UzefzZkHf9M9ZxyqlG4MxSPK/yKJzD7HQAZ9Kc3w2GbQr/nv
hzItHSKsZf1RtmjfT6qe8R4RJM9qoYmMn5cdjZpEmqPx3afZmIKLJFxubdrikY3p9flS8jCz1o00
NMZeLdU2j9wLihhCtDPfxWBcgZzTEFT9Hhoz/w07mXmWMSsrbRmMujdnvUFx5pYuQ3kvIEnrW1ZN
g7Ud2jAA6JkUa8Vhlo/KKSrAND2yyEUIIcgUSinjkMl2SftNyCQydz56hW/Q5Y948rjdcp7VI6y/
YWTpgrdS0cU7uWTPFo599Z5zYrvsPpDvr38AxR7PLmthRXEouhNHmnzvtgoujOmGhpoli/u0h0Bo
TM467TE3rMMmCi6e8gnS41qs+ZbfNvRlQ1J7VEsvA+Gv0M4QWILrZ/HWgCwTXN8mxtM1b+5aIGaI
hKqZmcgTiHRQFQIZqgQ3xfMcjqocE2CRhi2wUW0XVgVKGtCA92+RsDoBRj+mAnlLtT8131reP24G
a5qNx/htClf/dqNEhsk+1ZsMfzAR12jOyEMLs33KykYLJkJt6bVww0c90KPhd5jF1D/kMlAsE5QR
2tSc+7w5g/COEGTCriIUjDubHQm4fKoyWtRGFnr0GObEzFY+NPbKLgszuTDQmxIu30Lsjm5LnFHZ
qgPfDRu+g8IqiYfGj97XWOb75Z8QfHSgzmRLJqb9avjHgEpIHXxlT1J7WgIwMaJT4LIgUfzoZc5r
RfaoZ56WJtRF2u6H43JGvY+Uev6e+2CPm7xQCRbvyB1Z0g16T4z8xOAkeraWf/3lzfPE2km0a3eV
p3UR6apr3oDWHeH4SMkl5kgkEV2rGGQ+T8gaBHPZMoN+vBhq6TfLWSisEwqfHsTHTlwy9MKs8uXC
GfQGJpHUdK9pMefP/YmQujrCxruntNlBaeHd4wduR2kuDDd46hRXbxYSdC89vssV5u+x+1IyvyRG
hfR6DQECRXpe09zfe1kRO9TgQG6fa11xUGbK6UB9uOTX/wYmNU9G+f/NJGiVUvz14QJiR2j2xVHL
jRt052BdtSOB+gqz2zqk1hqBA9lmXxyCcPLidpiaPCbSXK/grV9rI5NIsVgwk5MAiXkMCveFW7bI
BbJ/kTxgTn4ErU2qgHO3solHXUSVCNwwFJxZbGmAC6zKCSArjr5YL0pQEap/Jar6xpTGRM0osSrt
qwHR/JeS4Ip9bxuK8toy88V5WTCeWlw17d9VsSLHsvDFkZGS8h7OSTT+LS32g9qvzbnYla278viZ
M4+7q0sSJBqhjy9WUwee0pIRasT6cLjt8y5y+CRQMod/wgnGkH7ULGsseU8Kl2D1U00uDADGyTNk
czRYSMlwLQuEzpUMcudc2OewkcQ1U+FPp5TK7ZZsfKF4vGoCe4yFZcjsQQTYh2R1IFFhSSVQ77J7
zfPjr1Y12J0cC3ukysb1/pXbASATx56YnOXTkeKpFSxDBo2lY8stato2/K0f2VjevDBKYt2DOagH
DQuBJhgC+bgEOqaN4gKhXvNR22y1wAr+m9F9WiRctlkbeCTf/9wMriLj/O5YC2HgYultz5oDn+Vm
jp0mQ6rpKr32uCu7Kau7yiI26+NVRy5HmO8MQSFVyC2mv8Dq3AUxTv0AJxkSlsE3GLmjVz897dWq
xgialmYROc2Fzj/un1QmEtjZoCMp1QnYraTRZe33qB0eZoZ4Sr+14NN0UynSlTRn0CA6svZtqflT
RPn2M6O4y4wY96mrm0yyz8RjIkjyj59hy8WKwP79kQ1LXSIbjJXdPiccsXvb9T7KZbY4AtKTqrcw
UaCqlJ1/9Z9R5C1oL+2BFUhRBBhp2Gh9BCv5FCOL5XByipOaRncQz3vnmdS4JOCCG1MxKZkiKK3t
jChBYLTfysJUHd7PtG4q4EX+6OwwdmqX8I01DtuNZ1gHgbIOvZ7trW4v6ErdpOTZuy7pOQ0dcyQ/
Gp85nZxxiBwIgA9KAc901qghow/iqPUna+DLSiOHQs7WUkCgHfYQWg2IIemlUnKaV/Fu5LKC9yX+
nieJqs7cfD5hFNhTMtxhz2w6cY/d75Vm2U+OTfdazvzB7Yr5GV7m545g20ltkY64Qq899BqsuxF1
AL3hOJqeysWXYPlWrqeaaQxa4WlsifIoLJcuxZenJaqBX/s3ifR5cEvJEUuto+P3aOnKVPYEWrVM
ab2SFlRbwSpdU3F8vAGyQdYWlYgtjlbi+12LHPi/+esQ9Cx/WEC6lbldBuBG+n0jSe85UhtzzcyI
y68ZAWhd92fWMwBDf02KiBZGz0yc3rhKFJlYQW3px7L4IqVM+fuwO6Ydc+CkBn7Kx3DmRRPMw6Sz
1MofRDhiU7xaZjWvd/rY35w3FxoEphYCCcenrJ+8EF0XVJc2mvX1AmJcPN8fKeYsOsyXKJXVbqUK
lY5lS7A5UdvfQcn3ec2Jpzafr8dvsciFhreUIqL/Q3PpwO/Sic/CAObZ3S/7KBG+9Uqyh5NQv42u
1HMq0yt7eNzQx6CJc4LY3DcnKcuH6JhXnD70j2NpnWqziN/BcUvHokHFbECWaj7opOrjGZ/PYas9
bChwN03SNJRd73mGvEMtJqWQhGxE/O6KjsvDJa6n7v45xOG4vFFhwiy08HVdPzgfY/a3dIso/App
/FW36tOQNUYwVBzXQze8wn3bWVOGrhr4qgPjfn5s8voMMBswjXP1ZoRYiHZ//1xa4/hzkcGTKLUx
+0OUk2PiNNafuEs0Xg23S5jjtaVaxMbyBn7pigFuBLQeymvR5gjo1lCa1FM8pBVf9BbOFaIxZecj
0b3fjAJuGKy8ABTeH/LYeIuYNqkEQocJML2Q1EZrJasd4O7pjhMChzvOsmObIaQU3deX2+oSASS+
/kbqcdlBzk+IR1JNcR/sQctjrY0ykxbd9sjCSTtAuf2smgEV8D5q5rSt//pLCszZGvlBPE3p1it+
Mj1MiMLAd6CqioxN7wtFj+L8FwXK47Hz/Cwwzidj0ZrjB+0l40UY0YeRzTTGAH2Nw8IakfucOjDh
BoH31TN3mgWCzv6gEMLgF9A9EcegE1uLiGetL4g6/iRq6mDfd6u/TUyNvh6sgGf/8JD0XjBlgHgM
FA+g3LzB7TAqFPoz3ep44UZr/fGi6o/mOrPlGgFWOfPS95JOTylXlQwKt/4XBt2U4Mw9+jhwMazS
5s7wy4FtAzA3nhGK27ODxS5MLqgextSn2Tm722fKrXEzMLFMBZ5+UbWSuGARmBL8rCrej7l4jRYn
3f32GEmIpfORmit8tEtELBIyC4yt25MpHV+ozZTtzpHNbC6MtVzoLLmb2j3ejQIJvxQwErpSAgDD
nGN3jni1FZq4GgVDGOCrczWpYjIADXciNr5hxY4S8d1v/KdYhMDiUw2Lcq840rfq8NH0QfX+r+es
YCuEyqFM9WNX+sl3O7R5xc87W9pVFHW8OHSSMnw9/okHxR/HxhAa2CMiQIkCV8s0/dscXD/M/lnF
ZN5PH6AkqyMPplYhEE/FAZiQfVOAYiaW7N4Sw8QmousZUWaKiWRH9q3kTd4tIET/Z9kEI9YPEwrN
RW1RcYHd1a/8g3qqR4/wz4gcelvTD/eVLfRsa/45V/iXrzTU1P4n4YhKWgSOqQyhBquUyKi9XFkV
r7qpoIp1vv6UZVRs+YFO7Cd4E/YdhdAnnu7zsl8cyOLr4Vv0yV37jXLD15lwvePDWsEkwvA4BDBl
x7mTJFjjAov14nIhEi+UB2sIyOj6vIN3Eh3aEmkoI5E1k9UnmKNtII0ZPpniXkBeUI5rL6v9KLeQ
uPTpqpNMk5H4no1y3KDtDIiC2OZPOjsPwiAsrq5DfSVeGog4hz4xT8upXy/d/50amzF+E7mQp0r7
RKF/c23XLWcvtXj8SBYG1vXMgrEp8su6co9vpQdz9mchPAH2S+wDZ+DgcLS8jrJi8TaWow4CfpG6
/SHk1K5xo3Jsaq3gQrPZXT9y7iyUXGpzJZCiAiF2i7ygPnp0kVg30B+FaJC7aHHhPMSnWZtLmI87
+zcM3aavOEh+xbbST0j+W9Ts1BbmLC6tvwTuovNkEsU5BkcbW9fq/lSTUCBPHQjny6e9M21W+z+n
T6RAaj8iT1S9p0LkXT/d1E9PSV3GVyVmZCy5u2sNYorKIHcjPiovER3nC/y7iuuoA0pb9Y2/QF/O
yD8TiLzVvYF81V8XGXQEBHNseOs/werNiTFAgvqpDJdjyyLHQHduREcBPrLVJX/ToIIsYh1xsz7H
YEpK9dWdjJrvTyhbXIQyolnrKvCFp84Pt9NxIDpzk+GiBzQPCpPFRQcU/74cAjsmVBjAAnziwRBq
Jkm4rQv8Hj0/rB+pdMOcd7cUikQQquBj1ftJeGSfR58YNwruExuAOtJ15Kv8tWCwP8zZWpx8ve8H
8gt9iSpGaVbOumNXte8FQsiJbax3YGY660H3SjuDy78dkgwNtg4sye4jlAoLLHiWgfD/hS22BeET
3yNRPsaTmmldzBoc9in26PC2KByL8nAVu/p1GXuiP6d7aRdJpXxkNnG65gDMrbkj4ZCj7qTnp/aU
NSJd1qJef1TvIkm0llLrhoHXm5580tBK7f+cmm2AO4zG2aAPR8ZK64XDbneBwZQzRQbTeeo+bu3+
7tgAygsp/sKs4ri3KvjnW+1wRITCDAp+dRqUJLeMZXwhm5S7rm9CZd8D2fl2jnBQq1UywUN/GYKE
OCWsmc09vdYM38Wr3Xa8k+loK9wV6ymO0hss6cwgQUB5hErU+pYJYn1tLEdlE51pI2ZExqsBK4RY
CAzADdTPc3MXKwHeN7qZewwH0bVIj2drhQ8Wd0lLxdwINndRuiXPkm1L0NoJVLqUvux7w5a68m5Y
iUtxoPqGXOviIiZ2dkdxCgCUpm5wx458XQr1Fxpzw44QkhhMtlC2GB5lCqSUAx8vN/8lk4EDG7BT
O9Bikh4LZ5AzjLvMM0yJHNHMtv1LzistwfqVmqSrfMJLMGOvNTfRNqCPDwzacCm7txBJA3ocIqeF
gDBOnHNImGJzwJIE00T04zNNtvWwYheZa011aIHZXPVfhyeGDz/iELTkoasKqPvIXpJNsVau93Ww
E3U1zXQovjNc7yl7cp12l3p3MMI8orToEy904yn2/GOdmlM++frc0gVu5REcJ0vHk/RNwwsNcgsp
X/O/mS2pnyjhKBbpkU8GUZIQZ/5NgBFoB43SmhBpFB7vNuc0WJDdVwWYXmHC0eukRrIZ3Qmcrly/
ByWDQq3hP9YaJtHRlJ9pMnBIe3Kwf3hHGC1m5IDGJjmAM1QpwsJ3JtzAysihgLxjyZRModCiqpyE
PkWfi3vQ8mLskiwCQHIlmgRdYTgfePQaoZBlS9H2T/jwxnoSL/eAgiAp9bRzVSkAjxfcLsddKpmk
tEOzGX8+nbzb08uzJCbI1vtVuQ8WV8i4PujsQO0Qs15opGLt+pekPfoBQsy613Dvv6WdEHTtV8wM
XQKj8pzDuYUPLs+sBBC2xuxRyU3jM4tDXmGB1GCWRk/Ieyx1WNSmx0DsVhclj18accebPwJP7QLt
cPcrB1qy4Vab2bjIFCcpBLVFbLmmyaji3YVLu9cK3cW9YGWpYK/eTgRRXn7WULTD5rXJFd2IjRNs
fb/0863t/GTzGLDXkwEZkTojCSM+w82qMz9Y+IbPxl2yBdC+IrDLJSgFU7y2IGTT4Pkt/MHPzlta
RV+WcVsCt/WvqELPtcLVjIVVz/qGLOUMuPIni9I/rilDlKUS/PiOis1b2PTtR8E5KwnFPAffuyEY
+Kzc2w0EKKQxkZsSSEb//c0feliOQfpAFC6DOJJjvBe8CopFl80ux1TullECw0eIuDY6cWamsDUd
zK5uY5uSKJsKK3sRAtBKmXWNOJ/0kDE7yO0yJlKz3Cxoif03eB6NwUm4o3Ro+PyikmYG2gg1EROi
vkpb5I+mtUR+K9LjqpBjdSwfWMKa4KRL44YKv1xYjfP8larcw8f5wZH+cjE34eMU3NqLFjcOBQhH
m55Ibj4+kU3Op/fKPEiNjUD9i0Ur3YB9mg7BGJdvuxvXAgmeyjvwXr7UiHxEJd40rXIuhMdq9swy
Baf2WKJzsg06Ut/L5umeJJNoUnls2Frw+PRQb4MCk/kXLIQrFYeug2+GV/m2B4HeimFEZMaJJDWg
fWeeYCz/7l3FX5eldcfi7QUu/vB4/L3AqyHeJHvz1aqlcJX47TB9AVEvg473prWmcbsUFOQuoSPL
lbp7bdC0LJ10sW/WkQugdeZ1YZHopLdrzzHpyHUkHaPefPKPP9XLlLJJJ9Enm9RDG8j5W647Nv79
MXASTPdA/yv98qwb/bxecCukkZ2EpBynCfOm5GR/G4FFylkRf6r4jrtAOCIhPThJaY78OEriCoPI
KJaJCpTgT0t9XXu7+8kL/FoCOd120cmKSJDRTJVOutUqcE9jDQqQySXc0Ycs1rUhVawcxRLHh4dM
c0CE4nd9vHAAaK16WFszMqz4l/FFpyhHFU2P34Dj8k8J3w6tkgnLKB8gNkQZfUL0Ui8dGBRiejrw
FtcyPr7TUMeRGqK7VgX2tqGPLY+FJ1kLpjzBiciyoYzM4Veh1AJDz3k0Bj2MZhCNJ4Sy9tvuV7ux
UtudNqdn0Qzm9f1YwEKn/PCZlzMt7vqlusKXww3INWeaZkJot/ZVTYcQwkfUg81U4poCQQzE5fbH
hj5bZTmcg3rmAecnggD2ygBgjNrAnCy5L+0YalgA4EAjRvsSQrVzNl80BffXlcio7OzOaFKNVZut
SDy9ltx9HP/pAmiE2E3poaQX+sL47sYPRjja93xMHkVLSS3IlcDOEOjbKglhW85jBXgMG6uDaiPb
7KPxCykFsrvTDPq7XsP7QrS9FfxEbzH5biedkXgFqrfDBzcHlKwZ7ryQl2zAzitflAAy97ddLLMW
M6Dwp1sleC6v6c7q+0sTUhx2sJgOsw6XCeDnntd3O+tf8I6H1LJI5hapnzRk6tVTzyzMpA6Xjbja
noGvqLXu5Cn86G8eQ07rIOh4Dv3p3eUB+mrh8PavlxBk+LxLZpptPbh4KUCZYy7P4AI4EG7i2B1Y
jhtg2nskk4IxrnZz/WiQ2Yyyc1jWa3D0Zff9HnYIrHjImq/YnhB9uzggte2jyZ9nw7YoTiReYXeS
aZcr8HEne4KrEhyrJmdTHjxFQiuY+D6EopN43Lpca6/4+TM6J0Bl6rx1uXZTNG8alZh2Wwg9Tf27
/oQNUd2qfdli6UHz4w4I6dIt3nMNOrMFZR1ZGkJoKzaJIMmM7JbljnLbUewKZM8fxemy55s1SDbH
TfZ9a/mpz/NDWTVBX+l203ISl64NEsdiVRuodh6djQTKrOfy55l6bUS2J54fOlNKqAetoG3NVNjc
3jtDeFHtWaGnaNF8Cfxt7gWnTtuOqgN8+FW803xvt+he8Sa9XbgQB1M4Rr6dwFlLvedrvULRFdFH
8RU3arfrWtpo0oU0mSqnlah+ep4og0ffc6aRlIaKxW3Iv2J/wrbZMmrMsYTLEb3Zd5xy98FE+8MQ
DL45KpRtsrcHe64dff7cDUqWaM0BEqkWNgzXAmFhY2ssdI5tvKpRHtWIyElu9j05lbJRY5HKvaQU
wJrMUOninesSeGrfXplIQu91gKC2etoAh2u1vwJ60bY1d/qLyHsB6CTvqS6/TFWnO3iRIB4618Kp
7wI1OUunxD2h5bb7GXTBnBgkLJIQAVkC+BveY48SVYrIun0MVuMUJ1XcEzxAdLF9scDA9FLhIWi8
/CZoKTdOsASf0RoLMJjXyVkGO4LVBXAYjPZ2pjKgtF4hgESR+3DT/2X0OnB6RZS5VtMwsZuXCRep
H16jImrtMr5uceqYxhQhtc0VLv/tsn4akR5CzKd2XU8cDW6poEKbTLzvmGHeEciXRNLWYQjWm/cY
Y4InI1ap+TXQe04zsBSe3hJlPVun19kAzimsgyviuBnW9pJIaNv7jsOiqCUcAilVT1epGM2nK94i
recBqrJCUeZW4Jxu238XDPHVwpBVZde+MYxiN+aD26cs8xRWTX5Y3jAun1T1+7xoPyt9CAY6OdMQ
JWLuhoFd2QoWn6dWWOIAQjG0LsyIY0fsflNlQH3Wqn9F2v6EAqLkMiMSXV+e/Hto53n0qKAIdKtc
aNwdTRvehb8nEtqkjT1C9VK18OzcYuk40xbBzukR5gqW/eIaoM876XbQwtR4Nn0yUoituyxFrk0U
qLhp0CyxV3Coz+Oe5PmPYQauQLfgglwsy6TZ4wpur0luFKO1ZkdkvsJ90esPRw6lDiatJ2bHQv7g
v2n6g2bX0mrSG4EfNl/bIM+6mQqJd0Mq8JcCPneRuejW6GM7gmRoaGOfdJjPtwYFQlt5wpEfxCjO
fVHe2JIWNsHwZNmQCbMcxHDhNhLgSIQBltPmf9AKu1fMDFpBQlNSvlZY7NlyOmNBmd3JjbrYsc+8
VZ1ZQuB+XOrFmo/7g2fPLtMY9f+BmGZSnA/kwmCGbuXYpix9M96W8ADtZeo1LVDcMnz//2cYkg7H
olhq5YKu2wr4fFaTCGZLCn9CUAEEchbNQIZT7Y5AyaWIUOJZIcAJy7L2tSWbf9g0av+F2YwbJKec
bu1JIPc/Fxh2Ts006bhWgRC99jb0KFU4oHlet5EB07inOvWpYzsIrF2i+pZPZzR/xGIzVsMsGuPG
mm8A6HwTKhmzfBavrI/IFXVjVAfh+5ooj/sHmOjXJWl4+nRTRIcGNSmkr2CJqMJHsApAnEuhPxeu
im9PO+JM6Dpu4wRgWb/BugLPD0X0th8qjXjHmcNdiMB7RdRsO0qcXig+Vu39CiDz8uUCeaWYOv5z
WZqAcpIJmL4Pn+MV7JCye3JWcMLUroy/MRbfJrjdnNtaxivkUjWrOoPL6v+hooARPSLi3xkx7lUc
q4YL42Bhhz0jnkUAciwG54n5XuatFJxEy+IgOqdfwho+QGM5ez08hv/JKLL47kp3miGQvBO6HeS0
cq2+OJa1Dqd1bR3KGgnNRJ3nPmzXkIbkPoqOGUzp/nnSyXZibbb8lz0yGuZHhNTigh4Y6s4jTjTG
GSDEFQt4zDnBfDIOJfFi1S3Y/Opqqe6wtOPXDEJI0ODKBrNxSLmrKu69LvmlvnhGY1Sb25XmTVOm
Ko1+wb1FnOqrJKYQQcMWpfX2grbXtWVMVtMvy14a4V3NRpTylnKq5gr+oWU4VQuQpMclMbqPruBt
t39rX+S0KD+7qZovNe8cGS3butevChdwpZiq1OG0aEaLC+K3crdAV1uGWCNI1mWO3RUH8eKxtHDj
UHJh8or6WEmAXQ0liqCtpb3ix8u4ZD0ft3uCs2uWlUljWJvN/TYpigqvZ6yTKm7VSSIzzrTrLWZu
NgeZeI9di426r3ZEThkuHBnNY8k7BgDFkpo25GG+iFL95OBwTbPLws/9f4gXGp6odXIM8LfaVPGV
P58O42ReXZGPa0zMcJ5COXO+Zx7C26bzSPaNsntb3D9MDEtkOMIP7BewRz2Fhkfj/sPB8NE2AeN8
exgjKjIXq4iM1jSSWLQS2WB9ymkrEqC2j32MHvVVicHQff2eXTRBKmcSG7rCgR6lY8fW4NUOwew5
0CfEt+9+9I77gs5BDuf3RXKMjaQp+FuLI+k/Eo4my9m8VYqLw4mev9WQMLthFxUPE6BAXQZ9EfL3
jAPWZMvBe8OIJpQqNkfucGGVR2Sy4aMJZm1/X5T4GhI5ur4/hbcTh8vIw/aAh6OKrRtv+2EEaD52
SX5IE4UxGPD+AT1BP/UD1pOapPKmm0MJkxtDuRJIxcMUtHRS7AE2rka7iI3pBjKAS+OU+tGYaWh6
g8x39fDkXEbKw43wLZsdcr2ZMse4EKbBhoMOIbw7TJFgXr88FlKwbTC2EgUPT+fBTPyCgezlQbj7
7KGxuzEULHyKV8zx+NO8R7ul9Nm980y5OF5/L9ZigUVWc6o+TKpiwL00jFHoUnbxq3naDkmrbrMa
QStcNVElOOKajJe/LJ5inxHIcjGcuATn2XSZwjejlwRAD8OgNOV+eq55DnmRS3tlQC1VkMpmrtsT
MQ0P2fUlGo5VQJZQF2QNDqj24NRj/hKsOIcZbFvNTkr7bx1MHeMUeC37BwNxnPFX7I+MIajFevXt
+TpUtF/yKUyD7lCvn7ogBawQHff9Q82MpWE7b32dvG2dBp5HaeiXTr0D9ciR466rtgbBNaHi+C68
DkfD1Mj6Bv5QWIPllKH6pSfGe9HRQ5HcGUjjsUAJKoBVkoPJziEliixj2Gl7+p9zBTPMU2PBavBo
udi458fMHIPNrucxyDinjJlbU+HQEMYfM2Us92RGVlRUw0HUKkRnR0l1+UasFe0Vbx/XpsWSdoBy
sx8x1J6tUY70ucrSeTUO2EPTxIObpHZBKX33DfnaZe04b6eGjpZlBpG7Pu86gjhIrdc7ksG8DRre
2hhQm3AaNPfmJvRv0NnUIpQvhhzayBIUZ+ttdDAe3sN0IK69jD2SrcHwTxPn/tWz53jqConR6XyB
UJBv4NVApNq6oAHVUieHI0OTOOsquBaRCHsZ85MyivdTiKys913K9Y0UyngROt468x8yhIIFZa+c
sOInfJy7Q6HTF54Lzu9Rk+YBhvs5yPEctofEQjgq6OXfseKoTO+5GcCyhagJt21fYftnZ1D/t/GK
1gozENf4LdXIol0JrFXt4r4G8gdtm0xTfQq/ajgjUTkUMf9A+QBYT0f/spxOlJXYsnFit9ObBvCk
aEsNUFxKs++bfXDXQQ0rXicCP2kaFLb4g6imHzioGlc7ofa2/E53P24lKZRzg/5cybuCQrMOqg6o
dUk63AUWtKcRzjS8RKo2v6FeySxEl9IbV+WBlVRJGzT0mH1PN8c3MwXwHpIbWpDPZHMeRyTc77Qy
C5aeK0hwi9Mqb9jFpA4say87p63Bn3AyY5utalmKXho+E8aRjckGNZ1IzoKB9aRTUQ/uztxsPTZL
t0Rr8KyxRz3EX8RejUNKTCQp/gu/4V3qrDbFuiQhgk/BoXHavBBofNo5k1NJdtHABkqS89bd7Ig+
88jlt9YsIqnh5mNiU1Sd6f2Vu+WnAy6SObhcTberHI14WDRwgMZGG02OEoTtHdAJBFA+E3jcRAy+
2j+gtbpoIM4GKgIkuM2gBt5aJTftIy5WDewXt2BSPqKBgXimN1i5RipN7aUy5lJscZDWdqIzdm7B
fWhl3zrIfg7VAScNTq9jpTwWOy5DvG+J8YT/46QfC9JecnI3ykHNygnyPq0bJgdfawg8cr6XMSKn
MJX/YGQTsJug77ifuMlA/7wgr5cl7HsttItHj3l4RklJLoBa9S9Ckke/GQeBd9Mohqb9bp+Yka50
KvYTEtPXg9cdMk5E6DHiquLcG123k/nOcGE9g/Fgsw0EKDs2fI89aVs7BuZcE1M5X8Anv4KUI7MQ
Mv2zEvitTT8pjUZQVcTJjo4VZqqPjRUTXzUADyfnrjDivbuSmTTB6rtd0DUsHHHf9z3qRGcMvL9U
NYeyYj/9tLTXlXTviCQVn9uXhYV1EKITVu8eXghY4tADRfzvlxrIX4HZRtEvxFp+2J69kJkWScQz
9TZIrvK1aCi6l9FZKhlYZMYuXEnuKVvjfZItUPky0UcCLAxZTVtjT8jGOzPFMltNIseRaC/03UAj
mhaM86w38EbXS0IcjvAjeXenTSIe+NOo5THLypUppVeVjHCLBmQ2UD37GKRbGtCk1s+EUR+x1Npn
sTWnspjNm59tGdxSURqccTEl2ljJ64y0V0CAjSUG8vr6lzePHGO8lE00PsrQqVj6h9gCIFaRpmFL
DdvpSs2VkA3WS4vz/ytbDiwSuVVg6JbrR2ZMkw2F27NagT1zk+CdaT6EWbn9FH4Wh3g/lPOq3Gib
tQBKIbNlFJtvmncOQa9zo1+mRM48QEjY5x+CyrCLoZTjl/kG2ej6G/+Hq41vBz7gROzGZje2CrJy
ikc7pM5VEcYOurk/Es43HK7Dg9jT0IzXTTtyMxldk6CZ2ArVRmR+f97HuR75R7bmIN4M6ZIHH55u
mTXqkhBk7xiOctVttKuAjQIGcIAFPbZoTKz5f5t5lFSjXJ8OZFGEJQ8vLxVO3w9YqbH19vSaiUJ3
EIMV9vTRVoC11b24dI5Y19Hfxz0EqFJ42jiVRBo+xh7xIYULhMp1CjrLu5aTJS5NMPPE4S63bZUI
ktGVC7H+Fj5Gulex/MAviUiBgwOp2gTkKbm3kw/fU3wiGoiXy9Mp7wYXFPBBkpefNY86Ci4UOkia
24Ft61IeGPiydf+JYxMGwK9Okc0IovLpKdHCVItYu+dak8aSOhA00skMviKFah8NrHpoVg/DWcdP
XDtszsyDXGpqBaBBQIMBl72wDEaBfnOGo/VGWti10q4NI8Sj0SAmdHEBCwP4Spr+sOGiiTGYUYxl
kwZ7E2esDPmSLJBpzBieXVRjpZuiKTcWbGc8nYOi/H+q3LCBZxnFllnQ4fxTYa5ERaRKyZsgcvKf
Sq5S+YlMHLuLYevvBBkXDUPCqvFtEGIW35fCY2Y6V7tAcE2BArRYKa8nu6IR/UZcw0aGUF4InTtG
8m3ITXyWy1nTkQxAUMolgnOWkDFe9X2kH9WNfhZWh8uWn6u/cFMHjmIQypRQZnCmOZRIYSX6Lxtj
hB0ZI1sJuOfxyDJtCPlxRtibhRIndz+RMsyk3MqF9U94O2xK5KLeeaCugBn/jUanE/67xP0rPeH8
mlZC30iD/bhFfca/dI3TxhVM0izR2rCY85EcUQ81rKuJZcBBvt1dH306YE7Bdud63stDrcMwx6r5
Dd6y4BaR6m1UgVFDLrKAhYVz9oCsHBft8QogNSCKhCVB4NaJfHpuXCsXUnTOB3e59sP9nGAL6PuH
s+fbHZPmrIDunitKBtCbPkEuDdKWzHqTHdCgRcm9AZ+Au9FifJ3iM3LV+Hiez5N9zujO1+4P+3zX
XcR+ANavhptp6Rla1PMhho6fKjpXWQLPMRFI/UyhGI4RxCXZflTf1ODoPfnvbEwblKwcPi+Eeddu
ROBK8EyxbwD1x4flwxqUOqzl4WUVWX0Gasklsi9gjb7/ZDk3kmWVNXpwmY4A1HtMHFtl2seK4rZd
OI26E5yEQYPaUIm/yUowGHKqUrGj7w0iEIZSCRaObJTl7zTFroShtij3jzZP1TKi8RFAscE1NIF2
I1uHkgHiX4VFzos8bJNatZM42R2hEjKsv+NwVhYtUWhgrMeu09VVqQr4lJxohtMa6PyBjz9JWrgK
H91WQVLbUylU6FX6x9p/0UwRfoq/QQNR/fnhrcFCBEJ/vT6ecdpCdGDa34Mg6+2bNYJeR9KxyiB4
pd8ELF6lWpFMsJyOmlM345CajTlfW3lFchYnguygTJU1vw6foy+YAktTY9AmFg8bx/hau0cXlZSx
d58WsT53sfdibk17njHoAhHP7BvE6njbq2bTvvSSOXsy+NSMx0n3m89e5cRde4ftLEK+Jh2Ai4ks
Abg3+8Rom81yf6P+coviP7JrVoGcXUUdYg2ki/hW5cW8Zhjccx6PClJ05jj3j9S4mPdp9UumyJ1F
Es1atr33hsMyFhxklT6xNqnx4JI4tU5Nk8cVqr1cxFOKmDJQ0qAtQCkAypT4SyGCDtQvjwvPMAGm
/xp7Fh5YbfZdQC8/rG2uNvaJv7nrs16FdCxnX56gwWEtsm3PX7wW96DkoabFEGSbXpl70ereIwsi
akdHtNXVDex8YCgineqFyrVLwDwHSblKn7SsNWJ0mjfdcz7UElzfA0Dkb0m4vQ4x8KhCZ9VJ0efh
HpAAE68oODOIwShNtPbU8tP90NAgEletxzG558naZ8YxU0qF+yQ/MFU/lC7LDrUyo79qJkDiRM/V
Z4hAGYKlIQxaLMw1svrZt26U1nHEbQN1g2hZXi0omgH2J70vH9hgbgxwXz0VBGwjH3e8465xz9ez
bw/lfVw3fLSExqRzM3pRTBoR4tjhKzpvsySyWNZSmyrKBkgb0zxVwnLAv4yOGdPSWJuMKAvp+Qgi
k8Gb2Rt5HEsMhyROskyUcJOWKOHMQP38HhBSVzXV1M3m3ay8zVi/NvfctX8UXwVYQ1jELo6iy5tr
P8YVVRJwgghL8AEGhuGAzbdrR2zgXcxxlrj1Xiw1fKZOCrZPNh2MzsmLBQ3sItXwVQck8hWoWmCY
2Rww9hNs05ZwCXuElq2Mwj2DEOM7A0TsaPwcY/ITctPcaDO7/pDyxMGjdI4bIm37g1cDD+rF+Lfw
FZ4yI+TcTTF0N6oH/12W5WmMv0XA59MgJCfaEl1nC1TScnXj1+tXk3eYHP7QppvzdnUbRfprPvXZ
V5GsRHAxQ6W/ENt2tFE+RIHKDUls1j2ZH5Hf+tkhY7hhYywbfzvYoRW2o8/r9pCZcmVPQ30/L8A+
5gCVa6tCNWwg20NfW716FbFBnGAZ60o1+W7udm0KtC9Wo9KfATh0m+yJOSSPbF2KJ00xJa1cJHEu
4meWT1MK+CNAGr42DmhpYjPmHBaPGCz5vRegc+dKKeN07FK3N0PX643CvPf3lelZVHTisGNQwVbP
nbPjwAle42c/JXUuqPcO+iF0g0g6MWWhRKh1TExRqAMR8l6Pmk4PW06H5wjCAwYWh48ELWbzIp2L
RVPK0+pRr11Jtm07ylG9/WXMsLlmfFqI6hXTLhdCG9/ywcMlDvmBvpAPGmKPYo6yAyeriQ+Ck/D5
OPxa7HjvriaskYIbdQr89Zs1Pw/LN+v9kknR1O1+1APGg3Uw0+roCnzArVqASemiMfrhxGjwtGMI
q98/i1Qt0FNHe4ie4Y/xVwt5fqc4mPKu7tKt+w1l7vsGGmBuw0RqO78LQFkQ6kQX7BGEbLjP2G12
cypfQhU6MJ3Qqf3bh4TuTHC0scUzpoOyiYoG3ojUzwIBIPiETAHY//WAzxgGZiDtLtRE8IDgnPRC
6Rs5uPzJ1ffn6NemWLcxUOtSBJfa1148Os60xlLTjyt3MPzDYCTIJnBnMBLvNaK6pQk9s97qEQWm
ZetJfteCeaaupbWiOFspI4lsBRRXRCPNXotVqYmxqdl+TBBjdKaACBMNYZQuUe5zYew4qASCcQYU
HL7UpUJWEkVhHGGeYjFtuAzx4wW37/VczWhJ94ho8vxYWPZpInkHJTJKSrVc0CUMI3rAD5zxQkmM
3FNNFrJOaRl/TniccigRsd/PVOsrGZOhSysFBfIXWo/wx8t5md8Xw41/jgVPAOUgJjr/Up1lZ0/o
CwZOj2BxljT7rd9CEoHssTfHBp7wlBRezHOi5jUCRajX0sk8k/K5476NS63JYEzdhF6IWQzb9o2R
zjTnbaTKryK7B4ZDc0K1T36ilR1tHXDuOK2tDhKMM5v2jzGYbENVfZQY+mOzQjmAYRaYKyHYvtsF
/Avpn25Z8EL3BjTJqpEaxrZI3H6L+bHL9mXIztag0XR7zzZEq6Bo65O7M0JkqjqGlObLR4/3H1B2
E/b6QXv72/Y3jpFMbQ321NMvM+SjFfvlofBaDAQRcDTyEBsSC4NlZ/bQmfcne/wMpqRcX2pxK0e+
qacuPr9djPAR8hMaRCvaMzWVSrjGdCOSOOlYamz9x35G/s6lsuIrLGrs49dXBap4wxh6wezcTp/I
lTHQO2bZhu5xQ4dxuXW5Yviy45MhTryskc2ILNIeT0BpyAfCDfrVkfjazzMrtuySglb95sSzBMZV
F1taMRKiuqXPJ6ZtYKepEzvOCN6+nSqjoFB/ru+owm0JBbro5Etq2YIu+1pgcSb+Qj+2e/+SzcgI
f18FrO9WklKBg3yE59IwGXjVbApHOuGA/M8ngsPaYpM+PvJeZeVOev1mOWt2zyAiurYxwV+LxPdP
4WobRvoRv/k/QAJJioO6hNh1yB2TtuwZARHBHVReFmSXg/9mv3GpMDPNqBVZDw/nGh+XB920008p
48exnthp8aThra1CnXJ/FmSZipo1LpJ/EtmDnuTqs2jSZ1/Zn70ydEFmCFNhyQLE5KTZRVekTg3i
jLo/yfI0uBPFERbd9ebpD6fJxy3vuMOAWuFR8RjkORkqXSsGDdYHP0ulW8ttRBj4RIKON8Ycvqoj
unGrari6FiAFAzHb6i+fvfrxLybVohcqzBXJvLyTkdavVViUoZL4IrId8hMrvHGqCiG0L7gfzoLJ
IB71bhUeUXoxV63bAZJOHQnVPvZZ8b0kUmZLCrgjpnRBbDIW4xSA1LzDJr/7gdeSLIJRNDJyBXnH
wO1pz0zIM51Qo6YoE/uhITRlboZLFv1INfGY7xkEdZgp1gabbR7qTLV8tRMDvYkIoC+mTcEilAoC
RLoSWDCmElbyzNHTCSpZYhxwP5zYEtGFp8VM9dwXWwleDeSWATbYbFToiOmEZnStkqPbgc8VdtLS
/Ku86XTgtpLvrVmEPLrijD1DgVGCHfmflkhxUujyaWF158tBFEXoUTkU3QJN4bqXT/FcJgesrGdF
4d0vosQwQ6Ulgg+e8PjhIdcxqDwelTR5IWv+Bjyn/wcTZGQQOVz5oFAk6Rc5Rehh59uz0mE1oaHF
PhJsKPIJOIjOOiEKjoVsZQbjt2jPoxy9TLesTWDgSVWW7v99xcIriH11/Tb/wrVYd8RCU6FBBh0Z
xfXF6Q55Klz4sqMpIf4xvgmP07/eo6QSOxqh4lXrGMzd+PL8vZ+PgtHQmgcwQM6Q6vT+/LT5mcax
nab/ItU3ujUKStQRK9h1JyiVOSMiff+2BVcQYu7rDkGxrpzqhfJbjPnOIRZmgQEbEJySgrFhn86f
3P1DnyZrO6VYd90umpWG46AGVksR+rNnbn2bSglPI5+Hd7Xj9x+VfgbkMmmIfV8gfK5tPY2plRYP
AkysoM172vzz/nzhiJ4yIsVyVMvH9F/BDsHK8euGPLwDNJjKIQhLYZ7pHr3Mw2/xHxpFZ0ld8mkx
PeRCKy98JyoEvB2/naw8fXfx63mfeGQqKrKnRnKN962Z0/MDZ34HtjNvkBjq692Qo/p6yfFba+i9
MObrcykA2sMtaSdxjb9PS8FnYcDbDsRbS3dneElXy8khQE2cGEoHI+UmOWs0o0fvG0755xDcJzG9
pLIFei9DpSki17nSCaSQl6sPGjtS0nMUQNP0IBcWk3K9EHbjKecTw2G8amGG0/zn5dcZcSVXxl96
EfsRUQQm5d7E17SnhrZNxHDO50s1J5quILrrZiZ6itskCyO+FnPExeCvMh0+BVnbCVr2uyFzCGDd
cYD7kDca6nJOgSK3Jb4aplOzExFhXHRQcjC51RM2Libaws4ZrfD+drRA3dpGZy2BX6UzwOsi3qya
+BHUYAQnWn3hAM30SiLM7YqOICGZHz3Y6dLvPsFo0gqPZNmHun7gL2EuEVEcCB6beDWNrjR1DvV/
41iyqnk/pJ9h2QrJ9jSnDIXpaDhfTCVg8zEEiAc+GUqnjzput/yCSqktre1Or0Wh/xb70VFwLou1
NdCb1xNExw57rTBbEG1kOfs+OXitE/egSkBUY392i89qIl1GdxuiLX+fTiS0XMREfKlZX8+V14B7
4oTIAOWyE+Gqx5cG4kp3V5Yn886P3BD+Z6aWjVbsFFiirtGl90h+b1uyEm0zjLKwniGj4iXLWt4V
LkbwKH4ak6E4CUG4VTtwl3A8fCiUuCdhj/PBUQjt+wVFlOaK388yb2EBNMti553S6fYdwU5rzN+l
JZtXs9OQcHhpLmKQ16+9/LAzy+6exzG/uEf4dx4VTn1TrYAKEeularv9OOzEExPhFOWbAnBNs2V0
HbVP/e/81dXcZgNKaa8CeczUIV/nECJ4I/c+IymX3BPqXHxKwthmK4R+DyMmq9oo++AaRg2e+Q52
4Oymvo3t5ZGFgj9BbR9r9D3r0fz4YfBB50Zgs57iJZpH9e3V2Iaf84QUTbFUrvBodw09/nPIdTja
yenTyfn395hDQmHSx/cCSXPrEOGhuB130oYeF3komO1NbzumeOzc2CGdCDE1vzTdnd7lrYdY9vQ7
yvJALdENuXKPm8O9EmFdSPCtTeKySnjSV5zf2TP7Sn5JUyLxhW6biFpKQ+6potAveu0JxapUfDOC
QPmoKfvAB2ROT7D9HUhdoZMGyBHZ+fzU+02iu2YWhBsiqA2j0eNEJE6wrpdmA2J8q5g6jecQVXsd
2rzdDoDIfyjDf2VKMHUjLUjwD+e3BYhrbK/Hgd5KkZ7P0Uhyggdt6/PI3T113W49mDmOJkP1apit
pEVYqG4uVR8UFXwZdgBsMF0sMTpwLmXcEMJyuiRqe4YORs3ilQKUYhEzcPxw5G7sYi7wLfZart6Q
/9dz1ev0XrFHOuH+vPxK/Tf6YcZSGWxDApy+SszaPHIf8Lydq/RAqi17+oQLJAXrTHErx/OyOpp6
cLIiSysz2gP3N5+KyAYogFo/4dVRZwpiNdMKRQdiqdBbxDmpdHP2qgpuI721CBk5DsWiBJbHJLbg
7oYb0SC+q+j2Y5FCIYkuY9bZvXGZnmS9OJoF31eaUrQaUorjbce13+GWeEFU19vkWmRkzj+B6PvO
rHK0uMtvfvIRk9GY3kjSYfurd9ebuZHpqB/sRghs7dtrU8tnjDUNwDNVonEuNcP8obudn9eQHpCg
m16sj3pzUtQYYUWhQJLqp1cXlSZfBveofiZIaAPp0SPRLjytNO0BHN1Buh4h0Q1kypIHcESElexq
6keVJ/aM86hZ4PG+0p+WxpSyYhKdruRUG1ZXaJWlbNYniArKLx1Tt9FvZb+ocbwpggpRONgA8ZGA
oyBL2jtJ2UioTF0XuhVySCYcEuBMws3Tqsr6AaZHw/jYwc7gHpgR2u8HUpmO0IzaexlFAsDp1trW
H4WP0gcPxo+WHBRLrjOY88Fyn+YR9SnGz+QLWz0nEksPC+Q0uUavs0/1NFqGJ2R0Px6IBp/i+wMc
/w7scGyamDdV+1Or/xrMmMASFvrJStDjogO87Pq3H8LO0dFN8OgkZKpap8qexrY00CGfc2x66ccx
dwWc3IoSmDMrF3cCTKmoqpnr7njZN3fbsRlHD4PSzc97kl8uvNQBTU/doCQly+uX5ih35lqbbNgi
w+PnQtdy4yhpEqW+SOY0jGkWhPk+tbMkdDhcShDX/Oip2OrhwyV482uPZJclxP8op4TL/SoCuAwk
A2tBfsX1W9sYyT9ZbfGm8Cn30qH9KlYf7FkQ1WQ1JEYQLc4lM/MlDdqadZOOEppbJrYgckZ+gMv+
nAVckc1Hae51/qMFsUaSwCoWkdmKaOSdAwmaCTpbzzAm9DTZjHaETorLzQwzn+IHdOtYAKBQ2vPZ
G4hH0tDXzIlqF5ZI5yq6GE1KS8JLhIU9WnYGIA+NCEzRsxFWPYXso2EXFha2Z0kOT8Y9Om+poceT
8IvE41G9iT0vAI/l7GOFQMy1qNN2KEd3kwhNxNcM69W+HB8ctf8rye8VvxeyF71MzYuhLfElegt0
jnXR+9bHpT7zcY/UhTwiRzRnLAIA9egWSfB3BI8exiHZhwInvGqk8furiQL7gC/xCyIOjcSMFEtq
RyDmWpmMPN9HzI41ZNC7B/Wpq/OdUW8klAqk8ALlOdPrgVaZTJ/AS0NoBrBu+QrNygh4rcKiGkxq
8IMpm/ZC2VJC4aFqhnyKKy1JmkcSy4NF/w2khLNaQ/TrkpxejYoqukiJ6D5tqzFISURJvaKKCoTG
kVKoSVzmkKXwf381UQ0MP1ZkJqoMtj0WNn03D/DjUy5UUyrz0Uu7l55nZT0qQ8KVbM4nLSqpGsnM
zElSXQNaVjLjojZTkSJL7rUwTmS4kmgxRt6lC0GD0gCpdyvnmZKFZpDZWkSIhpwlJMywCEro5lQK
58jd9zcomn3yYjtaqayVPWL9QsmRNecTGc/DLkvloTgK1PxreRcr7uvgrw+HfUsHyZtcnapWgKG+
h8W0MH5BQA0VSyexTzqwOwtvX6skln9j4wpDgYnR9Jnf7KCxM8RmExnCauawYtTDJzvm1kSA8iJ7
iuJvAKhJ9GZsFDhGHhnjS45Hw9NdLKiRo3mNfmvsctfcI7hvq2NRbOI3pZoEo9nWbdDnniJ4l9qe
kJHTZo5PIn+b/rWGYj1LaauI1ExiMwECbtaPyAtK6BpAx5YnBQo46K05RmUBC+z9CeTKONmaozf6
YpzzDpKPSidYBjJImC2B8K0R/yBBOMLBEre5LhF6LJw5qSXhDpRGwB2ldlztsFvxPnZI1kkObM7T
q4MIEaEsOO0/ULwyM5jLAmB2WC9QNzBInkRIZ8lKfCc4RxvPb1ZTC31sp/QkEsLRbBt2hNLm7QtI
qIoOFh3f2SugUiC8eyzbyswdzMJpgbKLykZYWEuMylOGwdnCFbDWJ2loZowfRGULEUMK1Ux6vNBb
ZrdxnOYxbfA+j/Imx1PePGIvmobgbJaZbxe9PmLMCQohYSiTDIMjgrItui3/NScwGRRm/3FzLfAn
esZMosrGh/QvGwvIf1dlOWMrblhkCsH4uPW7iqE84YLOu85pf8FTryfhacKDDQ51CNgDAGMBVYH0
XZRDW+yQBITjb8W289jZQknUyCt3WfhqrbWeRWFi7gL8I8iIZ9DFe6cSNMks7JZIqmFffVedqy/Z
n8o9qznqvJCe6aSzkGWZdkUeTDEI469uVw4m0bHLemWkYdwvYSpUsS5TqbWfuBHKkv5A8fBCevaO
tW02Q8YlnP9TBOpih3/1CZC+HizT9/81qUU+J6UrUz54LF/sN4v7xlWVtVOU01YnK9K2KBvvYyA4
1Wq3tliIFL/PF6nGRK5vMYqiE8s2o7MBV7ibgQM7TtrXRoYePcz8xm8ZCFXGNnVMg09SB7l/swwO
RKtNDfNU89L6G641EEAqMTqx8g8HBdxJreh2GB9X2gZLm87erE43b1dnCTC4UZSJi9ywNKwbRZyw
mlwBuQ1bFVuknN9dFXJqNp3nHPvy+8gJkUUMFq7wHx3MefsYfrJcPaUcPHUmCSpv/5Q6vNG+Is/e
khnRVollwBx3+6KmRBBpb6zMwgcGT1sjMgwMGhut00JLUxVI3ppKKn8FCtdnyfUPYE3TX6Mh2wCl
RZKmxucF9emI8Y+BE7ggQn43zFJ6NW7Nl/qkipm0m7nhmF4xvo9vV72j+txwfkh6m18P/7Wwrz75
WhdMDExYcTr/Q3TqDWfuMv2F9EmY8krIslkLRi2ysaJNHwXlS4+NB+NiLz+iLy0/HW8GbczMtXt9
3YOF+nPtLi17MZsLjDQxdrruet511wNfxPYoh1obq9VO9+BCqiKWXTdXHQqBTwxkO6kxHmPrLI1t
p+YWMuQ8VPSQbuSUOj3Lc4PyasPFgj3mcupaoauEnr4ERao+0hbM3LjIUzOqf8VhyQLYGFJxf8ZH
/qrcrI5d/8r82Wo8pIv/rPNTMHJH2TBwJhZdUI3RQ2DVwgtxsbsLOxC/U3K40gFGvofiYeXOjO28
0YqWD5zOLVSPgJlezPV05ZtMt9rGBmc3BOekaa10L9iU9c3WMR8020qS69nlDTJZIaCEcfYCs7nh
ruMjKymD8d0K2mQt3rrZ3/z/ndlPBXe8NkF1NH3cUUgnROstA4wnItVceyJW1gMwwBNyK2/JpCVv
xSpvKTZLF2436q6HDav1/+jdpaXdnncLiIofL9wkOOZeIsKZW49FXrKYnKnKalAxrSE8CIRW9WBc
VOtzoVhJpOTgJJURPgY1oLO5HjDukpsciXjT3fMSjP6zQmC9O/8erpS6BT8pDQn5dE/GT/Fcsq8x
3xQqSFgvpeWjCgSw6W3P++XMdq4NgJsAIOL8w4NTew2qXydUOeMNq0A0YLsPGBs9Qn1lwzmjp1F8
RfI05Xb0Oo6BieuBX90def/0GieZwzppsj/7bFWYdVp0XdHHlKkbi2E9PRDxllZbAT9VhM6oSm4k
YADocRBZ7YQ+mwC+yeBfSdH5yLua9JDLEyQl0qZmKHEmRpNDl6xX7oCnmIMMgEJulSwgTOwcDwgy
ECdTIfkbjQR4g8CqdUi4h9ViyvrrRjXL6muOzi72GXUYIeF1Nac9r2R/9T8oCh+HMS9yhx8m/YlV
cdiMMd5F7zbPzScHCC4FOJ7Jdo1u6a6adUP7BQHVfYngCoySu+/EEFzlRc98sqwZIqj//pHN6IRH
P7QJs5DxsRh2pv3eDPIPqnSgFJSLDuH0b3PlFyH3vk1GI1Y25ybUSTWJDu/OO9JrCSNhHiGEpnks
maw3DTNvPpxhveqww0O3ptNFzZPwnyix6yz6Wo+j1MeUAz09Qevzx4HOzXThYYMI3Z9skbgUcGg1
AoPYTvwnP798/mzgAkG1NV+dMM4b3R1x85WGiwb/97suVlQkbc7/INEIPgBKLbLFBn3nltv26bjt
jx6IuL8zudzu7UkpMAj67DAFJCwBTQ47mH0kLc9Jope7H0Bebjng+c3eixBb85D4fcYGoBbDC615
beMsTIm5Yq5XZhstIEyhQlodOMyZHah4fcSLJJVYBYAyioGSqyab4JTIuDDQSbI7D2N+vEq3ijYl
dNtmQXO2HnaNnLaptAB7MlJ9KxakixH+iiZHQIuD839M2IJNSNY/QiY32lQiBuiTuuUmiPnW8X2r
RfkV1LkHbCXXHflwdUnsiA9LnrmOUSV2ZNM/QGj8sBPJkIQe3WN9DR9Hakb2+shIpCOfJu2HqIS6
Y7cy/+7Yya/N+wSC7dQ+jGCFoQG5kECblGR78C73RyzmatqKUVIELhg7/cvdwiOa7GkvNlFMuEo4
rfkdyPzKqBPK3uPm3FClKw0swqGPTBL+S1+KDL76HNxN4nI8zQ6bmaC4uas29pcx4hUg1wsz+VKU
e3A4H1l8D4lg5vWcZEBMAxH7Wb8A7yyu01L95LgPOENNqopXgtSlB50aKU7Eze2PR3z0W0boUkhj
KQC+wk9K7bfYqVOg/C6stNDlzOkry9ZcUe6HuGFooZK/o/BOVaNCzrq/hrLQ7uFnP6y4fgn9OX5n
FKjM5taNKH/QaQ5dkZOe5N1RxfN0NA6MygJFWNieEtgeg/5C3xiktTlTGbBrC54//IUd9No3r5Ks
Qi/L0MkdqBW43qED5tVCFKZwMTW5e9RWcSduMe3LYdaesMb4t4STXgMbwL4BeNHfiJ/bg4v4TjUL
jwGowcjIIM9PPYNE7T/y4R8FN+oiQUspM9q0z0EjfwG+Y/h8gNmhoGd7R9a47iVbPZ6iKcJakxA/
yo0c1+jek7ZyxDXu4oKOB2EBHKdoK4tmM/zKUZB6vc7WMzoJELQeBTgPgWYQ8iSnzxFZAPHAfR0F
ZUqG6g4+uBytY2WI/BRx8lOROE4efbqku92J2vKeypo3oXfAe5P21VBjOHkuFqGFTAfQfV4rWUnn
Tob05sxrYOuYm1WyiUaVSGYSzfIpx697lFFMjsvyrVj8p7bznpxzYWqy19Wx6oHRw/IvFGv6XiqE
4+6OcsxNn+IZfjE8IwBzfEC40ZkerYda1ESwcZGcrafj7IYsCtOrEKHiE9AEZP8xf5tnJu55m29d
juVWpP71NRzfDjKaeEpRIx1FICPekkwATdwgW1VtyDsJ36o0NDL07sWq34u39t1e4222MWwYMu1p
BRXew1hzkryWFneZwoc4dXyg86l7q6F3R0WvubrhIov4HO99gipSVtZhKqVCOY1Hgezf3U2N4qD9
0LbfPn6nuyCOSqxjNfPKYetCmyChfwGRDPAY583/RehBDKWxbkuG2CDFobItbACtkP3xD1zXdfk6
4f/dlQT1ashnQ3E4+ao4Y7zmGIM/dR3e0RE6XzOamQmr6TPF8Aw3Z6lnuK60hEdQJV3qd71wVHyF
eagE2KFGmP5GJBqQioXe5jIlxohtnagKTMxA33H+t9rFPctCOcN1rlEa6WPT+vUhbdvcWzQL5INE
iPKvsZWLOLZIqC5JatAceALhNYZhf6PRKPxeuLmpvsQu+E3w+8vNR4n4X3JgJEY0oVNqVVbnYReH
ATSio5lqedtcDo9ZdZsknLPMgRLZRRktVTzqnHvJbS6GkJ913GdHTc3fjuiFcpu/ni/CzNMwgGG+
F9Gjy5AZsLBZr3RwKKXD57C8GUutgvKX+PwYp7M90ZX7XNynTQka2gUmQVvHh3TvL97UVf0Xo9JK
xRVe9lqr9y20MxW+FPRkDSYFpC+DO7Ar8azLhn+4NYDErMP2iFQxqog4RTcElnPiORU5ZqgUSAge
bSx27+Y62zKLsscn+LTHESRDu0XtCGi+0V1xxUB7A6vOGa8Ol7sYAHP3bYZl/UVpztiBv4UifIAy
lCkgdN9Os+h5nu6gY+PCN7BlDjPOLMKkkFX0ehGASB/uJLQSRAnu3YaBjyNPH8OmWW/voZm0fUVW
m8l9p+Wr0nrJUa1Uua1xVV3rjQ4dSi/rOtzT8QDy7P3YxOcxN1ZUDE3ua3aaxz28hf0XMZSHifEc
+wZ39J07jjswQ03hePhjIXlJw8t2SABxyKtDqgrpAeRdUGzNTpbf/nQYZ6AX7L+P0V1DOSYQfkKM
58TgPqy0HE2WxKEKY47zL8bfOEURrOcUpxnQRaa5yhhSf4eON33HKej1Yg0YlSE+zKahN77je332
NXw4d03PlAfjMljHZ+AKghTmIbskklJUd0em/zVuBOE2qz1hnyRTdS7e5ogoevURRkWCGnPbgoVM
xxTHEkJLXmKCo6A2zlXweXF0i4ABfhjdX8+dazJGoojHRAsXuI4YrRRXWXjEhQiRUlqS1ybzCYLp
p0iCFG8vt3+YLH+NGI/Q4K8mhnDSQ56zDrSCjwMtAq6It8eUl/3h+tRVjuETfpfttwKwBpaQvcgJ
NE60mhoUyyY6KnWEM5aEhtZZrMvETqch38En0N8LYpXxi3N8EkCLwIZ5s9pDoHie1aUC8j7EKHcl
/cOqnAI2OcpBM+2ivyhBRonYMZG0hdiA8rlCC9Zq0/s/Mxv0ZPZ+LeOMTvoFSBmJXtIGA6Jfymik
Qe8upXzjc2I0yqGExFZmTcFs9pjrDZO33x33MVXeOj0TbUuPayJ48JR+IeZXgeKZgM8EuWznZmts
AILWCclEIhoxYwJ/6wlm3xBXPxiCfmfB+OkIu3rrbjS3srJAsFgYYgOshRflVKEnT1DWwSH1vAFZ
4NGfP7ATzlah9KcnksYUxWQpE/ZzBNfwSxFj32cLynehSJbCzM0xayVPflAXlGj9jIT99hb4eIcf
ntTiBaDsmWH/aUaFSwsvRxQkEmNrlWxOL7KJ1CvJ8AQ724WCVVF633WuzJKuA8b1Eol9eOD7DA9r
NTd9lRs7XSAys15q/kSPlgEydfVdAv/85L+8O5XQ90DA9T2tVisTmYg/pRw8Ns6bbSkG65zpUY0y
XaWTcjcE/DLTCuPOA6+YxKNieUqRzrqTY5+3F7YP01LOdODy+HxYTXnWsmgQJc0qh0SDTdJeDDKQ
LYWYTRCY2mtvRgjovwvR4R8Kj71qKgc096nZzqactdfHAHRZ7b8q0I4SkRrwJqbGR2ZjlO7N4as2
LWLUeOWz+OL1BVclgG3Nhm5lEnFTIRorI7B660RHnDT+q2l+1i/52mfsa3kf53bIWXl5JD6uD5DI
9V8nQ60Vh8PTe3o0LJwfEemP2y9VAQP/B+g1cVvbVwu+d5ATGq2NiBn7wckK7MBDgJvyrYjv0Pvd
xv96rH1DqJB8t/0zrpIbwcvrN6oDoNLAnxqFRej6r6bUJrFubWKd4u8mfEUimJkJsfe4O7hrnlFP
0Xg8xwcCN9Cvoe3c7F5I0JppUVlW4lw7ztsFPbhDvvp/C0pjfxZrAZoKVokXJxtYsuGeGS2eQ7W/
H4IK/rPfIto0L7K+udhzMho1HSpQG60mdax2LQobz3h3Gn0bD1F/W4wKu0SAavBPXX2lWhb8kZvs
xqPCw1zjk766TojDcXhT9jOiCamDjihPNurmX7DBy3rr8+JCITW0SRqj3R4VGsu667w2OEE62WbA
dsMnYGvQ7AbALNqTP242nKMeTseOBaM6/6TROpUsjQfhM+1cDSCemJC8KbVh/0/z/IYImp09lqnV
hEJYk6cx0ukziBcrHr04SOO/JJ5F89nRKPDkNc40WgKJBuxdPothzXRrN3a64SuflW2UA1mdxR2Z
WGotAGZT1pUcdBLt/OUtACC5q3zaOTArP1D7CosBHJgeGrYjLMEe26wif0SYd8lo8Y4LMNy/20+o
e6+WpU59ffdMyrpg34gOCHWokcZjeKIP7p1VgHXMkAAJpetBHMR7xcoumBJzc9EN9hu0GQb/Nu2j
yRvkUY/4uRRKCd3xs6gPCnrcBP8M3syonZDNzWloZYllfCuNjwxjbNI8uTkG0iszThVvLR1sRjEY
dSgSCLeAx9mkvGhVB/Tm92MiSXtBqUFBUEgikutlE6NrmnWQj0+Hv4FxNxT8SNJ57iObaQKCgRV7
HX+bIoMusBOFTRmIDs03bXApT1C/QqvOgbOtLNeQHOYi8fsiJMUIpTxLw4pBAtFdHd2foYucV1RE
1SqLcIl7SDiStGKKcNdRfVN9G5fj0GxhaMKXalEQTTtTsZF+LavhxJTFVQswRzT2uw3QbDUspMy8
6nEDPz+O54jP5HgICW7Q7QwkbuhpeOdikv/lwHKVD6WCDPOFgursfi3/B3j0YsRCzeCiJsfMX98z
oPUQOw8dwx/0w7cYQpk84eYEL/lKMBsg+/a3orlNblfGO90cAe2nUJ+WoM0wt1hRUr0Cw8l+KzEm
pb24WR3hiJcmCDOkqq1DYnv1GWbgDPqpED76K4I+IqsoziPnk/HBmwVwUqr5l8zKAQALe2oYn1hz
VaQRSEL2zb48B/fiklrxkD9JxcWDZuvYTchbDFn8Xo4DAHg1qAU010eOMR8zSgddiLo0NOegBdZH
wGEZ9+VM+9TYEEQV2V1mDr6wjjFpbv/h1ONxgAdDUVkEXSaKSrMSXZAGDL0OC3bT5q8XL3Bqto1b
Se/GjLmBhlwT3qoM8+YnT4/6VSPiSMwdXudiNBWdrPGeVgOAPYE9VzNK1470u/M59ykTYet69UfJ
VOtwtRP25DqIgR755xIoc/U12CfOX8ToZG1jaesug94moAUR96oNNOQqcZz94JB9sanpDY/0LwkW
f7PWRSpyACHgRkuUxjnHa1cSqUj+UIvwGBQ/8GtbbDDfQEGHFwPvUgYhBuEqe92Hwbss6vnkO9HT
EczSLZdw0jxqqs1mfd/Cwucy8WLRCROh+jg1Z4fzdvNXBMpMwhWvitg3LplYWNWXxfheqVzYXoR5
wu8O2P1f7S0r/+FbDS/YrNkQpIjvVz8LL4+m90Ubgg91B7v2gkfTHpxI/+aSEyPFbrXPXY1QCOiI
YnmruobOw56PiFGxs/1SzIocTbArqCygKcWXfZIX00PYETC1Cm3W2smWL30JbaGaHfS0s8j4m4qu
Ur6S5a0zS6gouuiiZcHWPp7k3ZU9YFdnr2sOEbMraXv9uP6EGQxyeSMdmEHU0VHhvO5rIrlq/G+E
Ia0EM2PoeC6CpJlP8zmFCyFsHmxUMvqW6jti5ENkH7GKqjTHiJNPEm1tQN+COLgZwLPZOMJfbdVw
Eu8NhzUCdW7j5v6oqgonIuyQ+3GylYn1usF0zjxcskB80NjQu7lzhzGAlXDZXk0I3dqfrC7J5Wqx
XMWvJEsNi9U3bvaA4+8ukF7eSwiEfxOtigbsyGgJMVukzpV5wcHVQFrlhDO8RfkLQp+JQh8sGnlU
boSzjK1ujSaB9sZrrGQ60P8PQ+GU7yFOO5Z7+wDyW806wtczjM3H8PERP9WiKfwI6gi1T8ixtkMH
SOfd4BhYP1/x/gu8NOlh/EmlehpUfOv/DLY7aNSW20D59qdWXaWB/uMDH4H0tHTnBfKNXxvT5Bw3
XpC/sy1PKmBlTOFyv9JVWm1+aRAd1I1eDzCAq8m/becz2KI0NXUWEPAlt+mGs2safYZHgFERbKxU
uzXl7V0dcx3KS7u7/m9EXvGH1ahLeXPZV4KwJZfKKu8uTISlB3KiaH5OkZeWvYXHnJE+IVUVosId
B8y2XlDU+ZUDDDE8yNvm8pjO56MKsOWADQlDkY596V0DBdySfj+y+WQXPzVXYYyChqqmq5fMZmxY
HnPOr1ypvVPDKVCbaNlzjUZ9DVt0VW40BY0G2tn6c63TNRqQVyu12LEoYbO5w6otur/dILL2/plP
xcb6oWo2eoL/MzMevv77IfqEVNDKHjJaTwti42iAD9mIOJ3n+ZmBgrKIG8EhIibGkQXfBQMvQ/EL
qQNVE3bJePWB/X5LVEujgwGagIZ6P6GZGUkVQ5YB7GvG8TRd9ubU+ScbL4kPurJN3bFhS6X4D9Lm
9aXGDy8pic4nUaTktqxVf2DekxKYKRP9E5hXFpNgnMt7MZ+q+AwjY4qIhuUGq/X/c/kCPD8obBxy
jQ9w+2ks9uwGfcvamwY+nmbLjwnZ4J/aj04eAsYlAvGKIVeG96LxsdMBGSIpsgylejj+wSMDhOLx
sLmCFIcdiKeshkbQPa30K5wfyApgBoMmmuxSJCbMq2573XBtfE2BM8mrDOg4C/MuYUdfH7teiQBc
NWisXIuH4XhnBAnLQNOMa/Tj6PqPZVC3aNmh3hTfIil+ojZjDc5+l6a7C6p43AtpzeC19yUqvH45
VHVktKfSERVjA3S5ZgRuVATFLTJbBHu1H06J35ijaxIi5c3nC9QWoGrvPE11agpy0d4H219IlhDE
/ceu+4t5BphUwybipxODLQrnEE98VMt0doOad55IAlNJ1PYmHFlG4BxjKwM+rVpsgDTHNqYV+vP9
3h42lMwbpq5tJ8JexCn/KitFbydeDJVmZXyTZLmn8Wz8KNW9QKy4WyexXahlcNSGbdwFQlQeXGOG
+slbdMqZ0BM44mdMzPt/jC9KYCXgNFbTmutVJdLO3kouv967kUlmmli0qZcQe15JVbv5qHkDYcfa
lbyXt+b5EBIPjo1L3ecOSWrmGvQeQ+6po03EbUcw3NlEKjz5JpSppXBmg8b66QUtNQxz/H64JQ7R
yirXVE4FetPWDZehIeuka8iTryEmnIvhY5MNF+esdu0VHBdZZvG8XF/4Tx3wI9npWm4r8V0Oe/Rv
M+3mGxarDOY5JBUk36V070gGjhd8v/hPgmog65OCxZjF6Vt25i7epXUssZahLBLmQVcAAp+8yhrQ
hIyJXcg/X5ULElkj2GmkDQk+IOinNSFkybPVQTqnEMYXs/vYzLyNx9yZT5VuFZDs8B+KrMwfZVU8
cbYS/zmPvL0vxWNVmlWuTs2g09NW9ysFgQnMKmSwOtQtRuOfFa+3RFO8B47etTm0GFXcH+ei0XFZ
4MeirUkgvb2otSqBYY1SAK5xYcbgDKjr9CYp39xpI4ph9U1hEMdb3q3i0uMpT/d8/yVKOdaF6gwP
7GDQyJxNN4ry3WyLdRjq459Ohc91ax8KzzQ6jlNiJ/pOZA0Wa9pAVXp4Lq9IhIYZHGyRyIjIOEPE
ilQvOHBowpJFb4zdhrBfDQXoiaDhAcIYAVgDWHM74emkuod2cusk436DbRlEbNkj8H9zvB9GQvm0
cw/cKPD2M3q1p97DZ+Ywt8kuy+iieZSOPHToDut+9VlXR+i0hUJEFGcK9diQKLySr7eyDHHDZAX/
aRGWCChB0k0KYZjkx0drHcqDtO57gyyICIjBoXwXv0TViBEGKbqFfo1vZm3Pl5xnOKt3XuSzeNJu
iZ9tDY8oP9VDYpBTKpW7U7MmgpY9qepyookAfDtP4Ab141GKXpklkmlten0aEh6Xg4GEp/S0iFml
xUjaytz2mEUEkiC+3E3431yij+Gt/ZaPQu5iANKjT8n+OBeCsj8QnN/1WiGAbqz1IBAxiOApkibO
9jyWdhntIJ8VMEQlNQPVfTFV12TeC6rab6DR13sB+9v+DFQ/1lxH0lajxRRkELogt921ljPsjnmq
xjR3aBoLLEOjwHAoOqpEBiP5IfP5U96NJm0Nid4fenfvLEoao1G6ra05GMCkyRirqTLf+fptG5v/
ZvonMTVRpaDJ5UaN4OnC1Vi5/KdZbkWevx9XUBp38PWuHnNdah2LPMlhxnyyKK98LUjbjzvXcmOm
e/QEJYREPOOf/9lnIIN8zSxviHP3Wvjzxt/CFbXARzQwkVIcg0nq87kUB3MFLtfs0ZBujOl2M5EP
3d05kaXNaRjk4cDRDgOrKVjmyTcjNHvjBUnl3O7iHwRqrgQ9P+3doikL3K6+23cIU4DEjuAycQje
k4ZJWJsq0e+3sVYj2cOY9kKjVBWJ04zEhG44YjNck0EG6JnBdnQxkwhn+H9Its5X+KsEWjOEXw6U
wWEtxq/0jbt6dapzZoyZQFyW1tUXslHAQ/FN5QRC52NMs7rxXCUfpiY/0IE9xz4QzQX+i7DdQpzb
khLXhhndQVtpIim4sKGuqcWaeRuRjrXMY7dgw2edovbLc+J/G8zqGe0dk1p5avWGeEyPpUGM2d8a
NZMkuYH+PVXhgYJ0kNqBRie4vCOB9JIcLYlF5vYGELGlaMVL0t3FR9526p58ynaGNsJiI2cWenoi
voZfsHjoxOT21KykmgiuXFdSJKGkZziqy4sC4RXWvnpo7FUk7k/l7Gkh4yv9dDG3vs7r7wN09cor
APjEBm5HjiLWJZonnjpYD1Sv7amYsh/MtP9G0IguFmanXMBbcHLPOCdn2iM7VjapsLWYlLxWugq6
Ah4sN1ClX5qH19hmZXo7Qq1LpvoWAbKk5Pwfpvtapb+fzz1/3KBhBUaVNN3VHMng1CxtUdIZYtqe
OYr5YsMUHP914JDvMajFeqlRCF7w4NvqLMOrdxcCR4RDRgH8dnnPUEn2FHYNObVEMoh/yOD7+EEJ
k8QWyZfzGdRUqF5ogpjGtRdZ795lR3gIuTCezVZTQsqyLyV93QOVmaPOjj0ueK96cj8KHNwlpy3x
yrySvgp7144QHhFvkAbicA+BFzawFjDutgRFwKxowKCMJvo72wngiDGKSG24RTdNgG3SEUycDKTu
PSttaKomj1mLs75A6I/aelt2Lwq8eMvdNjiRtkW293MCK5I2W/vpIX10pclO09KVeCjicW/LAeYC
NuHL8z7bbWTdHo2I+yCgX2fL2MXLplJLg9U6RJIyjh44e1DjiGwKICnsvDo+Dppvv/QtHtJuNEc3
h9JUlKNCXyPv3tnOIFZ/LtChLQLeUw19GovX46HLMZjh640U1tmJcqwLD+iExHjqWbOblL+NGSF4
IzAjTkK/J4PTPYGOukxC4yCHk7oeL6Fw2mtbhx2VXY53DykosuHvZwnFjDKHTjpqLzCYbRuxo4vC
O/77KGFdlH1BnX8JnCRI51aJFz/xUUHSBQVw7DZsyT1DLs+lAbBIvCIEeQvBMMJ396N/HjNNIKks
cwdz299sRwncr0M5eG0IYOtC5c6JhGKrm/xP5ez897lUizQPMgyMCelJdGgCgWc5EDVvEM/YCwDP
F/TuwXqATU07wPaUwFLDJ16uNOVcqXVVZOtwIqOZzXandSsD0vU2eBgNXcLsjQaAvDCyFdRAytXx
509DsUZN/KxfinQGlIQFm216IT2rrtuyOuZvp/YTQ+b326orfJ/0TZGHafxswOsYjYOI3SOFkNxp
miQwi6FIzuS2qqOQ56sGtOsVULotWwsanclTaVsk6vSi+itxG7rt7ztbV0zg+RThFnvbCy4d2f34
URV5N5+YfqtYRRpZyX4Yfgy6W9hTfRwefOmiP04l2gi71iM9VmgHMWsxEFtwytrIdmWzRgylFh/l
DuHj5mFZYLAFzEPH8jcuLA25LRQAf0AR9zZxX/G7nK8bxu/bYhW4zuzbWK6NJ2GSVLOjupTwWV+R
7j26jX9u6qPHER7ofhOsEKCfmnbE/aaBl6sUTpYnj8mpFh0sWrr6ef+y36H2vp93awtKiRQJcJ8k
/rdBOIQVzZtw8vzorSj8tK+X2bgz6F3o6rywVk8g5oJ2CP+Rjb0nCumIfaYyes3GgVAaUdkqHoNA
C7liyIWVlD6ku2MI0xcawMlaOTADbUqJMf4gIHARCEp+4N7gWexjEkpx/X3vJ6KmXus7/bJ7Er3W
mvVi7bkaixovR5DHL9Ece4fHhSveskAQYL7lxNImJm4OrWr+KbjMRCYCs/SaySNWe20+wIQf7C06
t4uCcOdN8ARLP2c0xQ8cWLTW+CpUWE7JKl9ga3p/1XF7j4zpqxmQq4EAMFAA7frLDgA42wEyEoaA
Bl5K58AamQDSlG6QZYQJzA5STMfPd9vRFCQu/KSV6Rgn3TWJjruD5tnxRoItRhyOeOfUQ4pVY87w
ji0OrKyTmTG155/0ULZibODUVdN8PW8UTo0kzv6CmRZ7RE1t0fJ4Knr7akQHb6g2DNizcHJ4yis7
z2Fn4lJoCrpCrss6+Uv8yPExziF8L9i2gSRIB1FIrHmwUUIOQ3N/tlGrsiQRCRG52DrbXljgTT7Z
EOaTu6cFuy0yg6CGrwZaZBbaRx9W9a/vau14uxNpRuJ7NgiB7Kucy0/IuJzwO6pvN//OcUMP8VM6
zvlETVY7UIdldQvNqCczeHg7mIUHmoi5URTbcSjbQouDetQ50MzMsg7e1Mls+fOFiUIfd+54Q5Sr
U/R9MU5Q4qdSIxxlGn041Yp9Cn0NRvBj9RwToKQQ4Ybl10nmYnzmqFSVklz1y6vYy/45PymNASAL
tmuexAGeGSzGoHjFq2rEqiQQx17Tj3GgnZnz5j8Utk7UyuJzNpm8t/WYLEcr6NmNEiRK9Sddcm5F
QMQseIexLBmZaJ7o7exqzIGiJOua/sVEox/vSMH4KrjHQkhit16bab97isZK5VDejo+VTvzFTary
nrij6BouNisQtQ2wQiB0z8vpzYSCqAYUvdoga9JE32gMUgpAlJDZAGP9A/e6Wt4PFKkzxpnKoBS8
ioJl8kmFwYTEPRQpzuPYkYT20HVD5zNyL6dw6Vde1I6zWXYAmLMxix1OvvoVHvp5EQ8A5/EGcuzQ
PVghdIHTgxEXnXiD4E87LexuAhxEedN9oXIYagQ6acE3dR9FOUMb+QXTvo+nwgQqYYOkzOeV3TdT
32Guf38dpyT5WzEQcT++AIBB3ey/OElP8417BjS8xuOE07SyFdqQlesyGsGtEdPSqWXpwUnv8j2b
XWci/Iet9HKIhPcZcvrY/4rTTBX15FaNzPB51/eRhNFDzQKjO+RDUZJVhDjEkpg3U5Y2DV/2VjOd
DdAq6DxkURyRWMsHzgpWG6UHoEuKVAycKEqJT5iQs/57cRC0hMoGc32lMZgFa+aaYqDgM6MrpyG3
1MHLw20OQcwQ2TtxZFOc3OKGTT1kzggfMb+XBUhUb00qkGQr1EJWIkQna6G1BhZNOBHVlz1wIea3
TWVYoBikK7oWnosHGS5sqgR69xmMNESA2LaVxb7zeQsA1iXfZgy5dj+YozRfKubiqidOI66u7ow8
9SCdu2FtyXbn1cexiAMQTg/DDH4zznigT3Vor9gFsMPFQlYZO70Jds/94zJDuI6R/dYNALHq/axn
lVd6Ogs3GwqbnWy66krvUXYol5cwnlo6BCrYOq/8Ld/bOseTrHN7OD1FWEMkAcDyZHv4qJGyNXJb
jJzwNPJ3qgiRe4GNgdB3wq06L0m3xPkG615KyzQ7ZaFHfAmoE0KIV+fiwDYzJVLvl2bem9L+tpSn
Mzv8awtTs4YrWataePqsds/QMv8z4KpOtY55LEpP3mMApUSLFzJedpbAzuzfCMAjDGh5WA61lVg4
NXdQXBAJ4QeLP46F5Hnit8/JtXSDneSHUu29vT17CzwMVqg4iuwNdMS6ns2+h2bl1s0wZnIo4ZCA
1VzSAf1ykrYk5xMAxukfysRh8fp9R/zsUd41G41q0gdrw6XNlLfeYUIpyfmfKTjLp36BRQDiKaPE
fA9/omFcmlpD6mu70W6rY5YxQxQ7qusvtvjEh2Rhr9Lkg0uBkn38J8Cj/h8rJKuwIG0CBqPSSkBj
hbZp/aGlw5jX/lryvK9TFeg2LibXVRuKWPidT8juuNf8vRutZFBVibkuOAGvdZlKzarvXlFikRpN
THvSkDg7dnJMok+O0WoHfEkkJLRNgeRjqnFY2A8Iw5LIMxxXjc9Y9PqQnO6utpSlahXD1r1VLpKv
aqHLVfhXKJZ/oKvIRHAjOK4AeGr7CrDdQO9uBn6LeTNlsKJBBbkIokmepsjwR7b+SLrY7mVK5Ur5
7TwEXg44Zg9DeCFmnstET+ciaeUHEv2deC69qxJ/2KAWP8geuhx+BFRItHVfoC130Vm4/OMZMVjN
+6X6v57JUEL7gm4w8u0HIkck1RE2Ey22YgLSf2Rkdtqqg6JITmhmh86qdAzXVAakzOvux1lW4vb1
pOf4a+WgcOwP8RI0SnRgYC2GrTRj5bPs84/hqXnipPTtK83KFqBfYDdcA7SqLcJWOAGfr8LFQmQu
Waz1drIboDirNNQiieL8OZ2udmKM+aAXW9RZxvyIrGyW1Ho8fHnuu9T7OgLjDiFpqpYUsICVzt3X
wgdTyroOb7p26DpvTKCW/17Hv3leRTbcliupeo/r2biMBuJvr+cwe12BkNdFjbUDhOFvsmdlUUaM
Ej53AKkHTbEb4iLZxPqoBSBWReqanHJ2C7psVfNBE/J5OLbfanNH9J+O+B79fHUBnxFapY3u3ggx
MhM3/+3VW15TaQHMCNoTSd1vdoc/XxFE9h1WJdRQCkUUid0g6gLyWSktkZ3SgBboA2roOiDJlF0l
1eE/LyP6rGbvmOgBDz85srmY9ESIdwzpw6zW0jhJ2E99OToZMnUkWLXLtlTmfeEX0nwFG5Rj3Ca2
mdPZjXxH8OwMugmg/NSpI6oMEt0e8VtCuLAO7B0zYiQ8tKTTbZoHR4Nv22R67+U4gvvMl1vO2xAx
XIhRE45c/pK7EjNTDYo075lM8mGUlnN94aeNzQ/WCzS7mzZQFOF/PxCUnvw+9vICQ4WyAEDRXkR4
IWsWcShysxQC6UGe72qDSUYXAMeYdj1SgK0wpCge9ei6E+1cQE0hJaAvhn1ceZq8epAoo4O+PgXZ
7A6gEwZ7WJFaZ9Nc+CILbFrmYVTTchbsdpJjTSi7/aStA6Mcomh23pb7YxzJlm/xvCdu4v6kgjfZ
buOZvK/XtDMraPpO/YeuPYjMz8CjzZe5xX8yANmPoFo7ADnMAaAwqOM2W2YKxjAoQCBuI42AnVFv
WsiXeLJ6aQ3bpM2HFqaletudMKA2dmasMimt5U1F8CyYb48yONIRVCSfwenyoBYoYrkoD29TvTt2
i9q6qk8BxAzfn1sSroibsIe4ThQjNDrHeQ0n+Yh47feguJ8e3mLE2wEqRcSkBm1Dbqsy6fBaaA1p
UjfmvVFUoG9/y2sw8LcyYMNvSbGnp5LPP1fOpc6vcaRI2LTXKBaFLAXP0vNC0laBUwJ5M8JSnDOU
2s457BYz2WPAXK/MW6dlZwtkI1wHAP1DfXmxEWqQmH54VqzXJhIuur4m/aYHWIUFtfVLxNdR4L3h
KV1pWQ5r6BAiw2fV8BWmykMLJIb6TUkdFiLKeWFrFELb2z1eyWkDZwNxogFuZ55tgMjBGphYAlPp
r2CILosNpi5Iy55cjUfliy9KvASByF4K6SIPmwTcHdYnMriMO0OL4UfF6kRE+c61cuFvbgmZHvfP
ihZ8zSbdHgLzInzlr+a5liQBMZUEHIvHXj6hFRHsEOMroboORiHO9cIpNOJXpNqEEeBknGx6SdNz
CiygXbnEiNEbFzDhfy6xwJBOfJT4ZGxz0/bGGB0v+LsOoolnybMyCV5lFaR8xWj7DWh9QG+xTo9N
7lTpbY6lLdGkt8GkHeoXoUIPPtpJRGXgdE3iDr/EKIfg6Ff4xdboGmet+iF8Qu2ofkNPteqj5oN3
e1YwOn7z+G7cnGeaBdwoxlyKuph1YjyEVUwKDVwPnXg2do3nADldVlj+IPWvRFP+OZtsMP92rpG6
JFe3//FYWD5ebpdcKr6IBzn/vVwWrTXoIRzLldbKsoj3lmcBuwx+BYsAQ/TT9bSwmHYCSruTgT9S
o58WVWB0bRJxvcFIqoYsw5G454dWE25Hi6V0+D5UDcVtQ2/iboSomoECgFRdNCm06Ldm0Ocn6o3Z
WnNqCENt1uxiIS5ob6MCZn10N6jh8vJUbdrV4pnmbIep8usfOUTxckmxcrZTUQBzc7PFQQ8jbrc1
ILL9+iGip4hgnj6pf86tdZLwJrWXkFwjpZ5sKDKRs9aEz/IJ0Ynq+02zYDNh3Yz94rVfAN6yEGUu
RtskSXC2GmzpN0B5ZhAsbTLwJUYUZ3NAfPvzsilIddA+USLVEHoy/wNyqm+NTXJrnhOLrV/jb48w
IbVUm+ZIV09kKgrMXSASelvq3pdD9gwWsTpcBzkVp7cGe0xWwkwtsc+XSXBHJZyKf3ZOTpmjo/ZL
sPPdZ6HmACO/hw0bF8uW1TxTY5kRg86dBz+CQ2fSFUWjMfYvEL2ydiXTbzOVHgHtMtD/jI0epcrP
JTUkJrDPxeJVJjkePADXe0DSMRr3rJDoW8MVKHXj8bBnfnqmznGC70Ab3gX9a2KwJfliTFmJiEIO
o4bUcvoGAK868g2pbh8VwBKxHHKUtQ+JJycCAlk5BKynSfsm4YYP7+R+5/0EhscOUxPLYTg7e4kf
gb3GqnIjljoRL86wNs5/JD6FaBsqIrJScJotSiXjLZatjvULjG9Qn6PIoDvMeL6HddCJAcgEvbBJ
Yac1Aw4nMDCy6JwbnjTIDVn8v5UM7KyUC6QT9/jpArQu9cFbXUsIIwrXqdq85LJ2cuRWtMY9zrlb
ma85JZUZaNm1LAmdB/uGmIJ0l8a0y9f8yeBKrzdmoGWKgC9CNTgNkffxxzxZsFbmxXKsZZ6F4Da7
S46Ld+Ief/wFFYfh+RVNXo7pTAGQFqrlhqE3r84lmzH3pCDNHaufGCiu0R40estABFvMIWD64VRM
lMyB1L3MVRJrLFBIfXmjmr860o5RMIaJTwz+acJd9q8ASusd3S3/rhzr9o44owWQkVBEtuvgy7qv
+uJJWKCfZ/AQKWcUQW6CenZXlmWa2dliHRmY0YUlgzq0nprkxKHvBQ9pAJjj3Bmxe+SOFEq4T/MO
BbFc7j9iTmO96QixOz7rTTW/4H1e9wJ92wq+HqbwpfFZbqmJpvrdaazWniQiOTjrWzlXZJOdpT6U
SGzSLMSG7LoNUes/9xF+qVPppHC71fBgeu8rFiXTr9l+Kou+85r8PPgMfwxQvLfzsElocuZdp6LS
iyvxmcf6Yqufqs5Fytc62LPTXOqRk4gVns9OcMFp8BCkxuOHo0sFYVSspCGqpEkTJ64G69Ghod7q
Xz9xCyh6oYeQAoOW7qe7uxsqAvoLIEjeeEMPPrj3RJ0Mfh2VO3hzgIsINUpUH161JG2EYhdVBu1O
drgPPKj8nTUsorrQnFWak0nFKogRzssXFHntx40+KSeH2iKHCn2i20tTv6XD0hbX1VyGv6V0LRQx
N79aVUlpiAS0w3xZleZCcshNAgFkreeIVq4yb9tJqou0PfkRsgo+YZhNvTAdEP7h5w8dygH9RNVg
zaMRb1zM7z6/4Ja+FO8HaeWkBiog6MAAdCRz7mNwMKo46Ee1DD65Y8pFqANb0BTrGjvNDue+bEcX
65ugL+eYGfaEYQ3rTBl4KgTh1udST0hVYY/RnwjKMa2j75lZLlxVU7hjJ69bJLoavvRPjq9S1n/b
ImIElXKFdca78X7DVRksJhuF35dC8UcXDlYBm0sSqUB8RQw90L5Uwop7faA2kP6mCoUnv/KoBZYt
AAA2TD25gUnKOyZFOAkWi14doEqFAhaFsa2Vikx/OKhERiPtv35q2AM2v/DwcL6gDTh9Yvnh+4bV
GVIacOlErJfxaIiUwiJhX+xRyjm2xZBeDq8yX2P73JiBkn0htqChiUNJqV4kVYYydhFqzORei4+n
7WetlnJtuwmquzHkL+JF1MXF2ci25Wevmtk+8UEVNzQYjQbcXGzao1HrkxyF+uziXbDYGY+J7aqY
vrO2+s/7R2Afl2PFF/TaRJboRP9UTa/lYGBg4ekDlgWgawKjrcdiPj2x5BaAW57loN1pZvKiP2Ts
GCCBpSB2Ow8sJd2yabYVCUlY22Fqsj5fkngxVjT3Y6FlnLVZAjuFko0IwdnpeP1NlvcgcE7zLP/P
fe4Wi3ko8zr2NR90AME7mDUtWLpHIAqULqJ1xTETfdNETYhfDTNyeCukavmezyhDENrP6OjW8i/d
RpzYVbxsTK2ujdlURrCRigkdvUNFDa+ApmbRjGRyn4Q/0rP1GUYZ/enqXnQHpga+CNZj5eecHh5j
t5XLn5pTu4+OFa4YZ6kvxTKvS2/vC3NXSYFMiyQ9/+lY/HrqeJfRk7RY8BB7b29E5kt3fDj6lWfV
TS2qlGao1BMPRDfWMMIWX7/mReiBTJ6xROGCXdjqQMNsp0OAxa10uIqqAr9C1qV6aiw2/ro/J3w+
ARDnC7weizWYgafak8iRSUWwIOit6jnSZnCU2huswVVcxLQOU53RKsfNpcflb+KgjQ1rfp3hC4kE
jup0y408z7hWh/mCAJXh7CWfQ2aU/IGwCE/hNLg02wVSIYefKhXd43i+BR7TVGcBlR0tVef9q0K/
qiGaJx/eCWzvP3u0uLNr66IPGHIfbCLM8Whod3XH0kegP1cmZ/wCmfoIoXJGZUG83sRO1HDWkPLe
dTPS6LF8rryP/5c+AO05WWiyXKvH4eURdPdqL1aXSuzPHMHbnp8VtjPIKFKjBlTzeg+Ira67AYAp
F5okyULFL9y/ojMO9bqvjWVipYsFZ0MqN537/uQs01SRaPBqjelUkF5TXVppCZ/8t7Brfz9n0P7P
nVRZYfxDjbyW9yGyIeqS478RUdr486U+V4oazPzkNB/khSa5hNEBDWL6bmwGM5OrOILGC6Xfjaqx
8WU4lnh3LGFgG9DsVcy6AiV4HKcqmrZngW2tWXzVkaeuwR/E7GDUnmbtSOoxw6nggu/Xy3X3Zx7/
ZuT9iBtNVYrgTQSeAjtyJD+eYvxWSjyNhYBrmGKJRisWA9Qd5idEUsTR3O8b3hCPVHTfpdld+Beu
QwpRqdh6wY7l+xU7CmVn9t6rmIsDDZW0/SNQ9XMCIzozR4Z+/SyQcvTHdWIAnyiA8FEOgq6OUHvC
bUqy+R8p1pPutM0H37IGNBvrxvY+fzD7IdS1GVpzSOQP9piMEPOTeJJBmbMCj1f+2OlJHnf+/gzE
WTKvAUIU24KHiOtSumeSaB6t3dOBjhDk+4XE3FZiChClos2p34cu3AgxVXVb5nJ+V7E95QXfWV57
Ybrbg1qHy5b3OfT+9aZQewICF3QCUnv6pmOHjcI7DlzzB959byO3WlP3EWFzNctVYOxfJ4GqtNJB
XvPAjL7j2Crs3SuW646+GP9zF4ilVSaba7TXE1dkkL+V2qClSEkPaT9hX7ASg5Syii+807mUoeTI
46Pko3pPrC7P0ifAOPgYGK/RFSqy49SKVi3UwF00snJoYTEtag/3kMVahLhE7tvHiPiXy8SCfu1N
iGbxeEq1eW3yvIpsUElv06mfHd7cdwqJoOiI4hyzG0SwXoHC6Y+nyiCNcqiM5vwbHbEKRdhsOrzH
UfOogeBI1PZ5m6FtEEsgHfXUrpczTQX0trHZ8aWNBtvLigFQCydhZiR7tbB7wbFzKAW7SOL4NKC9
LzZ0Ra9rdu6smgX6pmFovrhI6ygthEyN6n/2PetKqusgGzHqPM2461ftW6/8Ia/A/RJStkcl4MJM
bhVxX+R1BSiAaHXZRQ0wBBJDflo+vMNeoScQ/cyYvciDFk5okir6rcR/ejttN29Ns+a/nONCI9Ol
ZQeRdepezIdp8l2PLbDY+fmummpZa9YvOtdebd/xwBdF/SfIJOFVo2v7ot++X9LQ+zI2Y3QlYxub
+621+dC24i6haB0gI4c22DoveB9wBhjlfiSN8gBfv6ow6xufWYcn4Mfj4DKjtxUhwci0+DzJWD2u
SxMYz69Ivs0Y/YmxJxgrP6F1R70Y9NT2K0Z+oZn2dOf6QzNqy8ILrr83Sd513rlqixZNEUCK5xbZ
LbdRfVukEHDe9U30EC65H8rCbTZJ54Mt9sXIKWDczCT/HC2HSaCCTLYzPS6V38cHu+1U7rCozp/0
X9Wl4mpKNMmyfhM2xdWSaczZ0pvcEEE7aX7GfkyttYgZfbihOOEPbZAIuAEY3UEOnAv/kCIlSPAu
kERkNGNr3dabe1S4yngjXv2dUwqH5V6RRf8na2d+di+OBVkQ2FCpR8ktWoh8iD8gqtsxHy+Py23b
Tp9PHD1w96HngdgKaz0/ZjNpy+Jk7T1NTVZrZcUdrgzpf0n7RWDDW7MWMIvRnahvUjU/o4ZA31bo
oW0bmPsHGT3XElaenPByRzQBGNdL+l/jaBd5GCtLmlscPAGKRzb4OBArsIlKRAmWyKsIljo3Y0W9
BNQOf2wsM3bWwvtLgWC7dvlZw8v3M+jmprGGTlfIsuiaSXX3kyuAM+1Dyj9tYdKQcFzA5BHin2qb
6Nbwtlb6Tt7pn5iGURYpr2hL0/RC4R5JBOaN9XOnM6F2GHHatHj0+tsx+gYmOvk2lMU9XzXPMgjD
Y4npE4JY+dBlCOSwMIYqFwhJS/IRi3kQQbegisscPdyrxfpUrmNgRfRHSQvg/zThxvTuiiR5CYix
5T+KlpOM8jw3osm7rXS0z4hU82FqSGccB94JCERBeKyRUcf/b3cCoY21HnB76GuYV9zqOJCntygY
mLudG/GrUyBiP94iLyh3gx1+MN2cgI/2fbzfldwc7x3bNiWPWv8U9HYWoMAUBRGL2R7NVwU0NTgI
8gRm0Mx2fX9W9G/utQHEagutTIv1pTJvbTfX6avSc7R9iBfQZ4DaXYScMi9y2FfWpnDFumn6NIMZ
sQFklMaAsSOolKrTtS1XEPH0gdUvVbtwRtmMFWVFsieqlEV2ni98z+p2QuVNoHcJgBMjt2xgXSiI
AjMIsOAJtJVvBFqll0FdOk9wN1hk4UJK2Rqo9m8O/swaY6+S+IruSHQeuIKZr8eDTEXolptKL9yN
JtZtJs9cHLKXXbNwYsJf6mgQybx8E1AqcrBfUiuY0lG3XhO9zyipGoYkyaEkVj+VWrDB2sb/5JhQ
VJnfDfxNbBw+UAqA/zQa6oW2Wi4VTBmYP2IYtFpovOERujkUnOYScMNcG5h+N0h5JB2styvvTgea
N2w17enbsbU3VHbs8bjBr5Vo/ulCKJVevwfST6fYlpW311S6QD/Z+4kPm2YCJ76ExM6r9OHD5RZI
Icr4nXYhlou1klYsay4N7PHNQQDMvkAWiHJkTgwt0O5mBbmPK7TqP7WOYKj8gSz6l9PaCFUewUPI
r8AR7M7JC95wcfUHfpdo9nXscgYPpy8PA1eVGvB0XeJ/U7xLpMCag59VsYSe1PFWiRo9CkwAe1lX
qUawHNxQUOuzYmmr+k7kwS0bWjiTmNHiulidts69iMtI9ohvWIClPsSq1HRFjt5qblSIJl4SSJUd
Q71Js/BHqR7/FNAhYMM7jySGLiH0Hh7s73v1l7DM8X8yvmeBFxtJYXxBX6pNbGL1b48UCalURh5S
M9hKLVYZQpeI00OtNZet5bSvFklca7kZFFtvdZ1+eWKv/AM5uyl18uYvPoqGFoSjXqsG7FvEe1di
0Xlt9ng53BGI0fyL0gwHB852K4cFZz3Soz69exYtAL4Gws7i2e9y+DQFVet3z9s/BKi9ZZI2S1WL
DR24D2jon+okn0NjFDE8zV9/FHZgMX/0CEU9KiJu2l/3NnAdZDqcdzhnaUb3HJPpUmRC9c8vUwPE
indB+CbW72zgGV4RmvIAdfrw3hISkDUs0o4U6+jpQpZT7kbp2eh1rG1R8Tml4cSUxHc6na8cKEh8
STgOWuhO0sbPW72/QeyQIk11GjB3fSLarJd+V15LEp5aqzRwRMX5zq9Dl3SlNvitSfQLbyvKW4Zz
KI61k0hkBU1VGAFdlbxFMEV7d2xMKZwDnels5NQ1E5PkA/HfzPb+CnQ+CmfFVm0vOGR/8uHmapKc
vgWmbpbVY9Qrew7MoIX3QglcYF4ErTyrxQz7CNacyNS4YZW4hgo3QuAZ91Z9IpLBSPWB0U0fGSLu
joXmwxqwwk8m34W8LaupWAQ2NocR4mWpCnm0ASI9sjVHsPqs77JJtVs2yHKG4ao1DUktNwKeBIr4
blSN4hxWCspYHZxskKUZ7ReWrYH+LBh3oa4cemBJyPIcwE8ss6qW9UYtX4xrfOsuooElJCdNDwj6
uB5qd55tPcIcL8U39kfx+AxzIheYW5c/9e/TvD5QahTzM6MwpM62XdthYKnE1G0/JFiDE0bvXuUY
ZEwXvJIr76yfTulm3baRSsj4D5r1IzrYUEeeIU9UJWeb1hjUq4SraLTqJJapZ0MbZjRptb6xC+DW
95pP6uRcWJSHW9etERg/FlXb73wJP0//f1vOuDCvSHbpg+QHzTZL1N38OY0tmhHpsJWLUR54nZ9Z
3hDfwjFqjFBApAGF5M2tGnUd/W+7kVVHtO2eqUug8E2EcJl6LjZ3tMoh0pp52JZ5hXiapO+5FkTW
nD1IkzU4ElZDZT6wE5CXiaGMTQqQkNNBED97UaVCodWPc5vJlc8vfGr/x/rKKIMC0mLbQhdbM69S
LjAZNHc12mMH2lV8LX3IJrbKHFpTtcyT1vgUpt+Hj6KrO/t9an64Piz/k4NQWR7nN2Tt3zL6EsBW
MhA+Wq6sHR9kNafu5TPGaFjnE/Zp7H12CTJw1i+BsPjc7eGSkUrH6WM7EVXI1xGIZU0yftncATBg
D9VrmWoLXaHGA6cvY1N55gDA87jI1CoxZ1NgnpDjK2Kz28JXigtWgLcoJ+pdj2gbWqBV96t2W6n7
n1aJH88BW3dnDka2Y8mcayKGf/H+WVULO0tPh8c3ZVTxQ9wJvBWMdT0EXUe5+2vd+/5T+wFIAwA8
vEWh/Sqsb3Nyp8jrAFK8tncWTqU4V82GBx+boaD4OHKTUuBHWfI1rjCmT2tE2Jqv8PR+sQ8hkaYF
Y948hPCV2o/o/1qFXK4lcAfNdG+5oOaRwRtOwtjWaobXxLHLpQiP0ypxCRdsDLb57DjOoQGVxIP/
ml1aqBKt6V2bghs/H6AREC06iV42s+ctferwCtjbF9AiDhrw1S8VoIifj6M7Qmg3OQUWR77OHiw8
YydF96dLYqmB3IZTBvNnJFHaFNOFE/HFyJdIMPZQMB2Rjhu5FW4Lm5apsONq3+Sa2FdJeZ11idA+
BmPY/vlBuC4N+pvmkEEj/SGxY2nSJvX4ZnyIz97jegzl4BYd6AsEufoquiYCsCtYeSv5XYpUJ1Qh
niAwFb7DbVwBnecytJiBg3HhyilfhptY++86sjtrWiYsRPDy3fPwb5lJsDY59482B9G1ePy4J6LF
k8iqcujlXHebHFXlcEQl9/R8xH4gnDZ8je8MvxK+VoDuT5oSHQhmCNiCWlMrQWrWga/aByYmRIe2
lkZut/lhn2Eo2qdd5suWNJaOpVrKWe0eu11RCXMxxp19SxMrk+MOOVOaSUj89ol9CC8C2fOVch1X
w2YYBTX5FvM5ahRtwTjQxtU9ox+K7FTFuSwestaywgxRiPV40CyBzn6i4zWXVdVEwobNT/IAYmTV
1P4XIjqQCZHNeYRqhuTv8+ksjUU6JDxixqRhMUyEyyWN07EDaAwUJyPJUxUZdDPH0Y+J3J9k85ev
EGwFaM8mk9Zy9ysVsX1cCevVdZQXXoi+G9fXV1wpF4NV6MbNla3Nt0GaIJH/I/FTNWXds/fCS1ec
aMejA0O2atpfM5g01cOtwMjeQi220cLjoiIZn+Nc5CxT0VDa7YJJ/lv+6B7swG1zxCqu4QVfJEod
e4tlZS7UW7bS/XzC4WQvE0cY4y3y887q9T9p+dcoL5cI4wdSsGWu25r6iqcl5RsxfVPO8EODVsRd
1yiXz6O84VVO9vlZlUVxjqqZuOsCqj4a02kFrOHqV9ePfXU2ayRvqvOrrF4N/TXc0lSK8kdND5mo
kjBbJBXcc+h8ovTS6EAr6vq5CZhaZKKzeLfCb8SsAGxt7lZC2Y7QekODFaHKOQ9tLcTyMBGulQU1
iosC/86yF9p2IyjCeLHFdvaB+zNKYN+p5kvCXkLr9IX5ZwVKP88FsQ1a/GTKcxHeSRp93xfQ7qfd
kifFbLXN9B5HBeaB2CjblZkjyfuImELXhSwWW+SRXy43bycfkIkdBwYQN5N5yZlVr0E0eRPszT4q
5KlJGFKZ8opf6p/Jc7Op0LOLp1dr3itaTEgAqAWOYnAUI8BC5c8Ej92gRPsT3i+0+TW5C0gSa6re
Lhyy8BPKPeztCKTkpu145LFXnV68PaQC0wIN7FKE7+Ra2hZMK+14liqnHbe74bIcTiEdXvaXboQa
3Ksnt5pQa/k9rwAw+kiOnwroLk2rWaFjw3zfR7wOe5SI0Y2SWszC/qmJMv9gl/S6K0YWmFCGbrdk
DaCHejbwNUO/D7WqwyiKj8z6KgXpsakyalz3MW66Y9yDil/9dyXGklwI+VS1KwS3/e1HcTKRZSmF
zeQC0bMRd3POTQjK6DwEmVRRd0hoUNbEvJizqzC+aUmvwPE3Qd0ynJ2zMePfKz+t/AGwLPOeURq2
urLiE06fe0MqZJYlXZHs836YeuBRJs/NGuqxvnpWAjFQODj2scy+F3hu9ZanmBwpCtzDbS0Uf3Sr
y6fQnOGgtlRXgfyszFYa/F2yh64+z0DTprP5dEh7KKMRjJv4Q714PeWVTWBmTd21NXTha+8mvssQ
llwDKwfIeb+G8jvcRxJ8ofGxvw86Q705UmY31zoI2+3bTppIuK+gnOopWf54uR3x+ds1MKC95Q21
hLEGzsBJMPKMHcjMA/Fjz+Br4S8jhcjgAiT7DTlmN7l+rcVOlKHCoz+oJ9bJ2brkgtzimIH3UOUp
2wiothSy6/enUYprmigFdZJYSu5qW8dkUe4i2epHNbBPNBgknt6B+xAJkXIFnFCkxnfXw6ybA7Ry
yxclu19HK2qFVE0dsbU/e82QXFXCBIkefhJbn+RMoIEAyouEdnx+Ud2c3I4oj9ru9cvp7G4mYUhL
TYOLD4fEwmbWQBKPzN/C83vPCNwZKrD106K6vNQPTTEnOBVB1xXUBfjVTMYqqzS8kKi91jBTC7TN
chAQRNrAqBsGhXYdvVem1Zbg2Rcb9sZ6wNjnjRYwgzMFHCxVCEu0+c88EZUxwxcRDR4Ru3rR0AGX
vvvJSLosEc4UEF1x4iFVBv+lFPbuZvvYqWtRnYfGeJ/uZS7lO6MUeWdnRRc29+6o8/VbQw4UuYa1
E5DQN+SZUvc7KlkAWa6AmSomReWU+Vv9PO6OyVaZTV36RkL6V/qu+pA/yxrKp6dKAKQn9u8h+crP
X/u1RVHriu/f8h+Z0goZ0/ofyL8bkUDLOJD9TaTUCP4kRFJX8QWTy8nT+1jPj7H/ilJlcqrHABgz
L4+b39rfMwk1KdN/6XuOWDj+CBwD7q1leQPbkt52xjSXz+O1oUp33TSUozeZ7DE3KTwMuEtuiSsj
e1SkPtvCYnvGpCK6VU06aebY4fJGnO5/U/bxNLt+mDR4MKHR3+vm0GC1VyP8YLTajuV5n/sJnp2q
L6ZNIrk0Cu8+zAFkSoN2H9F+ygOiT3Zqf3MtPkQ2W8uf9Wkh3whCx5Xh5DYrDNvxZaMSGwEhFqv5
yS/N+l89xU/NynYp+BbxGK+bkywIwOeSFZUhJAOV0yIs2cJco5DA41tegvSR2sNEINcI64O8rMiW
PZ7+kmBUwT793kWh/MeG2n2QSMltZ1z71Wn/5rzUDUYw5G7voZfQor6juK7NBz+7ung2AT1eb1SN
voxZkIIMloZZpwHAzeQWEa6ssCqsWI4qRX98NvocMTYpWfXmundtcqF4rX3LRGGmPidW8Y3IbEur
awItl0+LxbhZwdJY3E7K2mAcbDpWip54fp+i/jnSBQMabDvIe/uTGtLTSBKglJ0SuiiUpRVEzDpg
z1Fn2T8ml7m4peHeAwX6Xj7AT+oNN7FP4FAtz0iWxDCOqveR70JY3Cg1709uEuQ/kCeU8joZl6Vx
NK8elYl/FzZf6fpGYIs6L/BozzM2TpFEBYP0tb8xEoEFIbUmrvhNWstSSBXH3zmTRzyafJDKXNrT
oou264GphscvFXWY6uB2Tj017X4ORYf3RRGBlu9RNaug/rvEFgDJqj1zxzvFV5RBJ2rAySyNBzjh
2TN0kPRI7mK0Yr0qmrSWU+kthSMpV+uqtnK5+8WZ5cMTESzUEMx6ecXBBc062GuJ524eUfj4s69U
kRHZySSYaEeLdqHgCaNe3zIkDS09yKhxlued9uRPnoNrxd8IRTJjM9JFS/o4YmJWG7LM0YIkeQH4
eSJeiyloBH1+eKXvHSwmeWS0Tx/h0rZOIzLc9YgoBGNuMJ/3v39S0d7jykjeSZcufuT87/0VRJiT
igxz7y6bdeDUOErkSkQ1/DjJym7TWZ/jCUnYd0C26lZJAdBh72xPqwYPG9Obht1xiTXizKue9IZ7
XwxzXt57QxI85RrTTg6CpqRdmiv2qU/5Z9n5fHueXYEHqOA9NtNmdLA+tQluyh2+rbhaJY2mVK+g
MM2yK1fsoDrH7aWcw38saHsdDuBY/+wuuZ7AePBloYLk542Dvt1ipLLWa072iTRIUKHPGVhcelBl
ccOCEni6ZnFErwfT27zlF8MX5N+zC3aaceNtUoV1N/q9dplmkxWCzJK1GDVeN0eAFtGTMDjpA9vN
TMz/Pw5q0Z1Ef6dzOtKAERw1rBHHpAmtzvm32RL/olKCj9BcrHu5plTlPvN0yRKYJD7K8ED/H0tz
Fzy8vl1nqhBSFXR4GUPjMdxBSCchAIS4U5vHasRsSUPxhkT/DIAEivASfBjeH1VhjQufmGmHCvMY
ASaKMKCuiN9dwJN/kgvmeBzJYkyPKDCnSr/JzSz4Hz0PCEgIwPwUX2xkzBKPV3BaIFXBuOyFPPNX
O2donqatk3uNSN3q/Losr+9N2fQOCpr071DC3YLUfMIPYo95AMRH1kBARmReS1DEBZFyTyBVOi7r
NIhHfBWvKwEEULwPtqrAKGXceAXdSKwB1Rr9gJpZk88r2JQ9vlOn38M3xv8g8qL4M4fFuUhPYfoV
TmdcvTzCGxrnup6CWQXnc2fUsHwtSG3zgpWidCQDOhK97tRI2RJhDTuKJ/sZ2OCnSdMueHzt69vC
zN8LfFwVUIeLay7uQjDnAlmmc9H5SOLlGPqIf1bfSn8N3S6GHfHk9wZdM9arbbF4avXCt0IMHujt
SzmUaNGcuGFkNJO4uA5N3gPwPA1tm04LdC3a5g5yFP7VX8FUSQbfeKJo0/R8Wjnp8GKuDTaYyFpQ
sOQ7S2daKz6KTE3VRkcV+cF5nLy89zFMgsdEgi2mvs1T2ENyyDoIaUGrKMYmDjuTW3G3nVzwMRda
6Wm/D4SVHuGSTDkG6/yrLFOVB+NudVZn//o2vhqVKpUVQNGpXCIw349RTRUMruCEMIlrdvIwL1E6
ff7pJJUhRYLMnP2YLSxIMLzQ47GfreH4wGq8zeDQjA77+k+M7BRHPDbbaaJl6m2D2EoXGkd1+/nF
T9M3GAmUvzwKQHlq31cAb6p4e/DtQFpRx54vfjNmU8aSzsJ4KpgzwB6MW+eFtK3erjwz9GbloCW9
gxqQTK3rIz0QbdlacNBQhO72geHCXKN5+i6MKuXgn9JMNriT8YEQOwUy6kWqtbQrZ2Jv4Ics6leH
5QmV2tWVkcUMT4USgUAsjlmMXW7mDZjv8ZUpJV7jeLWChtsLyAEss6PoSXzDpwRBVNMpqaqEtEtO
MprxsfOGlif3NVBNZI9JgbFXQXWX4CEQ6+uSVg8hkJwAyvD5/ZsRn9WSwMbJkWkyeB4pEe/eN6mh
SuwmsOvE6e9E1p3b6ZQdLC3SP0MDb1wIRaQnP7Kr+tcnwgMLXPp/pJ/YdNVQvXsU32skBGmGbqHn
tTaZ29mCm+lqkkTvHBVIG8/OpDqrBEUeQ5c4H0B8/SOmjQP2jhdp0a+jcMZ1XSaBIK1a0rUoLoOn
mSSMGprGh9rJgIbU92BIYd4N/F7EbxZWZpMtrXxqwSWn3OiqRQmBq/3d18kGDN8eCA9n7eU1Rfz3
a8FyHMcYedAvWTt6qdPoicTWDseX3uKI3Wkc7M6trHGvr/PALSrMVUhPLy1Y6wcMjcAnp/jz9Yl0
gqXvRJRse3uB1gzPusdgieUjvVVJMzq1PSdnZMkfZgWn50VoSpuOhnrcH8cMDDPOfgBkRImKYL8I
ZPjAaK8qGnLvTYWVXhImr8Pq4sorNCsTFADBG7ZghcEDcxrvtEAHNJsa/dl/IC2Vwy89FqnRNGpk
n8ZVFfwqjzFSxg0toWJTMNM2I2vvvS1o9n5NWhjLO/YboQudV+55yQhczuL5E0HbA1iQ7hDmosYt
Kch/gklkR24h1f69itZXFq/P6DgjjxijDnZPUVqNHcerKjupfa2eHETYgzQcluwy4QyT5H2kYKg6
gNdQ5eVSj3eP2L89+60/PMWizRXdhRTY0V9ntxQo2KWa4DwkahXXluXYFQgqk7nXC0bl8Bif7aVN
22UXsc76h+GMOV5A4Boi59zwU1D8qpZW7Lh6rqj0auvoDGHHlU40dP0H2BqB/Zl0Whk/ncmCwHiY
BlkWXkQCA1EZ5g2G1Zkt1Asa3/yRssirXYV5ONVdFlBodMVjNMHDsqt6jmCSp5rENWz6xser14J/
XxjiiWYhg3cq1PP5FI+0EWVYZuqZwOj5dTCPjOy4kZ9J3pBaopswY73o4ZT6PzR9QERbutbiBPt/
wrFaxkjwxaqdd7yDlYMg7Z9arI+jUUcgxBftzD8InRUy1A93Xj/kKbkCnFrVmvlV9uSE1zL8DlWP
x105HEJrJ7MBwqLVMCHTN52gOtbygpvf9dVttc+r4PqWaZSYMgjwPg/mE2dTD1jfWpiJkALB0FBv
bVHlOe+0ojJByyU2J9zarcoVG/pTcfcakYnJYwDdKDsS95iFo41jmgrzTQo/4oKs4OgaIO7RvrY5
FsETasmE/yQXgXw37EQriUfhduOyOpaIiBKwGmtgJ0WVRBrw5PczxhDLQO746PVj4zv1FDBy7upy
sQo83+M9Lf7q1WtHhaP9Xr/csIiXXdQC7gypPs9IpMOak5jP2tkzqqyOUog8ekPx0ybzh44jCHQF
3qTINiW3pAp3QZNLPDkB/1tOnRBO0TRLScE+yAtiKQ468r98kll9QvNl3DGFYa+kWstMFmV8UH0C
4Zs8wqfmNEef66y1aEptp/h3gC3hNV63ERSiYmQkNn4Zlghep+u3ehA8W+RqkK4dJyV23wpEkHh6
u9MlsVOnNXtYakXt/Xr1a2R2/CLe7uTBXh2sK0X51TippyJtfCNotb8Ege2EDGzPUR+LZ3n+QIsw
QqYvOVnl2u+UIEYKe5yTm2QKXOUZeRvFkzGU5tcz3GiO14tMe3H6mHqogeVdU6h9B4mP7a0iD88/
9plj/MNNLqvVj6H71oOwWFXhmfsRQRsdoiBfaTrCGmWaH6Xa1+cMdN+qNrP4HVBc6VD2srKtQJTW
Ww8LLhWiSyQzRpENNz7yN7kkm/Y53GTSh1zXom2SdPg0nlO8r2Afh2xl176pdd5LnltQlqiKKQO1
TzaIpaEIfYbqQ377ow/OszDNCjtNxqD6tkBGvwl0W4DibgKG8y4Ubku1dF+brzL4CBx6GUKLwzKF
L7HxiGhd6uv2HTCg1n5Z6IhQvJUx/jEU7bzJnQmHSUcM2+IUUnUKcryGkIoqTuhuhO5USRSDI8Ez
a3rJp/5R0MzqugvbEDKXtmk46eR5PUfBB8nzlODprBVaN5YTRRaIW2UXnVtbVD52lJwdLeoWTDo2
bUHY7EXfNYpaUbh4/+jFSAnwHHVVRwHv4kJ3DYm/geqXxY3cuczAt12//zGM27ihzOsVfILhhzII
SoAmWt0zVCiQJg6C0PvBF2ti4hMFld0Rf/bP2PbPH2v+Q/SHzD1rqAALSeTb/oVPqXTZSyLmQ6id
xU+a5IYjy/OFpnXk7Sxo0ZPFW9OA+66vg4o9miYd0VSOAGT8sXts1P3r1J1S+Y9H2q6rH2wUJKiR
va/F9I3PPgwAHlMaMNIvR6h8WIA7FfoayQ9yH1HyQsERNoNbcMpRSOS9u7nV/r2YS4Dd/eXqLbBL
Bi57WXtw0Le/IJa3gSaZP23VR15BXzePKO/D8Wi6FuTZ3p6PDxH38B6ApLUvufR1RGyOh1i4/frg
CF/ARAaZCvx+2DomsaBE1QGrZQFjXDRlm40j7Fv0ucOadvagc4rcFFFXfNKV0sTELCTwfm0iw4Gy
UMaCNX2lcYsb4H5MjbF3b04+PyssKvwnmWOvrUXQburUsTYTNRNgy5HLxIvA7JYHi7JxS/gNiiCV
nXfUJV1vJ4EsBTHV5T8/Sq1TEg4xZipx94YvYuoYBcXshsysJbIN47rrOjk4MaiinPxKWaKSOCdt
mo38+VGR0XatSaRX+B769E0k40DWaN8fXIt8kvoJGrgddK8hls1wKaARkeRMZZmiTcOGMsN7zJP9
Y3WgdUSyCqVBOO1YakKK4cnrIj5pxMALxFVzN9EXPlNRNgBRkdoXXsZbraNfthCrdVRBbo26ggGJ
WsAprxOqnAekT9l+c3NYW1kO31v6YsnCnT6dpU462mgMPfFvs3zLptMTbX8O0gaMT9e3uv/dPTRf
ET8UK/pNBnB6iKg86E+jFREfUZJF+69bAnuAvdbErCETt+i0TOtQL2nC+GTl3GYLuseQzjcYD8QG
+/tsXM72l1a/Dn/aR+X3YoG1GYu2wTaAibt8JJo4PtoICWwmO7k5QbxuZ4WBM28sy5y62tJI0Q9c
IvgMaPAcma1lcLEvSYPw4cDm+dcu3hQj8Gakg9APdkBnuYWnUiEirbKyvotgK/5TKTVvJ6y97mho
F9F51g0LttBHlnWxV8DUq7FypZatmwcMv5fmuIeFl0QVtT1IyWVRdfsqbcFKy8OjA/YyJkMoBcr9
5FkGejsePNwOmVmpODwbsPfji2Np4UaA9E1/rCywRLB3huulcdfKSeAmiArYeaz2YjjEDD6miIHG
1TG+yNl2zYj9ix4A4Qyoi9shVmRL2nPZs4ICsqxOSxWTYauhe7nbZQczJs5ClED7oDI0HdWQDEFV
7sBp8Q6ZceB1JxrOwDbyBwOZHOVgiYkM0GXHn49jIQ05zTb7Bym1HrkHmSPmHmUjvwOvmOxF5B8G
ZbMXU8TF2kjtJ5XVWDXW3Nb1EErIzh4psz9ZnBnAvisZ8PbMXAH06L+8gueSGoeof75lTQRqCYP0
poHWVmres6YZHcSc/Ll4hJmO9O0xNsc248twnSTYZG7w6eMIFysboiTN6DuEptk38Y+N3ZhQz7v7
XzQ63vuFsQN8Xa2mDO+jHpF7S/5HsJyxjF/P7swDCj2fe/n8scJ2D4quEyVBEamZuUGnFguK1uOV
dKerz4Jln6Yfy8mSX5nsReOj5Y1WiyAIqCs3lddXV6oosHjpQZqs+d6RUZwKlhR3TamilT6G+btf
JB8ZKHTtZ2tE9n1qMZ1JYgxTrOnkEmEkep+qblOQYSATYcpOauv1chcxYCqlmu2QQmQW0BXLLbnw
cuAXEXGkTQc5VRjfwvgYS3dHDS6czNfXUxSCS1EhE0FyTONnTKu1xBMlpUJozzzTp/6anwsPEPYt
rTq4OaxlNxieXzWdaJQhSSE/kEFptLRpJVuI8yHHIvAPJ8ToafxFj7+zgLYv+HiQu+GwMmKD4581
RipyiYCdbuv3Wxi2EY9wI+IFyvwtOZxEyqLQQAyRIid7tICOLsn/xRsloDlzLTp3sM+HGr6V/Vl+
y5FDBL8wib35S6/5TtoFhP1RHyAkCFkpowG3HBFyMKYjlDfrVb1lgHJNc0MA/CSXzA3n47sibIoT
NQXsVhNpEm2JuvY7csT/7pvtj71C5+6ZuveoGJexOqHxgacdwVtWGQlXqgyQIVg7bZQt0K+o7KXd
y9X3HF8FqWIZAopKQfhMgKpUP+M+rulUfo36CQk0qMrPJRk5+XOwlf2hyzmHL6CtYTKk7UjqMSYy
CYOwoCzS7CMNHpdfNFasITEuy4vGsKBFkVl7Zf/C14GaskhjK0dti3U2Uj0pxclS9ibYfgvr9NOQ
LycmD3zkBk97XE+QwnxG8eIfN3dLKiHl8KrEjLVJq7n5v36NKN6gaXOvM9zbo1dSL69bOiE+Rkfj
WOgkcQzfXiO7ThdeI2neZJpRwJMAGGMb+X2WxOKisccrEVPB8je9t31O+BYo3cBKRUH1I2udTZaq
aST2c1R//zbcPUJzuNkl5zw2U+nX2gEzO656ZMDV4nDHtZx6ryN7y0ANKoq0aH1ge+WUe6HAk7JH
Hh8MaMMcW4kl6n/Vk4/J4tDr8serO89QwGuSFDmMavraLRk6R/QAZSdTtC9Xl8nUk9K+5ry7mmWx
nTfpKmcKVZpQAXccdRDmRYnf/w5Rjmtu7SjCsXdkifd7XmXR84v1zJPcH6ODX0h9tmL179MCW0OI
BmGeIT8AKiLfMtFucE/AqiXJbIyC6s7fJUm1cwRP/br+CVfy1VC5cMl7ljnPwdSXdnG9x8hjthUU
RxZuWbvpT7c0KOS+2GW1pUECcwn9S4yFkEgxUPQzHedB64eYMpojkWwBwBZa15rWj5uyzk1U30IZ
jvWI+j702RKXQbTAxTXlBMW1XF0YluK3ZcEIaKaBcXizYoM8TnXqavHSkbK/PkOz8AL8Bzqpx0JD
1aPEqG2XFNagy2kDLElp5VuDvXKkYl0v59DFBepBmGFMJ9ipwoywvifWsfDErMY0mXXAZLSG2Rhm
0odugoEFzf+CuqXeS1dneMc+6RcSCITSPxACjdcpmqrYWfh1e6p77/MMOPAw7z8UpERrzo506+XU
Y9Bu7dgUk8n58paFuFIK5GbPKQErFb7W6NQCz2KuvWv/724Twexl8MbiF0tD9tzvEzvdbW6ioD4Y
92Z7T4LhiUZ2oLHtuvMm2G2c7yKUw8D0DLYf1X3VHbLG31B4X/YLNjSVgG7E4RIIdmVpo7ZnEz0d
ujptjMjuYBaaGxF/0tL4NPR9sbEmV4JuK/kwVqhtJQ5UA8789xPBHM04KOaneZU5F9T83jdY8hqW
i27aAKCuYdd7IfIS7u5BMkUtFz9SsNvFIKCLX69aeDypaGWZzO02ywVmMHLi/Lk9Lru03u/xFvCo
/31Xwvy1vhkYbqYg1FXOjcD0LRCXhe4vkTINscQP5UqWRbPxgz8nb2ls13IIXB3HOYSMqn7EXyP5
+gBo2A+KCvJYwB8aWDwCL/BQfAj2ZmcHeiaOtnPehA0BuXMSbUgCDGjtk9AmoSErMPlmGTIc0Xo0
n5Up9Ky/cclZEqwMXlDT3Li2bSnyondNYpqWBFvCTLF84tR5NR/kuXFtdUqIJLXThxZr0PPFGqei
xu/ecgrgbQc6h3SF4grk098rLqpCqN9B76HXoQ55zaQsMP2QV2ZO/B6ZqxwT7CCl54ZXY1wd92/S
3M5Cgy8q1dzaOZoVVhU9Ydj5GKrD2p40zp3M7ySzEpGOadcsYyDpRvOUh7w1ihgi6yh0MElq+0mc
p0kyRK52sshVe38AQxTE0TgIWosG0K2Q3WQA+QRpQJc6IHjoQe2cJ0cLL2qnrguttAlRCkx+1JYi
LocAewCM7GFbEqz4T6Z3k7Ax6eMBv5UBugG/N55WWS6KL+C5x22dYFpNocm5n7D+MmN0KUJcdfnK
p6PD9i1GncNRvSlhEWZBDuaAhxdsA5OPqOE5eHbyct55gRuUgOLxk9Z5hLXrMCA/N4ZZ4E3slhCQ
AxvSJFrzCuwcOmbP5+cLn2wkVCOdw6ymXwla6049F8JJpxUiUADPJdzq4y5GpnBSnzKQ06tLDp32
iOT49xyIgQ2tqZJUhOkAY2VSnvTntItRyBl5kaPFwmuqtS26W+fesuTk0WrDoAhKYcJLLGdHANE/
mTpfGJLlsLuiubzaPcKN8ktdtjg48E5LFOGSyknWyZbrPTSwlCJIijeJdg1IryMMWjdZmvBVC70x
9djC9jX55em5c1auwZ4egrkukY+DdKjUnheIe80imZ83f/W1lli5Jn5Z8OtjO++/J6CORAeZyJ4v
UYKOtT47uLxdOF+aZ/XOmKbDsvTnd56iZbrUJYBU16Q76wiNa/VS+qH9dTlTBToK3FsaSP/NGPIp
FYfBtG0jp3GAniGXBn6xXDUYYOQQlf7c9/CMy/ZJz0OV+YBjtWBP44lUsE3DTzy2EQkISWJuCySN
7AMg57o8iW+2aHKUFxHhDJJNa62yDi1LigtjldRBat1WmmKCwYX6Jdj8OtZwlLvv3pI1+QfA3pOT
uIZ6ft7kUBwrMDH1Dcla9NgiOcP48OJUbHmbxrF2O/DFO3HkeQuXPUkmbiNVkXUpuqKqlGW5B+Ua
k2CmlGmHhOO4jWnBDuB+dWdJcyvaSOihFYKAu/G7Saz+WN6VYeDuZkvL1eJBm+xDLgQ4hxcrVyGO
F+smJ+/yP1jQHbW2Fm9WDgZFvM2RdcsFIoKoLGzky4+t0ACvTVY3my69yhllDc4pnrlmz1Brmm1N
2PNNjznD4WkHU5znruruRAFeOZtydMw9Vvszpq92hLimVOSMNuea8PsRuxNAG5Ryb3Lnp6zxTjaq
edH996wBszYXGedWIlfQVJA8jKC16rDuA9d/BjvbhKzZ8ZueLyKv3uJoNsPLjz8TuWRBdgqDbrSB
0j3FrOjb+OlRiryWbogKv/R9uOpu3uar2ZVluj+7B/EBO2Ouq9ZZqozJlYCmhJ0VR+iTHwPUzeRm
vE4Xc4QfO8JKSUUqY5WoDbnpftBQv3eFAKJeGHAyjl/PKNzDX46CCPmZxR4aLLD9E5xt9owZEn8S
7FvOclEMG44B2W0MvUT5q3C/bVzo2/HQlzPgx8U+2HzLJnoyuEjyrXCz0OGcWixiKtLZOZ2dw0Ji
Srqe+AF9mtPO4Pu4oZSlgOhiewl7B520CWTwpfgai5c9cQSJvob6rfopgTPr3JXfFLcm2dQnysH+
MJfgKNgUDFeHqSbh+nX+HQ+lGQWgHrYzIqLiQgsblhbOpMR9/abIVfaVnfEmUALdGI1xtphzriyr
e0wHgUjUXgkPrOKzzcEiZSuBW8XRizQ2xccr4R28MQ5jApyT1E2/UGNSv0OXiqohfjF6OIeBLqR/
bqu++0Z1YJI42LE4bTEGBFhdQ82s/xe8FNvkUrHYKK4r9W0LGg5IfqL9xIf7M+VK9pojGQ8mDEgG
JieNbLR6cppgrAK9dzcEwRMxZ+gpW5HhHU5kvR4cHyjmhrs38mU/QYOZRZa5fDHHPbhIAeVQLE/i
XYjE93SkwVhP0I6UV3ne5fDSBgELa6budhyR1IcfPBJcMQxAqiUBxLGBEh8kIqEIrLKOvVOPnlhU
pNHc81/D08e13XPUc51m6EO88ZYb7CS0hta56HlOVEK1z13456w63CRe/seJk+indf8DPbcqaqHu
I6fsVh94vdVWOSo4ydA++aANWD5Ijw0g+j9zpZBIcYUNF5jjSwapbsfnTg08+u1nXEdeq4wjXili
5pjaH5navH34H6iAf5cbTQ9lcpbnYt4W25j4vMlICnvYSy3NEi1Ar47mZf8SgEBW3Pny8l4+VYvh
psmX55W0jDpOdBeMhhQGK9mfeYilTzA9h75vrClndYs2mceVlk/N5Mz6TiWxSN9q4WceDoRrGOup
eVxz4/fonOKff81vfW7pyJxPibjNyeSo78Wuh1utZ71Vy257WGRD99zs1vi9/9aqCtE5d5ZLv5/L
x5TR7t2Gxg/O1/aEgb3KyR1IatdOobCitDMAGR0Bahm2AKKrQwgHgqhTeMeY2THVE+Q1sd/j4q6X
IbwAm9rtND0Psg9UU3yKcoMRaBm+wYnQpgMfP6SOdi6sKyez9k9bNdLUm9iVWCEMicQO38zo05Mq
72M4Z0Jg80TVlQ3pUGwFarENjcV6G5ZR1SviOrNBJewgINu0P5VNuJSzSYRIsken61IgO3uKFvBG
UjbdIPZZDDjII9yfoD7dUpE6///w5ymMsqmKPPf6Tslxl/LPhOCfkViwguZd8Q2TB/8B4Ze+xzft
BiQkD7gpeHN0tOC35bPKhG27uFEYS/6pzRgtGjXTHbt4OO9UmxGPVzjYNPw101kluf0M3r/gbUaR
MF3u0JcIWkPFct418m9OQfLld+KSHmoeQgQ5a2w2hRxEIW0dqt0L6ip4n2yuo5kgDtR1ehy4ayyt
26eyA7OTqXnyQq4YZdjd0VnS1ZSDO3yAcKhhpa7Z+6cILX/PeUbHGrvydwAuqh/9WXMCjK+ktFOZ
MnYmkSAk9OHvQHUqm7CbXQy22aR7qyiIzE/7l2jYWUI+FQxfVTi9FgA4Z3tdwHr4+YDElqMqaZ6g
N6Fygqc1ZmLTR3seuZpoZge6XKO1rqEaQh6ZNmfYRS0wzkiCEicBpzI0WVKXwVYMV6oYRmct/PG0
vNFueFbhrBqlBb4bvYrtgNOKpOz6yVjIdbdrwEciENvf+xF2J1++oR15MFMVLjm9KbIBIXupTNL5
z7W/VWej9nmoagq2ZAxW6eT1hqg5eTCEjejeRyn6B82FhPf1beyzcKsoc4ULdc94SuupVcDkDFEq
+p0+dX2mAFjwxQNXc6IKApEtbUa06V9s329Uoeo5XGh52x6gFmJuBAS8mi6zgxNHPWYIq4eqTu3m
jMlAsrthhHRWoni95SdkOUrSJWX6TBoOBzmYR19aJ7iBSqnuLbeR549tFJFNvS6zf4yFICEkpfi/
vAS5pUVGf387m59bia2JhZPWWEHSTvcXRf7tiZRVHFL3NylAhahpYHXeSpM5fWAgZwRN1eJKZvtY
zhoeox89HE2mmzIwBPHuDSjJyPWzMBojprady7PB6DAQnWfSDvl363Ht8SWphbb1yBsF5RTBOlzB
KjrmQTQ+FEKcgx+vFtw30b3oTAFIIg4gvIA4uWN/mzq1UU8amomoM2GQmcmSuQRP+NXfNHveKAt+
r4CTNTAPBZaPxP+GSknKCH2PKluuhgt4EDwEkQK0wolc5MMIMjpVabD5TcHR3rQgC8XXggE2lXLb
1U0w+KJ7YGfe5xD2l7i7JliYqn6UkNdZ+cAKPVgAAJ9ne9nWjhoaR/rwpGZuYY7IFXubNClM/XuX
Jn9m8Xop/Q8K4Aaxtw+z1MEwBi2kKwNaGbUnoIYyPoNhLHaKETydTzVOtAQ/1ZAcPL85MkVb/h1n
5h+yYmsll8sHJJuyvm3WnG/+5TRZtZgpjKj2n2jbUru3QY97V15n6L9vRci2xhOFdocqorRBkz4+
TdpqnHRRN3nRtn3VDcpJZi04QJe5VVju+wKsm14GINKunVauw1V9puAMO6Yw58OFtMyRK5ArMIZx
uAEpVt/uTvfhAFXCPKzSNwRwNbYQll4IcSXHpnUmlabqTjAmShgQelwE7jw0YJZYEqHMT1xrewXv
5ajtnJNuLwIUSv2zxQfSGYdUW/JDIYOMwnIwxshjmliXo5wOLWKXX22/utBb2vK+RaEdLTZWo1fi
gfosg58y+ZDsLZHbw812sv0oRfnUuSyOz3sLfcg7MeX91mLiQXy9hqO704BYfKQY8AjlxPBxHU+O
/wp09QogUXnxW5s8xj+9fBJo2pvIj3bQos+WuEeQn4BNtjmIlCwfRtpQDrgRvVstr5LN4tUN5vDW
9VLsTFAdOZOlrApIJk5NHuGSOTgrl6L/AH77Nt2pvnin7bm5h7MeYlqf+knFZFpn1ESrKVUeR+UJ
F/iMuCj0s0B39NcfEfR3ywp3d4FB1SDcfxJUhhuCnn52hBTPcxPJGZrzCnudgUVheNq0lUkOOl0O
dFO6Rgw2wlWMRj8QbiTQEOHTq2kbqWa+tMnt3DXmcST/TOsBc1X5/+X1QptDy5hmiUx0rlMGUhCR
StsJoCnr2ZO3MFCoQz88bZQN7lDFNemZvvSQKLxEPeK8jOOYTGmDv5E6Up0mHZl7u2BsYQRmC0i0
VL7zZYForv2ZypjvjMLcqT9vmtfa+1C/WLkuzuL+sy5qsrDEukFT7M5I4e3/VtFDSBFStB3Fgpmh
zKj+EzSTwcZMuNcqzJiEwWxxVvrzRp1oVOU0uO4gz2gYiqpwAiWbHQCHblKBg0grfIIKb+7StBHx
7byT6HG7OQYnDARsyrLImfjBxiiKxw0gJD05ZyUBtN288kj63L4kDDqpJ3Yj9FKeq519rDlW6oos
Brg9xYalVrPZr/iQbNJdaVhoEi+8M9GqQNE7wqO9nYOeKC4XD7Sb7BX3iO3Ida5OfGo0+Oeqk2Sq
NORHtiMLi7j52Z9wsB3rsm52GQCksZz87KfbUwXk8ovIw1LGb1UpsywBZy9caxKFINL0bvfqb39i
A4coJmQh94HUvEHkrtQLbQr0b9Qrseh+cw3mliDvXlaqseSbIErYKKkzQhaH/ETnao+wvfCa+QyP
yJ0ei8SH6kczmEYU2yflb+NiPSUk/ykKv7/HyoX9apXrfW+40TKVcahgv0OWN8n0M7jKsaSOGus1
m/DyjSGefyPlOiMe2NT79UOGHa2FFKYqzWh4p6zZtVbHNFcwaHZsSU0r7wkzme8147yp5lWmisce
iNJs8wSp1IeLzlMyE1NULdzCp0Xcizx3EUMISWQCGIQtMmFmN3FCNUU0hFTLoPGTH8vtxAiyuNvT
Z1Ga1iswtkCfibOWosxxyZj6beceZAdsIL5TDFEekHxTeE8BY2NBKuc/plpo30agCto1nh9tNZP/
JETgvbbVj9J0fMbcvQQfDRZ+yqzdTln8Nex9S9AdfSXLGC0f9hSaAmpt6rn+B1Ee4WD0O2AxA39k
oRC9TENlhCi+gnM6D0QuHUaUgi0ggg7P9eLHBeT0jzVP5pT+0PgmXSKp1RsAffvAh24RF+1lQN9B
wZ5X59m0/fEZZl1jalv0J3WpbXXnpWKSvUvUlhpgu9jiDDM0BfLgP83szKrVP/QqxTDU5+74GyYR
mattt5Cwq/Q69rNd7vMjZMSNLbVS8bYrXOcP8JswJ5+8afvWXZqZKSvMFVoubXNDs2N56hvDxnAn
U9Xoznk1dWVOT0I+1/DoK1d2Z8ygW7hRELBwuJI9slM2QnbUZ7IaG3A8VMVWrYfa8YdYkbDPsMf/
rElc+aevYtYaPURKSAeVoPWSE2p6tUl0ql74nG46db8Joqfx1N2nZTAFEJ6m3ocVNyqfz8yoeT8A
nC2s+jUmj1lYkjzfpVjL+bkf152uCahOQDt/+R3yhZRtiGLaz27VlnqPlSpf2KQ1aRKAu0H1x1hC
s8b1TNbk7QvsIptScpF/ehvNCFKFhIojn8HllcNjAHirYzktH5ID1PAx2/O0N/FZPzJgPNbBtxW8
AMxGmRltteYw9pn8tsPevIFD9YGIN6knlM3TLEhTbs61AzYTkWR5ra6OcpBrB5Jyfhgu+h6W7aDD
8ivp7vWcOG+nmAs84vWne2p+ZwOA2+7t3Mp1tBRlM4U/yUelRyEKWQW1qcSKKUheb8p7h41TuUME
AnJ3UqVczlaZh+S2BSXj5KvJjqdVLcocYXIriM6POKE1M0/UBiLMJ04GyMSZhpRXXu0vguLmrfAv
w1Wdn3lVOCcy7y+l1FNeGOTaWCZkeSYgf2tAp/5pDiLo5CrPBs+M4nytbOJ2mLKEnRs/bQ/8JXSy
W0OClT/zk5GItToKMi2ZsydmdrrZxnljQGII/7dfEuKV/JIpj6EQwLyB+TviOpQow+HdCc05QpUE
cAO1rKQdNl2T0N4QsTFnMfpegMkaIoHJfr7K7kESzYWWMqc9rNrUv+CtZ1l2SbwX9cTgARIp6OFy
sLNi/KZZ3+pjCBCKDOliD5FNqqRXBQMiL9s/PvNrrpUawUPEJ901GQHs/bz1LdP9y2U5/QLfIcOc
PtSjGpR6gr1jDARcCgmrxlGt1HAr3T4AW/ID61wldvwI7CbFBIcMBr1mJB1JD5kZkGjiFl5Q46ao
kiR0blyoPvTYT4dEGXwqHPziyfUIYpHi8jIGby0xLg2vb92I1iAtefJSZA6ckvEQfMLWZhvkPwj9
Abhq1MJ2Utos4cgnOxT5OcoS84JtTbsgLEgH7MP4HZtO7dW4LtGP1KGAWwtgvgRpfO1V9OnwDyOH
kwVn1XGdINAgs8maO+IxZumJfMqg3IFFX+kDT2plR6mnInXZBLXONoHlJJ4QACRNnuZRb6HK/5rO
QCu8SgAZpCISrE+/L43/91hxcW8Wi8UjNXIK9b7WMqdL4jh2vedxjhQjFtCsO5ZswKBzaCnkF0Vy
nh/bhfEvkiIxJn4Ib/SayUMbIa8JU3PkSwD83iGWquKEocUtnq4EWoquQfJeVhi6PhNe6ZzB0+Cp
lOBhr1YMTTgxKeW74i2wFca0PgYrHLqBBP9NspJFwhcw+IAI39xKCKV5UniNetuC9Q/i3LWs4ADH
zTMCco1ndHJoO/85k2INfZR4Ti18DMSSVcyOpLCmPEFlcbw2/B5HVri54o97zVQLU+gJuJiEAylr
nmQgell62rAq1miczYJK7Va/qMdmdeRYQRWpFQzhbvi2Cg/d4N3H6L8df38hn8xK86kWDejENq/C
go8CWOpWmqh6vNmy2XVqHZJ2BH2/k9Hji0NsCFgz1pymFPhX4aUdL0eUN0euJCwoHWit66rxg4Lw
IGA2dSXx03sIMiTkrsUw0drU56rrF8wx+tq/qHmhufByyxQWL+No/Zbq9n5OxC2My9YOpnvO5cB6
s1ovLKKzyrCbtftwCziF05gASbswF62eH2fB67K1N4t9S1TzCZT+2Sz+BK+Ffzrc/WGgdA6seQWF
unPinXbcj1a6wHKVPWFURpMMEgCNNY4z+3hJvsRhOehmorRz1tEBKqrDNHVuSGzW1lroH4Bg3TKp
ig0F7fo6hQyC/Pf+4DXjcofA4YoeE05IDtT4ZjcrAB7tdYHFIHpZBu0OjF6epp40pFBGs7NRM7mx
HHGulf7IDHAjqcOfQdIOiUsCbsHdIXnhk74mPYYpBoXWLqhRZkWsSX238rJoQRKw4OFYGCFOYC3V
vWKcEqiKqoZedfFCNTr6XEHc4RlH6gvHyigWqVvby1arxUycSwc/ROfNUg9QJudfVIuI1+9/Hc3r
i+u48Qlk9Ah7F8fygSUbNhX7DAWjBlVm2cQoMLmRmqbmI7IWoOucI8dAWE98j88XU9ZtNIZkggK4
0jgSra+G+NMKJmUzyxRrfgyqF6xTq31HsaEC5isJWZX8pwo2aBb2RrGpn0xFYdsACJITq8/4E/QB
Ja601N79UmIu0ZlXDqf3K+oTD+Tr+xpMxLrg7TYtB+PpTlWossmizV61DwtpcxDqlgYrGJXQymw4
gisBVsk7+Gzx+MTP2vVWvYHl7oaYSr1C24lkYJ0GLSAWaPouXU/Pt+wFjS/UQD0Q4uzhMl38TxMG
vTsJq508GqM2gPfXyrOiOBAMjjStC0yvnf64WKF+YixABWdwMIRd1Lh9whL1Fcbnp+l0Ut1w3wF1
hiGOBzTPYSh/l+aDP99Q9KA2iLvHKCDXzMX6gXvCTynoJfoBH4exUiwtQ9F+YCE3yJmbn0ZIx1UA
BwZ/pOEI3GsunpjvdcgDkDNPfB3tSroLzi1wfmpDKnTUn1s+mMggzoi0fV+Sf0TMIaxmTEu9oW5H
iRVcASSTdMTdCRDTBYv0aErkSNz998hBGPYm10Rm/I9X6qdhwlgg1iQElqJrpyL8pkzLcHO3xzyT
BpidW+JTmykkSxXbQvmBebsT/0PWgz21HyZSa8qD3Djq5KA3eHs6B6Zm5arqJxDoII+O2F7o/9NN
AljapCtadHCHC8xoxaiKmj957meHzQBSTYTPhHM0D6tVrjxn1cPCj1gIID/PUzsmMVSckvL9tTNR
pUhFC76Y1M8jT26pCjt84IV7c1z9oP9ABgE3QWCVGcvnozQV5nmRqpGFXZlYDiBGYQg1WrCcO4Ys
HbGFEEAghHqSY8tTWnlVyaihkVPbeU+mMgoCJaBJvFvzsGL+tM0NeFJmOGctq84ANxWybyyIH8Uf
rt1aXMNcUvZOvKBwEw8ZoxkAi73zBLIcnBJ3Ir6x7lyS0Vyf3M+R6trUt6KfEVI8gGdL+DkL3GfK
hB1mLk48pQgCi5Qf9w8UYo5gAhWNlGyRle3vo211f1vCTDDoIvdHALzMDFcAD/kaaGR+DL0+cRBy
H/SA8sirS7RrWvkUpo4kbEZCWawl6sbWeVqQVYKYIGT1M0/ua0+86FGNnsKk7qeEQmYbNOmjFhGX
Nn6GJfa9kS9eXUNWLoIPbv79Txl1u5/1RYlBzDhmiLB1P2bPtUq/IEkduSAQRjv/yUjUA9y1nMpf
+dTmpb5p/n7oCd2NSTYxKPWsN5L3+0jF+QZDUZudRpvt9OC3UFOctrID3uajlNfGQkL9/Tu3BgVS
8bEYyxzfT5Zgr4JjjwsNLTjH76OIfgTuhZ4+MMWzy745vHI66aCFSZoVDqAQ1f/ONLlAcjQCWAmP
51GVV6SVrkWinMsPn66FBaOE8SXP6xIiVpAyyflkWsaZk5Dvuiao5lpUKWCFrctTVB19SZXA17kW
JW7lI1Jf9zDn6YB3WzbDj06+ytpftM9M0sFrkyei1ObazIfbQbd8lCkopXjUezFbSdKDvZtpR4gl
HKkVBPNmWW87KRkPrWeN0y35Jzjd5T7ypWunkpy6tLcyfOE4hcfo2ohKpyasPw0eXVQFPXxecZAs
F1CMZXA+rQH+LZw3CXtn+bTFWG13q5IZBwcKLO3ryZDFwEogF3Amme76skIzM+Vh+qqJQyyHH5hX
EdiG5+mFXO1cqx5cp20RN5wdRZjk3rqPu36P1ieqVmoN1OGmfzFzv86VRVlqXclQRuhJ8cZ3Gl9d
6XukmASzB/VQequZTjjVbSEhU7301m1folKf3LsB/jTSvAb/gMQiXGdiiYpP6AoXJGwP9yCYSCFI
26VogjU9hsPZlsA7Lkh6lW/iYUg6fSO1lrHXOSM5w7K3H9vXKSGM0cE8Nd09ntFazi/o0PKbPr/+
7X1HqdMUA2VnzU1ZiQn0hLSnnr2Uya4wBlZpE11fjgmA0bvOhK3Qr8FD5hJIbEyB5THJ+YbGxKI9
C9LT957l87l2F2RmXQRAfa2U7lqfasRQwyQNUAmT8fC8ZWpiiKIve3ZoAWi1TKUzCFQAIDY1y7Z2
sgLWbLmQVR4iIPxZAbEy/5oYVGOHU8GcwsawEsHGk/wMD79dVRNKeSBA0KQsamQ6sZ7gLZoFYsmc
u1dNs8eEmwg3/n91Dh2cI6i/HqYT/KknzUen9nvPocpE7jv7S3Cr7u1W+PrZcy+M3eDIqhxXZCte
2l0MRoKNM006/DkQ6y5oblgvctKTEWyhYlr+dw+6oaUom1CtdQvmCzWjqVL8+yJFwtC3JB3NFkqR
LYKM8CAubSyPnZhYgCeJo+/izMHMB5064ewkglQKDfSki46QEhLnt8NM/vS7/Ouh/TL3Lms0/jRi
Baanw91BbSI8RBJTUvG28MHteWoyZh3k75kRwp/YnKuuEkV00u89/X2d4cQLJunaTqKT8oL8cMQL
qm+TNt3KwMSuP08aB+nLvZy70pGxnpNaOjhgn4rnQySXkK1k5mDQnOBQJAPAg5LOBmXoZzKiYNQm
dmQw8rn8lI6InnmdUMB83EsFTmQbCpm8P+dhmVm4+ygxou3k6slGZeZQpfBFCnO23KXO3VF5J2kn
seus9wf20zXLz4YNl7kiyT/SfBwhEZv1ozCfc09xjg1UZp0uzXHicj11dMeGfJHNoAurEb6kJcpu
FSO65J5nCBMgXGes+CsbRWN0ZQ7UhrVxCTpIMrkWTRChii0Xm7srdOQXMxjh3M8qKBtO0fKcUyfe
gPZ/ZxA5ETiy6dl+vSGJZKJPJqD+rmrtYFTCWioaW86hjsPp87hpMlyJUtykvsXlgoXyfnNgKjpL
BKsPqyhNZ6Sx7FzzRyA4753uKQYt5qLYUDo3GVUcMEJ5Um5CUSu/jowL4o7JBqHQ7/c2B1t+AZQN
cl/IEBnd0bnYzcMVeoQ4Iucbos9L64K80K8LJnIZAYSbspmh6teHoI5kC0fltvdMnRvDj9bc8HAr
JF0rqby6+cwyb++S39p159hfQMk8qgUeFzJZ5MNeS56H6TdAtD91LzF1MsW6Xfqo1ErjSYno/B3c
UtIoxTup7NHlaNlJUjVfUc+ovoLGXmty9R9n2TSYBlEXENuQ0k52iaJQzQ8eBcBraE50595f2CFA
RcaGtP37BtETVwgexV+E/J+pXv5ExDOc3OdA6AZjUemdg0hEeN3aK0zjjFHm91lMrEIBTLvSapte
slrxHKhZA6nWxtGhQ4ArHkWXh//m6Y73tmxCS9f7Ge7aHHc3jUDjMpxOc1IQO1cUk/9vTePfdz7d
p6JiS+fT8/hg/CS6kUwWWbMIXTQRYXl8Waz6rxDRz/x8aMkxf7kyUW7J2cAcRSf0I+Ztclqq1aXX
rRthcfm32NTwlINdDszJKUkphZPH+1/LpkpDCx2aWySgfbaR/fJKwV4lACnfsJl/S7OlLAAQ7S6G
u5Vq4tdDc+PoCZKQ7yiPBJXddtJ4zE3LGV5Pp/zptovywgTXBVm6E3ziwKwaXMh1rS2UbH6/d612
19Zs74lyzzfaphXYhdga84/Orq9skdjKHl036w2eVXLR+vMibmqaP2UcpnW6DlVz/6q0yqdkpsRJ
FQadZW86th7let+R2y85Bq/JxJO25/1j6ZVdEGH6BvQ9s6Dfx+bwKey5heEjeeBiUyZ/qPi+cVd1
/khJ4pGjyQ1dnjElmuQZkj2k6RF/LIOiESuXCUQZ4541fTlO2FsxMYYElkXzbeRl1hM8vgeJ4ugo
cKvLEIto6WEfRyD12SRiv5W/Zw4Ji4hmR8JJ8VZo7bBQ+KclluiNG8Qz/kWmXayvsPdwBBjwHZNE
g3BicpqLrELHRXMuXX3jlJBRR1ThXDiC8OZd0EZnTLHzfCJ3JxbaAWmV88rXY5lNuQQusYImXPXI
6dcND6qpibs63nnGE17cNIi4mjx7rhf+6O2dO6IsrVcjjCTFTpgC24C9evKmnlKorSEPp6WWNNDV
wHgLoLK3ctQk0cxXO1Yg/H76jkl5LsPk0xF82LsWR4NNb76x0lVCuZg4GqJ8hF+WTbwO7cS4y/c/
fceR2/P4KQM+6DNRBZ6tt1b3+u6nuEtntmVJhiF8Ciln6ArroI/4IIXua0PzCuZp4FpLXWIXcLzF
1K1YD9WjCen+p22uNg6tuEJvB1s7BMEMI7c4jq2dgw2KRwsRZfl94t0Z7+Xy/tCPw6WP5MdJE34Q
+Ig52z/E/XSI80xwoaJLHxhUYF3zajiJci4dfiVwylwFV3gMIExtamgqq/zwkAwPpltiswJKGOIW
T1mQ9wHBjSW+PJ8zihYf8569mhHXaEioVuwGAQGf3pQZ/rLKutaSDU2q/rlfGTnImpovVVzOZMec
5RbHmZMPBFJxYinffsGxYRpOo5hD+k1Y79laFxGPSkHqRLWm07xeaZ6dQ2sMfc1nEXzkDVB10x5z
UYFdt1DjIWXQIPo/I0VlPYqTNTc47RwVPPKhYhsrquvpO+GnFvJLp3mwiBUoNo8Fw931BkJXmJU9
N9/4fWkUdThGCaoqcVEeMn339ZBsbBM0Rmt/CQtZq6Ru1O37xf3R1Eq4AEkGofJ04Rfi0fnh9WTW
tDGUlSSFEPbGhCUad9Vi3/XWGelSE96o3oMVD6Xmrze+lyah+HYT/OuK4IONnHg5h08H6mJ73lNE
vfvqbIpsX9DflRM02nEWkYOwSMWf+VRDevYNiblSzqy/eX676RO9ClB1c4OzTNUispkZyOjJUo8j
qwkrhL/H0xcFMeqBhdDP0wEhNi/XCTXRmy5GprNGMoxxY1CrubqEc8YS3LvHEuJS5asWYjJpBAfx
oznRZliEqMrojIR7r9qhVqrfWJZwoMNx30iI3QLeNOupKXtP83Yl+k86ZBhzHlDUXHJx9qiMJ5tz
ay1C0r4HFnn8F1dDPc617N/aYlL/82YHq/a7A/WYQsuIeDrRI8NHI6qeGpj+lPCMs1y6iJAa+uyQ
SSKxo5UrLjwNRKYR4jVXsjWhbccGmc8wB5IuiwA0dR1ZxmNQw5Bu5KqZ6lDpBgSBnjlaVSEzAzHY
q2ozBB7RKdoAZnvYA+5Gtu2lVSsfIyHTTpdb8hI+DzkNWkKzWFQ7njZA8KXKVYXdo480qbA+Tua/
dAMhbA1Alb1MfxZUoZc4bHwUVR977eGcNgHeCl9fURbv0l2yxVyPeMVXDCAE9VgqeUE6a41n4jhB
v7MT6mDzlBJhBTMirI5tsDK2pujDDd+WmYyDJ3SVJz+DIYTdlb+xQNf8U3ILisTiXL9Ph/hohJme
MDW4fAEJt+jQ3dAPs7qdv5CaTOrCp1X46GFdKbertnjFjW3Zi406Mjw39FbKAZFhOwbGT/a6PmsU
g5+uK5Qo2Z4aCjFo4/GzMGunsF01OijY7HlTzBt9teqeveRTc4/cuz+qVyR86D2jtZFlV5uVH0o5
htYwqPm/m47+cwDkzJi6dMn8ivhR0iaLzr8JiFjWZKxGqrspOuasbbSOj5Ooq+ydTvdI0SVf4IfY
y97EHcqZjZBac0/QqqT4mF20Y7UH/l8etl3Y5f+3VD03SB2Sb+XJAZT2IveVsSBPrMyj0JVbyJUV
xtirNlJkQjAbGpVyqdO6lBEHtE2Eoz9qpVLU0mq7e2wEhgLRbhrY85TYOTsXkR8ue1EWdYoCI7Ei
Gxfx4pGXqq9tYjyn120A1IO6jW1YgRIIBy+q7lXoOPbojQG7uykVh2rZlNPaJLhwwMJE5RHuqZ8Z
33ZhdyJLB+lzL1tm/eMu7RRmdAjkcuxZWb8uZPR/cvqgkYwJqZ72l80bpKOuNsAZHwTBg0hSe+dL
GGLzZHnFzwCGjHbvusdjJXSZrwQht38yQjZAEpp3xjRmhQRGzkxHxX3uX2Ab53jYPPPsEG5hRqzD
2Zp8pVI3DN85a8/xkM28CXuSG3sKFHM2CDRkkFHpdwRddbwN+W8XmhEs56vKvsxjqMzRVM9XdlHN
8SjSdLrOrnNqgZs9Pz0NTs8UzOlyzsQgPaBh4N/t0alNAMQElES8DbzF8z3cYr3p+gs5dS2SBJhC
Hw+U/tTDxY9eUn3d4yYOYqyJZL4MD6zOtjH392uObLnoHojlZT8MFY2HDjDiGxITIGXKnRwh184p
AnVPHWooHoNByKeZCjEr7j+NyXwEhiI128xeejS9KkIAJdGnyu+xpHC3uk5lXpRiUupFo96b8Mml
2LqZ91o84H1WBkiRxxMmxPFOoZiLYF4AWL+WDFDZog/yg2zkFYIvstxutsy0/B6OrhJ2U9O3b6Yz
wA6oXZvdsMzqinbo8fRNdIvBcageV455EMaLnM7SgpUbz1AIP8+oCsKGq/ciWVFl6wsoIcgHbV4s
wP39mQkzg92nEESt99nzRqFPICws/iVvKelVtCrs6+R4RQYv8yVJR+I2JOj3H8u5O86uVJ5fjrWj
DTjuGWTDuAqXX3uJXbpb9ZVWmebRnEnBQQj06Qn1sP53Wzcku83DH3fOvECCt1R6jRvhKgWTv6fU
e54zFw76e9aBmwAtDgSMJ0lvmX9nqiVhD4Tgy00aK9/2C9tYwUFcJGtPbUijHq+3oxq6dnhj7kiA
i/DLPPHcx3ScWlSiASo104mYVKKQNZY9ezUTLtOYC8Cb1GOIUtXmjlaOYxNZbTa6am6xUESkz+jM
B1uLeXJciZnpNHCVvg6WYWVtpRVgEIiz1Aq3bp0AHS/CLGwYBa3XvjL8rCDZMoZxfdLwlojeZSwf
sohsG4ClvxLVfYZ7gWgOmoAsjF/pzCcRBBd2Jon8E354vmIMtp+ONcBGinE3G7VqgpMT0L4vQroI
CAhD8yx8ig9AvPpFXsIOziBztMHdqHoMIQghGl35ZvFXdDfmymX/AYP56jnIkExEg9F2OTCwBUNM
VczW0VxSVCjgDAlyy3C08v0vfKyHIwGhh97NA6GowrkFQPN5M5b7xfG5IL/EhdJoQ161cB4ggZOj
8QKgCHG5wL0gGzlU6HyGCnkSk0YL4YbbKwkpOGyVSc2toGA3HNrvK9Os06zVLeSzxWJC/cSy38T8
Td0aNxgRsbre4iOw8CLnszdCwQs+vi8qiGs79DdfCJlO0teEqzg6/lLJeb96WKmAOcggJdqHGUGS
YrT+MghKjnl+gMbyD9gwURrafShjvYUy0cT69bIwZcbwz0iEdGeGaGcKW2p9AZsMmT5POSj6pt0a
nfulW3nXUSxDrlabs0qS4aqIpMLhc5bJsWpmLnotWgmspJZut0T25DU2k0Zlq7o721bvMHwr38Ei
4evU9j4CfwpqYCOfI1lKT6MGooWsnQLDvf89hL4Hr5yTYSxJMVUi7qWoxFr3UtoKO/ZAsjud8wsw
SG2nppF/cJsEz9yc+2JSnJDutb3aTP23mbzfC/5G3cA2Xd6ZkS8QJSiWNXwEQsXRtuPDQZwIFy11
02g1wADMwYx/x5AvWqVTFpyMNuTC1Dr05Rg8hP63PlgROgafdpZ1gqeV1YGwA262AUg2IKZIDNtJ
c777/mvidHneQmaWbJB4PFiPmGfb9qqEM9s4ZY4HxXikDrJvsT192jyg2WlUysbVKbq3Z9LNrz/r
NBA4OIGzCWqP/XLaGHq1yMe1dFqbI5fYzYnYiUv5DORtmFtRTLFhMw5eiu+HInOrioPpsJ2grECe
ssTvnsGbthNYZkrr28e8mnTo0mm1iAjvylP9bfWqTUk60iUdP/9Na+Z3xvNdUwpNQDNJJ17BAgus
dliRN5JBxz/rvFT8PfrYhiJvQx9vD+PNrZfYK+qV4EFQxHVqh2E+m2+kSK2AD7AT8RTI678+lb+H
ymB6RJ1m3WR7H5g4k/ERkewZR6VhCk5iXr4VDouiCcHhcP7R9ltczmGcQp8NvGd/ZpvbMcYi+UOK
DN55DbpVhFfHKeM9YpNSgMmG4O81vvr9NSMjsWJs+UgN4do7AVBpTzaoJcrsTACbH9+FCHess/FZ
0mRrmsCpxD5WZsPMHjOfQK80M7mkBpXEmwGbX9ZydXHIhCdJ4sEJqHr0nBnEZpsRIKfZBqJ4iUlM
ZP78dUdGGc5LtPk5nY5ecBaPSDEqTJtvS/dBte9reyqcUJER3D5DBhS8+a2+MJSJTudS87nq5mwy
GgXyKVUMq8bK28tqeRtHMMGuXQLBOfUyRco8/k/ur2EWXvlXin5sbs7STBhgiWbdVvF6EkHMA8CR
bEzgJZIqMdn4iE1kfbQYYBWmcyQOS+arMXNZoB8KC0/tpvEl0BvqUC9k2LBMBEZLREp8lTQ2Ca1F
BMJ8KZmJsvX0YyASI+xcqy54llVzadOxxK3cZGEsIDNmKRlEXTwxb2ELdmK3heMXuiFJfpSOGfZK
Y3rcP4Dpal2L6EXLxggUioZgsurv9E/5epFUheZlzElY7rFpbdI+ZPTMh92Vh+Lb9bHbYF7L9GR1
WjljGrpmYabLVTrimwqjxfhXFRwczug41eZqLGRqlrVpRWCghOcpCI7knVFPP8y5C+W1zdilZ4SC
aCasASxrNDUqO/cX6vtxV6bvXJ5ULQrc4HB2tPzxkKqwpdmRk92j8b+iu3o0C9MFlij3fQyDmmO3
8QWkDE9ftCFQkbAHLpm0j7SDF9bMowmfW0nJrDfMYKHw+VyXXg6QEWHxEYHaONkwad+TnJ+4aFIn
QpHK4gQEaLMpsWOMEBfzdyH3PhgATE20xubNocQuSrQvC6DK34BgYiApgCYcwzQjonwXGgbMi3Qe
y6cyF0/KKPm1GthDSzRytbwsFpKiokCKB/87PKoHPZXtsm8abeaJbiU6Wf5Nkgkw4fdzCynXW9sR
clX1zsNcP3aXOF78t1yys8vJfRolT3PNzt0yv2gcZ6WbiG3/18I3J0Qdyuf5egMEtc1JQZOq8VmI
QLr1GwrcgfQmjwx309ScIdK4YJEGGvbhCRtNs1hrTb4X+5gcrAEAJHit/x7YYITlE1zTfcgocObk
rGcn/7645NICHOjoXc4gWneo6YXmz7JxYPac6JJl0RjJDjQez3cgcMOzfVB1D6uFtQTuToNDFj6I
3fIujp3MqCi00EDskzM5SBYI0TgmK40zGGCWFFDh1/psvePjF2TjcqftEAALFbSDhNACXoymbYAX
be1sKrWien42UlhJ2rz1bUn5OF2g8yR4KpV1K5rCfNw9cHr8Y2kpOplmi0l55qw9oFzrmVh5+liu
rDoFJFuhPmDs/Zmm1GMuqTCdun7robcM9plA6oxJhgEVnFcoBlkNvy7NHhO/X4a9W+yvKrNxMHmW
JfhYc5nWprXgpTo7GiIQg17YQWK+eW1Sqf2SABAkoN82E6YUt0LZWSGkEJMQke8YO5fbcN63JLUL
O92c/l1vgJWiAQbNeYkVKJDxJfZYoAxJ0gGHNZH+4vuSjMBVnrOMjIwMX/w6f0blCEzuWBQtfyut
T5mi29jUqy/tg2KUPrVW1r6Y5dcOKZr1gAS6k11aAsnLEK1l4JO3sFEvz1uOCCmmkAxkf5+LUN0n
D4QWV9tEYB8cP7Ls4xx+fylnqjHxXZBtYo5ubmsi4fyWXJ/ERMynyfbZ4sWkH7ZNPCwZ+IUXgqzd
3v1GjeLIvScNbrMch5HSTkRCF6v02V1kfa7kiIDe3F9wSTaytJjD4a6n0Me0+5fNO5tSIzn/YOaz
bpDJhuS2h1zk8G2bOhv58Rg8agEcvbc9YzVs4chWzwPV9KOooymVIkh6ElTKh8TWPwEtSlQwrbr2
gRxCEAiyha5H8kA20Fkrl2gMJ0ABUFGGzYCO5xxLJbjWA3N8pDqMo5YBBcLMVK4bJdwwBxCJCOu4
QmXEVmWg1NsXMYJ4b4VOAyLcF9rsUissHzgtbABg+a4Y30SbkAXY8kiJdzAkqAAuTd7xYPZlKZmC
GGpvgsj4fqKrqKhEBL6qzMsFy1teUhfYUzB8dUZgFNoBV5sFeQPANL3gsswI10W+CU4sXFRF7FEv
8YfEd23ioDUT5rJCXOuxUxR47jJEONi95yaaSH04vA86S8xpyQzpK7l7N2R8E9Xtkne9bSky/T06
3PM5rbGWZj3MS1uMYeqbo1SmrtsRpnl0CNg5w6LC1fGVsPH0K5doPn3L7O6XPONUbcAvBIz7qT8k
apoyvw0vUq7lyRBhzs5uCpvFzB8+UtGbWOS72KqhjWy9yy6o4gMpULajpQ+dTTT19syk7ZgVDFD5
w/ofxvq3MHvEkpqnwCbXkM6AKVOYwq3AtmPuFyg1997Lr8eZ9b93Ci/t5xmQdIDYHJzwCXWGmVjo
D4EhKNH2Ml35NJzJ53s04+/gqfnsHDru0YD+GvNqmpiaNXeiLavODVil2jYFHfWj0ud7F7vVzc4I
r+oaBcNtGw7aGKV+t6opiDjBNW8tFcmhI8+HW/XB1pvxLc6uw54KLHvm7hwWHD1wqHE99fGPI+4k
O+P7qXPSMraQaYpt2e0peOk0eXI8JV9zZbBTUApx1RYidtnzcGyKWRRRt0jDplepkpnMEOq22JWD
tiCEiOW/3gKT4Br3facbarI4vMw2TfBnskmTocLZf1w66rZ86LbtQGLiZcFKU0ZI50zlAhQ4x/oc
kgxSzb+1NDEzbIXsDSSmXtsd5uKeCuR7h7SqtKQKA2LUyIm2o1/cPy7XzPeLr2EQq2QWLIZ8GUdo
tz1sLQCNt28IUx6OFx0i4TGZruOkBUDP1UwJUEk9y0UjIDttXwlr0RQfC1+vPkJUsifxYTXL1Zgu
yhGpaT4gShBo39xW0iynyiRRjtFN6zsbMbGMWMCBN+FnwjePPXMale0muFVeas6ChokwKaiR0Il2
VeOs5DWUYD2BB6e34YdtQmDnDT0j/C6uCuDyHmgMCgBndgSIiw3uWEvWwqfsnFWIwkW3sd60qYxN
2LtimPWz5S9Jyc4cOfspxxZxAHGUxBiqUZtH3qwiiXNuLA/Ud9HhlJC+Um3DSq1VbB3Rn2svLbWm
vvR+20HhDoqugw3EMDgojX5DR7qcIRzjjLztheQGkDo7qXwNTQDHmUmGCOm8Z/ApxxCRq0YfLcu5
v9bALtXKF5QK2dI7GBkWz9zTkdWBCgyHQujHkCIYgnt6MpcCVR0kJRo/ukttilGtStHwjOmB36ne
5UyxWT2KYPBYn6mr8gbA/uyHAbNwTcVAKyjMy1AyFQxZa60axnjaUEHvLpqzsmvWSUE/uog2p3Ys
hrccqwF3g0WwRg9cc8PqmEoccaOXXjl8qWD4ZMXMeDXZeMQ4EiF7ZsfBfTEmcaPw5BbuAfuUJcxp
wciQYO6h0ELgn8XZ4q5gnaxiDxMM/0H8RV/X+ofaQRyEtNHK1WQDjE0gGFN4fSq7V7vuNEWS8d0Z
1wR40LVBWHV4RCpQ+T6vSx4cdXj7j/gdV6UQcgR1i5FAHYjL2TGKLrL2IoSyY+jPTkMp9ortPkBx
9FKSY2g1WPj9DCG/N8fPZ+u+TjhzXSjmrvLAtxj6vF8JM3E7QiSiYEZwOE/UuTNUxaDsglj2GeG/
cjyNliDfmoMkuQ/XQa27sc63ykisf3uiHwbIBy/821ri46PgD6tkcRc1nMTmPPCcIXTyUG0Vzfp7
rN9mxPfaPmH9/C3cNVPhA9UHARFqH/JMLJcuswSELyBgUhVD+PteEjzndctmLR10ODVkkpR9Hn93
3xSP/Y8qqWzi9/y2Z1OgOrty8lNczq4I2MsjXTC3nZYCIMuIxcniYaUPUq2vU53oHSQ85sB8Y904
MmqHnM5FviW4y0CVLCZWLt/U5FXBOLP+nqVk89v7XSj7m2aiRP+3Dyo6AvdiKo6ThjuRxn6pOUJt
8iNUmY1Iq0SzLwTI2ouHPTmTFn4Njp+m1GjGuTovd+/26C3YYlImHESMh/Sx2a09jC6rmpn+3E5D
q3KgWEC49/brJ8oTCAFGxL9c19CxmHS0nkVl1WlaMavFtnYvw52rIuAvF56wc/FjvZ8C1djLwfTg
p6i/sRuCqMTMBfnXgl9cyOQqWmSKRcVvVlp8+sERQnqcn+c8pXqizsOL9QeZqyMz4LeLHtfhcLzS
OKVGX2TQnE6fdozZAX1y0fNfGqAygI+JPyb8I3jLFJnDfwnNKe/Kaw9pfq1goc283dcTHNIA33nw
l1T/JY6TLdIwD/rIBONqPVhUKEcshFvJ+ZFD7syoLsLQZNtCFt+mNffXEiOav26Hc3uwxlao4S/o
J3N0XL42EgHl7lSdw7UeQ0mLA1rDrGJh9Sv+kiu+f6cwCs8xOOKzC7Mp0if3Ysp2uFscpyBLjOEp
3aeO4Kt52wo6Fi893efK3ayR1Amcps5SzFCaVsS7jac0rYS3+xjr0ChkJ+d5uIWAgSCqD/mkObmV
6Z4b9LnDylX1aYVBqr04Hvt7BHM/8tE1FpsQGwNnvIlhmS6LYPOzkobIlngw5hc9T79tGHaF2YNg
fk15Puxe4lk8C8Dtnaf2em/jxup7yT7OzIZHspAP9DpdG5aRWHUQp/5d8jssrwF5xNUQqul3nteT
6321YlU2HtE5NiaaFx7xzlBiU3UvYShcp2Xh08eks8tgFBsfgH8JaxnigFuL33RjjIx75gIxMSMY
TXlNeYguY3pfBtw4Sz13xPVrpwvFUSmPumJxi6VFeKxA6dbrdrtbKYdZLx5JlyegjdHej//+XhHb
Gn6iIAqreBE4zPfaPalNM5Vn9Nc3Lua2qQNuqFosYAMY2p8pVuH09r9/Bmaxx51SaENbBQuAmg2P
N0ehS6UNd/+fM6Ti2V5uuan7Wx9VhNr30REJ/3qjjLjSXVKs/q4Pfj1CAjvS4/qT/xnbVwhVOYgJ
VVmlcMVmS4zkAKAtFnIKce3K9dnDqYjF6WF86QAnC410RByHixpJpmnZDCtnDUilbgXJx8zLVsFX
7wFKnQTmGwOJYL/so9vsjrvk/6zw2FyUVF8X4hEVO/aFc60V4EcRfdvGOWuhDebRXFsEV4VGIQwv
umug0nzHKoRlkwJC90t8a8jTYYdZ9D7l3kIj6nyq3tWyrY0bmfbm8LsvdLb9/Y/bAiz14nO5eJu4
+1hVCT78GX8G0uGwNo8JbVLCm2skES5719VbgvSbpiCpf0xfgV0Uq2T1UsgHJ4Y+WQBr1i9XFAMo
u70AIHoT3/1WIayYxtNZZ9JBIUy0bMpyOyprDqtvUxrzJ9xxGEA8gtUGT0h0rA9pejfk2Ngob4/C
6sUj0BbyKZQrMI0OBlQ6F8HCi7KuU60Hq6mX4JMLlVtpcMXy0hf8zgjQ1ESGmzAwmu3X0q3Trwl6
saV97wM/y1ajRGmIE7zD8GVzbI4zXh2/OmwmdFIFNpAZd2D+YvZCRaWeK5ywQSyfYMl3g09Rb3Wc
lEhmyOCkEOokEe4h1ndNYK64z0V3qI0QrxHIrSQKzPUg6NQYTNs1+cc6euQwwwQWNa8qlFuyCm+1
GEWJ2D5vs8M0h9gvJ8DBR0P+RjwCz5NvEedQxW9jVgCrh/jNOQAhSCwhwKe3TKEJDkuS4YYMVhJ7
uRRrtcn49INXq2p2j3U1aE/Ohzd4a5p1AgZAfnJaxFSb/vjSUDJ+JpAsCYXxPV3ARCvohz3ozNNN
CxNy8q3t/WjjkF4wDdXz0z8myO6NDDg9U7mzOb3W9UoqF63SNo9w+dXoslbUCPFulV3LJG+TRdYn
fIqv/k2fU3mt/hv0L+ojJ8Pv5siTeI9NzmEQNbfxmrNdM4BG8Aep4McnsKySkzeyz3szPDZwXpgO
eeTHFLPJKL8+o4TJU0Q+16KZoRuJ2H6czt1DEf5rr9rseTCAApAKPe3KwccROr59RF8UT3NGfCEr
8n1GqTzCANyJM2tW6qwic/OmWvYsnszcezP1kobwjQ5hwnyVcEL3I9CEg4Oa26lYe5q2/fexc3dC
ZWtjAuqZDmF23iwoD9mZhMFbSQWpyMaeaFbQtvgUs7PO7JU9hVS1GrgYp5gMWAROx4D2qfS7RGKW
igeY87QoS0luJg8DNW2QDvN7kaaqsehfcZFWW7/yHKtOfxnk7RnJqb7Qj05sumEmfnGAmpd0pZOU
olHBLixXnjI6HW0w1CSd8A+R9OGJnSDuDK8kVwEqetsgdGCgYbTP6q6nXn1iN61HH7rdOJ9BGWua
XNM1N0hq0a+OMw2gmgIBSlfp9QCcJw2w74w6rqCuOR8lWcwxXlaT5U65V9punMO13VrxmsewBLq6
ryHwY0hOFj4g2sokKg9ZgQLHGPwgwisCXav5plFpqdMHwGRtbuxrxxbvsY/nLsNKcR9aWvgSW2GK
7DYA1qe3WtoJBH2CEHgDb0Q9IFBxqx1NHCN2pK2oJ5W7p6VgtJgOjyk+lIJKxBF99+ZnNuNfkHGB
ZG/UYe0zDC3I7FD45x5S35WGpHZs9buTMAJx5b4wsKxzfOe0ZxRIOc6y5hnuZS5Kc1doO1vRJ5U9
1/ESstYp2rcIFa4vR3yTc5VLD+6uLgWZqM7NQ9H9dqIDve1HnO1gupNcRnfGoPYWM27kdfA8kVzA
idOIaS9T1dNekq3hOTv3lJ46OQi/ZC7t6lYFt/QVmO21rapGrDT+6BCq6RPbpMEtEVn4RmpadZko
CCamJWLQT8t+T6yxwsQ7/KB7sDHzq8mDinOZFtaNfaugnAssjKoPTJ0OdO0GM4dMLw/4JwcvjGbJ
/YW0yv87yjnUbTeNDmnOyDYx680WVX5/grSdBV6e1i3CjozTEDG2wegznkkUbBZxGHKo0Pu+N/+S
zpRS0WRE+DGk6jtq5Qiyc/4qbrsaDTmzGFLRn2Wyjz+U8tUyRqOHLFe75KQMaC5WRYqTH+yFe81J
qAi8WpblL8vcfOPqxt+OUUop5u4uXfNQtLDioP3TYi0/FJysBOG34eWHJhULgtFBDIoayEy1Dis9
6HmyBdKJwhH/tJRafkW1/+qHow6yoM1VrQvBkiCOBzdl8SVaLLsCoZnudHknYfo5kOjiC/gzPXr3
oR5k4j8AoGLt3H+Zr4I+0oIfeWk8GTmcEmctC18DZlMpeubCqS9QlAE1u2TDrEkBkxY7Eb7s7mgf
ppSJp1W6UKpBwyEKD69VzghPjFISJWYrqDsb9wa/sy8HjrsF8hBjDZF/geUST3JzHSraOSu47e4R
SqemlkpyjH8XmUPs2NdEfocnIuOoDX7ttMP+TN3SuePIBEsx6Vt1sxdsc4OM+psE3OskPxg7Sl8m
KcsbxqTn1CrN+61MHirjGqmE0VBZz20cIkEwnSFDw7s/A/GUErFDjD4LvvLTBqI59QGC9i5Om5MW
tLLCwp2GR4CLxUVAKJtmuo8RvdqjoHZpjbrc8O5bLc9rcPpPFkuiMr3kvuj25TbZZSR5Dma+5X/Q
MvSXcswhEUgp6SUIwa3ZhERMqUMIaEVKvyHbk8Ul1770zuL+z+OIGnkpccnLfJjqtvO9jjgCQ3HA
Vdgp/MQkiD+2CDL3KA1JVFfTcFd+Vr26YztmQI3xSHxXpzpUM1jGTKbnR+TN2o+r953o3m3cPJ0g
80bnHQwcjxI67WHXqqK3Fqrz88L1wYoIDXqdkLr+UXTAN6Fml+E0MEsN4scCHyyPidMYBqFAYE0S
7Pd5stINFl2Il0ozhUDNaQnEoSDJOq/8f32JiDU7xxxoVBDt1jj8PShIEbUyC96YZZHX/wMewkSc
651rfIEnyJc9nkcp0uuGGg1l4dZBQiejtnQRnpHGSkJNjQH3XicZ5GMqbCPRVaDTNRNcIAPOSV6/
fdZNXLaP/PFrNPaAwOCUZ0q5CA0sbuophXyADsfB0qVLLjveMRAmJcqwS0s+PpWvm24ihWhxxzC0
aKES/H/ZgMpLHyXhIC9W4e0Iqi5WqD7oJ4wAY0iisGI8ZXlVoC1F/9IKWLGhuyTAgJVwcd3h67tM
KDr1tqNDBIkMtKjUaECLpOwV2jf7V1OEU5VF2o6avVS6qA6pcdULMhlxnklMEyCxiBtpEr0Onmyc
3EOQ0LQcY/5Hu2Fax/13KQ2la9+NGsDD0M9jS1VWwEORonLv3JoJWizwkCBsd32RWsLtAsLfK5Zi
IpF9tv0swvAVCaCt6fPlr8nWQ4KFCUJNVGBIXArX2jxB2TStH6ii60gvOV5t9t7bsscApW+Z0N5u
eeWX5ZV1nr2FQFd5X9upPTDjUKXvHA3vn8TjCcjHfvQ1C95ELRigCkZ0f4/p5iMOzUNv03k3GzTu
ElVZD+lYxJa0tPikFBKgVZMCqVyUGJwJlJ0Kw8ROqgMbEYbWFJIbRuY5UWDHByDwjtAK8UhQbHv4
Q3+5I0tAlniTI319zXM8RJWzDVGsKNNvILqMFQDGyhvgZISYkOAJfX1WVrb07OL9o1ET0kK2L6ky
cx54m56b7zbZb0mWEuCyahWA2rUOXoBH0t6bCnI6X1z8l4m3Xr9XWHI3+Ypju0/YLCPpKk6alemg
XEKTZTaT9ePUkB05zDpJT/URndPppJpe2pCBKRPr6GNPXAuxF8y6SxNUEYwfpFMYi4VTWbbxUqlg
cXqgldL4IYxSDjSU/MPoGJNpM7pPnPTAksYykJe8vTQpM3GXiuzkNTc3o2JztO4s1RN48zvbAohn
u7sjo7jFHbAAK9jXcpL23VcBJVlrRixTYik+jg9jNMxAZDMh4WYKDjak2NNltpuQzq/hFx5rUxSA
F/K+bV63A34JgJD1F4cMddUTsr9nkUKZ3beIU4ppMS7eVjBHVypi2ak405tcbUu2mc6AOiterITQ
mLMDxfMZDQ8yovdBiOL1klysiO6RmVMHefleKFX73/VBvmlGHxVjJt8cuckTWmjEqbQVe17Q+kBv
NAfApi4nz88ARN8qApQQ+zWKq5hjzOdX2b2yxaNkO04Wvssqfz+zjdKIZDk+NA5GSNJHsB7M/y/X
Jb8nQjFAd20FgVNKmrrSNq6xXKd1feqT328/bRel/O421SKfy9h+zHzXKlKnQC84Ya0UJ5mecJ15
oQiw2l71vTPKfoSFFQy0Vg8lUW4WYeGZObE1Bm5OCMYQ/mDZpzJhq0TsTESvk0MosdZmRvZhSALc
s0eAFjwFCoKJC9/aJCODjs4BshXEcSR4bexBsjaXimoSv/HOHNXnXcAEWxpqUPdIeKfp4ryrE5Qa
BAEzl/N6HJ8S+5I1TxL2GG3b8otxFcQpIItA3O35Z6K/4tLRHPn9DZB5gvez3Vnx7lv1lyu3TK/X
BZ3yXjx/lXugYhs1QrVe7wc4DpQW7Qzo3jaq6CsCJ4swnDELqFIn5fw8OEA5FKFghOER7y0tFCy3
gL4O1XkKS2pHDasIzaKuE6V6f8efijMA1I04e4kVvCfZIKRc7BTZ+6BB6+aA3RUPFemnvhvWThEG
XhRLGY1Q+JcB8muvLkshCUjCh3AyKsZ6TCWLQj48oW1Zx/OwUEgGfQhtI/qi41VTn/UNXwGxtqCE
lZIhm3ZlcFK2KsYI4ptE3AzgqYbHfx1T8zAO7jVtkC19gf7ULJwegUYBWRcgEFh6re781I7hKWF2
3AIs05LBxJiyru3harapdHhHG3wuWMZZn5BJRkCFeIV0f8JWF+LcRhr6DlZxpDRFK7wTgtVikAl5
OpX1/2gp9Dr0TYaCaBRSkwIF9iSusgaXqvp5cdLnxEVdg7JLcUQJCSobU9ivOwFIGz8phCvqT66Z
/yL/RnP7X+JfWAkWw0sztQWszi5XWEOsAPwoey9oPd7G2xQqVsTQPaAnUDUdX0wHltl4Sv5F5h/f
1gCKibIq1T5XawV+ZDU6Ep7LOqQCbiUQRQGNm3XxMp2hX/Nf3P2zqOcZ9n46UzrEYcZThoJWkAvA
5l4s8gveuRfg1FvwPD0sQ7fQP+75ghyEEVp7EDkIg8lA1avjiEnMbmaLX8EUn8cIISG1TO5EJaLI
0gbEmNohN5+6ramRMD97Gi8kAE04H65Kn/f6BPSCGXuLNMxvFRdLdMqO937GQA5obJovyOslkG8F
m8jM1XRxLfF+TpDqbnkjHn26CvZM5sCjBe0Zzvo9vrMUGCfxSaCPk/FybfdcOZeAx0whUgprMoVI
oUvLXmR9/f2bNZUEseDAmDR4NypmNAlecUa05MlFT9fnU68WENrmXNniTz8QlQWlSyhhrxNCaaVy
fhAPUcopc2MeISjnBWAr0Ge4wZKLG51jssdbYyeSNqEMXHbRmr7U4pPd2AnWgvMxMFeA3ZP2C0/L
0fnF6szhAugHwQ+w6xeNLPmEHRMlpAvVWlc+uws17nco2PobGCu6FBYGRPSIQtUkKBro3r5cJAvC
Gd/35LrDpr+QOq/ybOKL6r6cguXVVu2i0sItR5E23XGng/v/LBU2Eb7fqw2zg874iAcJWbautwi1
Y367BWxCmD8VMfJceoAyXSRxZIEEmxqM2vdHpgQO6UPjx6fegxtNBY/u2hjgwsO87+zL4Txwa4Mh
DZse33xyimN4eIK93iS6MrDgOdmyl7W0D/U2cOjGekAFXXbMkhi4mo5/gwfxeGqbpCg0qVFsX/BE
wYCFrbhmdyHy5RrUV7G5WFJNT0LVU8ga1ldaJltV8khl0QpiFRgbr2dtNQm1ka9qBYXKnwNn/2BG
eiI9cQlYJ+RvHRmLZSbZB9/EPbd7ITAN/If3zDJFwg3xIoKKFOvTOgbq1hyf/zi68iHl4IJxyosb
s1dy+d9wcHzryVph2sOk2LPPOn37QvfEyUlLEp1dAVEHbWSC3mCo0/juAoRM76+5hCTWvR4gOnV1
yNIfCN78+EU2yEhTF04gYnPvaMqxMuXqoU8q1DNuwhkIemD8d2U1DqXQDCsPkpSEGBtNAtea6XnB
h+LqmHOZuHQjuwzghKRX6d6tjPU26NPHI2cYBNffbuWg0bhmNOIjxbWl8NDaYpSUqPxtTuTC+04v
f8//yWQuiYiXOh3FFkaIJUZvW9a9yE3FzwgGJvzCrzNXUdUHSbE8pNSjDhBs4g/nUS4Ora9y+ZDz
mbZMgasvVEdQ11lyS9XQ52cqaMcGIv1/f83oDXl3cLKWRaaz6OZwwH8QZebxuxBk0pAemqqalx40
ve8HwpfS1enoC2RlCmBWR+P+2cGbQeSslR5XFkK7kPyVrRh3KGP2Av62F8XIgnqwLnYcmkT73ut6
M0TWw8WS20QoZVIJ37UHsx0lPYkNK1Gp9B4DpenHoPFQ8wRGcRwRd+2Ym2cjQVH76/LgVHFFOnPB
qjoNbljGK9rfpK9l+MYBLpp9Gfvl/XVIhUwgwhWX8JfaxXpg064MAz+bDlHth8OzeIkyOpC8Z+Wk
cTbCX2Dd5lvyjcN7cguSC3ZGHo3xKwVvkpyonEg46DvutGLdvBk0NNWs2Z/00eUjSWoYePlepyEe
VnDA3tpqShRkKNL7fb0XMNEdVX/dafdkBg4ziBpjQ6hrsxSpEQeLfnr12jfIbztsP9oyNIQb/l1r
OjPZahadXSNE9uRzhbRSCYNWlyD4JYD54UXnmRYA918XMcgQVVT7EFn9uSMBG31COghdC7PEK9bw
AavfjpfnRcPbzQtxKgU0Z1UzQroStwqDCxjDK2rahX1VjrQkxZC5VzbBnEvR3XZQlBFGShvcOKAe
K/5jksBTtlRerqps9+NpBvcWUEvdl+BcwsSQWBSZ5VgunvvSR4hfw6Ybe8ifRZ9LF83dDeDyAWKK
lQzdyFGTtfe/Fk0on86HnpcKI5WmyCEC+tQOtBsAarjbzcq2M58eJ8L9CvQQ+x0PO+mICRf9V6OO
Dzt7GD2YVYEQcbquoxK1kLl6rBuzbNnrHC2zF91RwZkP7BiLC74WEgzIIxLVOt35D2LZEOeoCgEn
zRxsN4OnA8AlswtexaqcJxYj6swUHDJhfM6YHrPWb4KXnwD3/OxX4xhR7JEN+EuDCwQEHVnm7voD
L1Y3ZQgsuDgPSrmVTjkYZ4EcEyMRYDJ6tFuxMvCU0xvVoduClzpoVfSadtaVE9f5U5StepuXuYE/
DN+Sqr02/8TdFP+VsJ27YU5PXsP14aIwbw3XAuTqkngQFiZ8jppCEn6hxH0HuNjaHCRCZK/Kb97Y
lay57XNe58aQ8ctHGgjhoI155HgIDTpgPs48ZNMtQreDdaL9B8MnizOZ41kiKk1GlXTg0ixVATkL
s4HFLKCHPLkp8NZysHVoXYr1HQGdC0fKPmi7LfQJ1l+orTp8a9Su1CHFibp/nNzAKB4+v1W27kqE
4B4fj512Hg4l+LHJwGkO3mD8LfUsAwdIlPYgQRHMha/EW0ZSVZYHAjIq/T6pzVz9gIXbMvar8mrE
CaAOdjZ25JFlTcDUm/AFuGXjseolgSCGKAgujrdeFaARkXoYOAF5oh2U51ELYiIb49grH8/S0UFM
4gNOeb3ZZ37a6dFpkDeWrxxEuQnYl2yKjeN5vnTHcM3eHmLUAGfxzixiSbjJwMjRv/cD4Q1naB4v
bzZu7bUSe4Mu+lp9UAAgSBvuatu1SrRw2FVGBq21APVrvHXn690F1QtwNAPpRHZkVzIT4+TGcQT1
hsFwqoFGoPSt/MnWnvNYgsRKhBnwuBKzPqvjOEk1G6VNOdIENyiVc7IELqrTeNMvhzplyhlGjIb6
EUW282KjUvTVsgcssWdMYGf90h0oDIzvdI45CZABjrsHwkkG1IKVH4M4NXAF7J8z87/zif1Tub+p
MmzCzMIjNLSCJ47MnK44Am9oVp8u2rzdSy9FT2kTll5OnTS7CLHkk4JXVhkHlpOB2RrwWrlIaXC6
Wnsp357fzIMkrh2Xlq3EXedIwu1h/UygAivV28lVNU8K9C/vdK61DFIFNQQOCiIIVY4UJhOvTxA+
/7Jxaw1t6KqhrZeEDWJFpSSnqO+LszSIUggkFBreyEbKzeX8dUQO9VRwRn9OkmApaXJd2ajJa1QT
dmHI4i227R09k/J/nzPtntU+shrxud4yBoerNq64Weu+F1oGMLKySIzTa/EQZOFUbuJ8lX+DRXbr
HjjMtF5VDDGHpjKZW7nbymfOoOlkYkwJkjA4XV3R/g5dS1YqxE64l53J8RWo2NyAZjIDRw4qcucl
Ud1C7SoVszYcYYJhuRFIvfc+CDK7lwkd/+KqYHax12h3eK4/cOqOdb/EiUoR8eJiQ5u3pFmcajsz
09Qcyej2DHGIX+HLSEy3prL0dBKGmCqG4oB1vDWYzg1MD9L0bNIMbYXXd6KOOKCs/wZs8lOiA73q
nTWbSMUNziLqGvUFYLd7Pizj6nHYaLgRdgMI75QXu9DK1Em58eMfdfVkWBieXKkbstHgn8wxwtlP
5yk5M1iOITSqLMKUHqLQhwyritnfjgd2hvmOeDD4Wf56OXCtGSZKsgJcawJl0wbSCxJN3fH7YXxw
CMktrY/GXzg7yllPo7H/cGBlSKSsJxLo5rVIyRsvXuEDBtMxThW229JdChWbERiq8e3wsREcvLif
EDkBE9eOC5ejXc10QqWZfiwniZJ+SRGLKjMx8rb9SWXh9TXoaZKwTcC7SUy7COvOUAaX9HRE5k7f
UEQdK3hCOgCUweCGIP1FtdIQ8js6j8zcGnOdhYabuhWHkYvRpOEiNN+UwwCF17zEVlGQNqld3OoO
vOGAHzLoHL4aVsfgMNG2pXfQgNVB6mUptQU6wQzQcPG250OmeIvYMC8mDiJdqCMTncIIkyOiU9g8
+E4uZFS2S/UBLmRfmLi7k5hmgc9TkqbJqosr5W85kf/kmjI2lB0YMK/onf6wi+IozMpj4tBwjH47
u2pqdXj+7gvbg5IJrATEkzDBdEoVJE9XIpoC9y4U4YLtYczGI4hQRDFstPSbbD+hJtsJuhnjg2eB
CGooapbyVk4vjB6WBdaFWXfwEMcwsqD2lNqU2gtLsfS5Ik1YTk4frZp9fBDmOSaNmfk8esdWvKUP
e/J9UHYyWUfVFu6aTm7CxKL+msQrZo7D+n2qNQcvpzxJUmgYccGtn95xxhJe2QJHorc4MFUIn6UR
FXam+De0JGCex/tnmZ6u7eU+4Mq54DFuRwNvU9zIQygg+XFaJtuoIhkyrVqZR23uapDZkWUvBvOt
21AddW7ZBA6otbd2fVbRCC8H8MBbGaSIEqoDJGpuDbtZine1cw2CQde1KMnxWZNY62hEi94Xj8lN
Y3NeoNwyR76QDBtv1hkKxpNho5njdvT77j0FDAv6WIczHHsBNrSgRf7hh1E+0h0L+ZybhvbK2mN0
qd0mL4DkTIni7+8oFaVWTgZBwiStpqRabaetHtmCE2GVvdH1dEfTiC+HLaoWDttBPunuFc+ByqID
vgwKq0KUToQQJJa8b+Q0KKQcLwK8yYcU/Mv0xK3XZJhXpdXL/F70c3qQ86UOPqJmKvzruJfCe9Nu
OUw4sFuRPqyeocZuGgyAx1eEgRumpfbEqdO3adLQah8mTjlULNYX8ZYfiC6X0Co4tKp1QnBD+mxy
6BeBOpJIht4W6NZDGGivQO1Tp9vkvTLNbOJdbsOv9xRcMMWCJ09rBJo+BjyGe3efo9UiSulxMHLF
Rxd2ylAlxuQsMPWp5QIRngdkHxEfTSPTXdofHxhtefpX4gtzmZS+HN3CHL5qQOcPpnVooS5TbjCo
vfw8OCxMbBFMnmEGAMzKXNbRlAIcw1E+UeB9TtgMRwaCdXmFbr/xP0otoDiR0QHYzmi4spy/Dkkn
lzyzMGPn+TfZz+EevYrPxDFR4PB/ig8Q/MCNxmCGIyPXugxbYyfc1jjOAculiwMrKjO2KNi9WQqz
dECiVFnnF9M1sne5w73RCNh7RAbO3PIX3FFtrZqNrm+wzBfEDeysl8PxgewgfmpI5h/rbk9zJJgf
TJcC9mvSFwlFOz/D+jKt5ep4CWV8jAENyXfXqYxxU9+sXLHU9yvZehI12CfAzR8CZL3amlad4JE+
zZAMjYu7uuDIYmQfC2RbxdqD7RfDD4QRio+N4BsU8pk2wqnHIU3FhnaAHWYFoVMWTBATWZl29A1T
dF/+rkVe+bdeycr9mkCO0P01P4O4nrQExHr4o7Ho3lfwSnZ58eX/p4BRYSay8jKOIxahbvFl9Rwc
DXc48rhM66nCAgIdGakaPxsdcByDRLbLrGfSAeT/2TiJuGLL/5a10dhE69NTwpd3LmBj3hRspmOH
Mi1KhrqsJjlJX96C8qi5oMeGZE2IqcTmc7nE+sERsSzfZNZII/Iy+loxYwVAYO0DPXJCgLJJf4TG
ilfzkXNkcKgvuZrh6lNOczVhUobRHrTjRB14U/Hc8s62zoKZG2zMommlVhiOzXRd9r8u0aBNkWj/
/OnhfK4EJK2IaPcwbtSBiT+lQG9mKtI+BTKmzsiBgPInMTATPteCnV56zXI3Dm+GCVTkdzUw3aCT
2JzN02ent+eAryFl4R7IdID1fxQ2tU0lYV7Fi6TmlNt3yQcHhW5lSlyKSvTFFc2orL/zEPRm3zQI
MGBk5wUCkM8YJ5QVvMZd5IbwSgXdIJL6PM203fnreT1fNvGKQQqZfdYhnVkDmJhnVry7VcCjthdi
1UywiDP3ZcPTCqssd84FdRjivxzTIBV1lNC3u0MH0jYFNIhcA0AGob65nf8zrJCshLjg18yir8Hi
CUJRq7+wHOYTz1oDBWIGqqLktPjYH7qanEEat8sy2qjMFp673UDBlEkTJaIaZyhY+dM0ZXidnrUg
iqnvcC3bqQ+nbFEyAEIUozbR9O5cbSFfUHu6oXEklUx9avQa0j4JFyxynsyiJbjoCfTOMXHlXfc2
ZTtmeB5/VaBLwu3pu+jXR0HuYNK8zK9z7/RI3mMln5bOnmq/OZBvYqh+XUpny1ttwFNA5+MwLAQa
mIbXCJ0OxKrBqJYvgGnimGV/JLvewYwXqLjFZJ6VTgrTTr92HqlIKtyDj/EzNjnoxYqOLMQ7Blp5
bvgpM5VAjKhO6WeftoCV2ffQL0K7EfOmBbbAb2nBDgiwfEmuEo8qRSp4Pc3RpmYw8bhCBwIOIJ53
kYW2mJV0SeF2UOUhixG2wLex/9VBjPQLE0+4KCOMiWDTkqCk9uwB0gwXjgDXuFuakDGneUzKACLg
2ZFoZMTwLiCml2b/apJXgc3Dv9i2tCX10vDcz4sYNdJum01MH83lLLeq3WnUDOsXwGfZIlWDVA/d
WJlnTprNdbmJ3kRGzCfwKoqUdoG15pyANaNy9agv1jxoFB0KEQx5KewSUkvmmCzct1Ht175PvU7s
9aD3Pmknu8FgTMTtG78rmDcTNEFT0txz5Eyq65xpVblG8p5tvXWPdv64zebZ/qbvi7YjtCisRVad
ys5UH57k72lTkQs8AQibF9HEDzuRVmBQOumIjzZqGZS0Yua8Vinn/s5HlgJse3QKcsvfanGNNmKD
7feG+iBnFLAWGNDr89bsqhVKMfNfjsqS/bVqLM7RCTN1Ae7AZw1jRetLz+9PmIBSZkgNBYqsuJlu
rCspjtoVoFsUDnegZNbonnzWEzQpN4ibiASgZhV6wFdX+a/KoNEw4XAwJ4CY3n+00qo4/LEv/Dm3
IZweg34vK8e0t2+84FM+Z2S5tURWZly2aHqDzZn4/hlzMV4tZX8bh/4e6Eg+Z2d41720ZeVgWjGa
kkwxLppU/CxhRCNLjC3bsTrMNA824HqO6ZIDq+ceA3bbDTDbntdTamqnM5XXjZZ0Iecnf5xen+ZV
txZbQQY/jEoc2ztZ6Gf+Q987F/77/uLQ2aFiTV8Psk9n0KDbReJElb/RLMbSyRhLwjWwohnQ2Qei
WikXOn3J10+t9rTC0hN4UquJxYdCv3qw/nURXXeHWLStfGDjTSUJQDojVgQRX9csYvzpP2pbh/pD
pdHiFODK1m5WreSFd/ztUbJ4l03jFk+egjxFscfSD+ovHJtnozcy5FN6CtHCZd2gDYP9PbKk1Lek
+tibx8eIjd06MeU0UJ7RqhMLYHlvW60s62r2LcJ3H7z3io1NjQatn2xcg/ZXsIirXEj08UruW7me
Mm6xKOjtMpvX5/4mTOAFAlqmD9StIQ0t4bMHsGCgNTE3xW2PvJ7BNsp6XBMegQTsP0qmivJRVuHP
sa/swKZEyKoBf9Wr4jhL1kXckh5/cQIHKGoISpR6lvcSOyh8XAl0RjX+WRl69GgYpyiShYLxOkQ2
1ITxSMejZuSokHvY6Y3MXwB+xO7FyFgDY/Z4ojrO5yZ3+FTG4RQAjp1+54Z+nucHEM7u+7l+UzRF
GJN/Wr2+DmQPMqf/zxPkc1xmDympAgA2srDRrZu1rXbDNB/FD7rCPWs0NoiSArdpRRxm9Hsz3t1S
zvGrWa5h0iMxQvW7Vt/4zDr4ITyJ0AfT21YFap/evq/MA6SCbRLMZvV5iKyu0/ssfGrz5nA+E2i6
MHBAC1UJstPY0YS/w54kSV9j6UJYJNaXVmcg3ShtQcK6luEs+N1elBe/H7OLydhvMTG96xhEO15K
s3rkH5khdt2kseJJiqwq7EoMXqpeHH1Tn6IpM8Yh5y3t3S38Nf5D6DYyAJsrQo2MPLkux1gfilcJ
Qhl46qLT41esANnDO/Hco7JSsxfzEJE73Rr9BQfh1YcC75AIvvkrAVHh7WGcP7A2Uf83z3xEQSCe
hqfsA3acll/eKiLt165VPUwxixOyKVweDd5eNsrlsMoT939sOWXjurJCZTrXySqu62/ErflB3Jmi
lgqLsPtWFac04eCUZFOF0BRg8FTb5aAA0bZSKeY32x6v4P4sCNyYgHjVEyxBNg1NV6WN+HiHRU+E
qItSlym4t3TuKB4VISu/aB2gNbLzjPZXcs13og0Kl06Lqao1X6Uf37cI1TaGxsVDkgMByK5Y7zVr
sQUMkj2e4k9SinS5VBi3FRugyL+ju7wLPoHtw3xpLX/UEt5gY6YxqvEep4H/f6NhCGTLeQ3vXgbt
3X2ewKm3VYPkM7kctjQyeNVa4Xg/DaMEn4BxmuVeqyE+Jnvt87ZVrGU0IabnttboESXg8ASRPyJN
5EIlDvrc0eP7bivx2tDDXPn0jN7vJTWrmh7x8C2wBXWe8wb1HmA5s8PnIRQt5uZYHLkFcL8EKjhD
HV6hnj38hNkkslDfmbYfbNN2c7YO6sz/D9yZLX9FGxU4iiKM+Maz79moO51cfhIbhvtMOdkaVgye
cBQXmiiTlDfKacElJccDSi1mU9o5/W4psPsJE/NVsVeziRvl3dZE3xYsJE52K9dS196y3q6T53SC
a238tyvddhB4fkRrfSgfduu55DvIUvWVaMw2LmIeRpDUgYG+N/GK0Nva1BOnw7KSYZo/rrNCz0ER
tAg2YlpFk+vM6lQYfSyBXokZCX9Jlcs1tuxqBE35zkLl9NkiFwNzJAjpfeTnErxrGLLvbBnCNTt/
Z4iyu3jiqxgy5kya6VHK4u9WdOCFSNS61WO859MfTShEuI+sf+sjVaITINYNXQMSAjZeeC+BJ81N
UOP/xIpYAEDAQIqFZx0X+2mm6u/8+0nkzUArAwje7DRnFtU3LL+3v/T3qeeq8u2ffq2GyI7FaD+p
eRRN/WnDYQZmJA8nUU0fmOlIh6kkKVRCjwzUgKBcOusQVIgK0sGNCMOs8ke7SL39EzmiPGxhExXl
iuwqcmob4rW2zB3QVeMW7B6o42za6xgQsPx4w1hLTdXXNwT3KWAaIWKKQ4vWYg/1u6N2buuOAyMd
IrZp2F8vAkzubWziWH0H89p4V8/gqzRegEoLbpFa5rW2Aqds7JqHlAhf70HkTNHHliELVzfvtVWp
pRcaUlkLFtSFKgXUj1o0DyLhW9UUl8nr/512pzKYT0R+2nuKNavgQ6vYY0bJEvyGYAbUe5gXw4il
rBZuq0o1gVMXL3kIZG7SSTkVJ1zHitHUCkU+U+PqbMdgEttxFP00aAblp9BQqPJMjpa9VtxkizD7
yh4q5EiZTNqZ0RP4H0F56+2QLz2E4sGGUisxmXKbCp52/7WMTj+ztLipOBuX2VMqpsEsFq5hmaGL
mk/rkX0poU/MBnNNS1p71mdBWbyR5UsTngcvYmCGUJiuBUOoZLBxZhhN8K7cHdZeUsRi9WtvDW6a
8PihJj+pFzVhmsUP1aIJk82snchWtXd4Dwitb1qSHc3u8rzlotIgNvjEHgBTe0UAy8SoKgAVwj/X
PaX2rEE+Pdz5n6v4GeaecsWerNZ8vwM5aCEKB38bnvMU+bCOFZZphoCFJc+vyEqGI0M9K4v//pRP
4aXjsbIxd98qPtbux/103pT6HLpR/tWc6lEIP3txeT03cHdGVs7AAEG99MyCX0PpJUbMLgww9Hzk
sOzcWrsos0FbWEM826jAyqnYLCZuN/tPkex1JiMfDUnLNxowGyg1t1vjEDXCywNuGJeAMx01Uqxy
0RYHVCa2LZw8+65ElHBCvm+24GJ+7sUZ4isitO2dQctx+llgsu6ZtTmvn1R/jRSkx0jWUlKeUPlH
4P73RR5Vb+IX7ztvYlih+/VAOP8jutHz/RFUBn7n3ozemCwL/pBcVWAgJEW3A8lzlMt+DYOUT1rX
YgIz69fIvjPG7wX5+Er4aMNQcXd7hvutkI2F89Q2tAGc/7DxrRm7jDn9rbApezCnScfc/mjWYpMn
7L2FOlDA6JR98UqE+fiokpZuNHSVR9/D8/aRhX5AXqkTecSSNVJ5S3tLzGr+QFiXbyWZ/EWk9fLK
A/P3xRoSx/IYL0p1QCg7oZ/GYWOeu1hhPs58YXKL7u8mmB6sZqnijWyOUqAErxCtWqnXG06EnmjX
scmD1HDh0jRN2gX47d4SjrnsCl5j2+8PV4AKbVUeVRkKd9GTKERFaD4oxt9vSFgP/depuY/BpZDV
qDLJRLsIkPrSNsayOhMEc8Meyb2lBT6E3esv68mNIvRk+ppLsLULwlVDU7IdezyG2d+ES8cxQ73p
D8cPzr/IGI80E1Uq6uYq+5bpJzQBXolCTNUzwUREnMOmegrMHwqWjRD10xzNOh0GAlUShN3694uz
xsz0zMgK5LQ1/hbqvBeBxKm2Rj29NUB12lEMmQv1X2XIlEafVU5utsW8oQY01W/ShJdAHYDQSl24
jFbT0YBYwjp7thve8YOZzm/kjODH4VVuU3GpxYNc+OLPKfdyoydvwRDU4UHOEUK7IgFiJ5ePn/DB
Ue7joEeUIzrco1j8IacYKlbS+X0RmaAAy+vPnPaOHbdUpZ6oZgsoW6CzHj7NREAH7HnH5c1OGVCG
yimaM9ghJ1I6C2KztYgKeuJNfJ24XK2uTHWNH2t5Ze9dnUweimUHeBxKbhTuWJNKBkff+nJqxFE+
0DkyjdxMEUpmKlzvhMmO3O01QPZ+2hm0jUWkeoLE2s6SZqtf/SE40PHF8FLpX7nPhHCFV+fAP1xA
f/zm0zdcUuSbt92TNgNlGtEYQN1lmq14ea7Jjwr8njNBy0Utfo/4chaZ7drY4SCgpKALrISkrBXn
q0zYqAt3DT83kQtGoEhlgPNH44hFd8G45Yxsq7XBh5YRMjXN/8yW0CAwmG9HTuL1FwxlzRqfiWQR
leX+bwettQaVdUVqfydl6Gkwba29wJ331yDNbOWWv8jaa04DyBaTnJzmPbNXofEL047zBy2P2M6x
sPN6Fcdjx7rLnUC5kZhY7+4ol1hGCy8QEQZ4NO5nLP8I5nyoZYYywRsqqf9coQrs2KO25QEN7jz7
Nc9v/4PtuOK+ePuCzWgFvMFMPwbuUM8Pdp4oYEjXu1sek+s94RPqUjSFPUqfLf945cr+bRl6dCPM
VyBzLJ5/P26MLHcclJtRc7OmNY6fmwAcIMswKx2NXHWZ8UVrvXjpb/Hq2u9mgO9b2hUNsFs4rlVr
1MEdnL94ueyB5jKs3BIJienC9yPCbwPIhJOaYMgCq2cJF13OerTrRtNC38ZfEu3DyF5gZaE60wG7
EE1EJB7p+nZxEboCiaj2xuGDQpsR1krSXKR5Ie1/oYtbNqavW2pYFKfk44aFnDLUM0jgfZyOBYxG
vOO4f6YoPahvOh5MmBe9TVkYCuBv981X3ErfiG7zBkvOmbdQekIYOYdjMv54pTJ22b1oGPA2n2Lj
23sTKokklyBe7ktHHrFLdLbR4dsCAY0zX9J4pZ9EU3fHurCU5RwLgqw/LFh8uQEP0p2sWjn0Eqqz
zohAZvt+9LN28lYNqCDsfCrnV8snFsmBPOWpBAus08I2CM+ayWLYXloDgt/lljylJ6mRm7hoXaA1
p/pSu1OoBxFK+bpqUEylY7nngXY6DjC1N/nb4OIrVb/vcfrMcoA+ZlaItYpKECRQb9S1VjaKhTys
lMLFIvGAb8X31yQYEQlB/Uft+Ny9XiXLzB2cD2x24ZLdJM1v9BgMrW5NBBVCM5pGbQe6m5ggIgul
nv/q4j8lhbi+X+BLp0PuFOX/TaUiasIreTAUCuNTM2E1JcGV37mFIkuMQjgIAAoOC/FEE8/uZCm0
K8j6APUQ2BzgE6commzyu9An0QN/RNe2sWIPo4q0vCppoX/KopqN2PoefAmkiNaMyh2wSuwqPI9R
jQ2XKiYDSxp3GFpYufmLXefrMmOlgoglGreBZz2XChNnF/sd28T0DuHqhRPREfG7EsnbNGi5Hq6/
bmjAuVwwhqn0cgla5Exn5Moa5H3gRxRb1iIenWhP5fsezOSxSA2tYBQP2Nf8VFL2zAxSAV54Scc9
pRMZqnRpN3XYMFsfA7JpnjIeRC8kLm+4nt7tk8xHYzcCAYQPjmjNyOS5HQDEeT0QQCu2P/BynkAb
IwdiVPbyu8SVK2xMMd1Xm1Msa5hgyH0l7WawT6/0HYCMulxhsCa0KU3cZ2lRy2zGcd1hCjEQiT3b
vF4C7v6B1fFphszMoIv277U5faz9ZZUqz91rAHroWKyRigsNFEo3oHFRU22WBWwTnoKEJcDM8rvq
2f9cqXPcaPLBdvTm2oBbG/JzIkJI8pX+7eWoApUjSa57nQD/GItiaE4fjLb7YulJgTktguXf+m4/
NV4LqR3K4sVuPYHIpwAG5UGkebBnoPCtnoSa4q25Qrj3sPK+KB57PdVFbTwaw4N1VtfObEBcuJvR
IYjeQmBfUcn/g2SXPSG9a3o2wx+9tQcuvAnIiDP0KkroJ7Y4d8rmIy/gyp/FtX2s5ObEgXVbQY5E
2Qeq8Zx7qmDNTGrdQ3l8hqzBl6eljxxEu5sWYkrlvPTN7Fb3Yda+E7lILrXIcS6rKMCi5feyB9Eu
rZkvVBrTt0AUt1I/7OMLtXW60F5QmtH0bzmrKHWZkLLv3HYUey9RZMN22Nwe3AyQ3071PNR5TIVX
oX0POybkkuq6jULGeMXjZixRzUDLZMqzrDLtvb/ROz6//KrLg2+17s30mQgj5ue/WxjEj7b/G/VQ
ndvnTXg1U6rQQgiKlUKJX+65M/E6/xbwddzBZ+swtHp7qPAJ1+38IBHd6iw9cXvm7mlbvYjK8gPr
fBAjMMDrQ+oTrhlpt4k5rHbxhbYFVw3MQj5ntIOyvMHr7iCFsO0+CSSaXXUpwU7SP6VowPU+TAle
nyLE+vhId637PuWO8292WBpCezivRqxY+WaIIYzFYuFhz69o+EixFJpQgxB5/a+wdarT0FHVRADg
EXNh0Nu6/ACHGwhiJw1Cg0TdDy9Xv9TcK/uXDZyrCVhCOO11Vf/repQile16mp3j7zlmt6etbTCN
pUCcRI8QjQ4whwfz2xhUAM57iSCABxsPpLy0hKteL6342k0XhvAwcQMocwE/8lfhqKGGIyShYl1F
nHjP+eR3Ja4oOaZyxRdCMi9Fl3Qw7IrdBujmNtME0HYlzkFj7QKCtj5LD+QauPyiYVookNBBH9fY
vROiVBWDpqwBrgJjpaUDE6ioy0fFeNVHVYWqA0SL0cV+t0Po+RgaDUtqRDMMdy93pRZqLoex4/VH
NTsxBC5P37SJ9Ebh44gevZy4kmpNRVBDl7znsM980Karf7NJmfc6ELNY8i9S0jLDXfFhsFEy/MbK
FsirioIE7iC2frG1fTpjTVhfK2e6aMsHUhTSF3F7j+e5kLBnwZ1EZOF5MFt4qHoKOMWErTnOmpqB
cZSTnDYO2+RuCRo6NuJL2SCuCdFg292Xc7d8S198z5zeMKLGQu3BeRTI4D1VL+0UG0SuGJEcECtf
AFMGoESa+aKliNBPcYwwvl7xJPV7Cp5/FYo5CiiL70ZUZsDx7xZhiqA4hDag9TnJWnq8BsD+QrTD
+151EtRzym0lUyCybZtknTrT7XxyJ0UgOwXZR9jqvsPYvUR1hvnuk1Z5YgajOPgONoc6NtNTgjwD
EJvzPzO6JHh5O0nJSaturGpIEitA/U9TrrE2EiRfaSNM9JYSIS235i0HYznGfolo78X33Atd9gc2
4NSIrYiI12WARxZVC6daUugwe5BjdWJYMlrVVM4SApAFT+q8h7t5XG5o7fwGbRKl8o4llDi9XSxy
OTNkDRMc0loqX2aqYyobU3qWsyMLkJvwYLmnMBlCFNi9JhRoJTyzY1SO8WevuDJhWq19jqeN94qH
z/aBs5aay74nkJiuIQzEwANWPDvV9Sjnfd/ieC/Qxriv1f6H6H2HPOmIFp9xDoKTFPp6IBXYv7MB
Vm3tmpYrmabWT8S0oyESn+Q1OQct0nlQWnNA5PuY/P7hxAj8PVW21S2ifwy4qQ2SSRe8Y595FEFn
9bz+hkXGYPqb2Zi727GWrQF3V4+olVLEPlWj715MkjzTcd12pavo5n4mo9S3SFfoqX5TZg2pEnHL
FIDh2oSOpYNFbltSoYNkkGK+ZvnbTy0gi27RaNhTa4hLk2St3ZFnsvQDBSTSwFGa4K/ldF8zGKUU
JYEaK7ve0kg5lWmL+OUMQeT/cQ2iVXSwX859XoQVZe128DpLJIV6TdWSTWrAjZNXEeEs/5i6NAP6
TjPYk2Jivh/EcNak/QBrkwI+p283zGEcvu6bSM+LkQAfs4lnyCoNbG2r5z41hVE4aQ8dt9wnF2Ib
gLBt9ML+M8XloToM+LWCxZ+Cgd9ZeDZVcr14HZGQUSv7sh8r054aky2UbjvYA9jo9viTQtKm9vM5
6nsGz3sCbhPIAjnP/ygTwG+e6gL9XV3YLJQR6sdR/RIPw79ZOsAIjiL8EaUeG3OFVx1UbT6pPvuh
yfry68NEmd/84zJj4DcC+ccPyInW7lKjdF8Jp/O9aYTmsTGzSK1HDWdnHq9Oar2fzjw+JjijE/Sl
GCaSWhkyQwlbROGU9mB7EzOBsl2w8L+hNlrkvKC6VzmMUqVsgCEG9Pbq26+ZH03eYzx8oqKCBKR+
xoQUHO0FFQ5lo9F7SYsRJHmALwIPBXF3ihSEM2o9LCAvelpsx+p0Akpu8zqD54AUvOrprWcTVhfc
uFepj/enPMn8BcxdWWyjNgaL4NvtEdmUC7QtCWG0KFC92ChUdh0hHbYaCvNeDAfFg2ZCs2IuXHaj
wnH6fzKv6GNVXnaPkk1K07wumbeMx6gm6PqDdkIwqvlwnmAxoFshwLp/M976vryJN36shdrnx9Pl
myiGb1KbWvcwDxuiGONFWznse9lgVGh4VS509PLpXakw8X4twDXb2Nhd02r4JLd3Tel4q3dm5rS2
LHsDwiw+IJLsM8HPD4JNyTR/kEjJ/EWgmRexPBbgU9WQab9aIbf5JF1mUV5H6iYnRAGS1HYGskh8
Vfb0vJjts3IjOIm5MpyMdMTX6wN7W3mf5eG0y2czE/T0A9Uk3hIfKYCh0eq9NhMSW8b4kpnd50vU
IBtwIBykKItPEfT9cRwMd/WlqGOVB0WFzzzc60wtkhuM9XzwquRBoV1bwFS0w0g6vg4M/bQpyNTT
eczhXVZJlgGlQEnd8wWgUFZhE7CSpT99nMld+KkgkD9nxxaT1MRq48E/5ISZpaGubmRb7a8XxABG
57X6Glha83n8+KIACuz0CvG26C+skdGIEBdxJ74YehykI9X7r2yKEWtxQ/qDqsNz0k+Hzd53VfUm
bwP57QdE7Bh3FQa7U1kBdxrLxph0HW9YacA0F3I1ZqG2y/0CULpOcPEgOtupDUoQcz6V3osp6u33
IxydsbnDg5PEdI+QnfmytHjES+OzlFKoVwiw9fzt/fsSmjEAOfFxIyTecAKaEaulcputYrLWQ4kN
P8t1/NVWzEljvgq41iUe0KewG4AvCy/8vsu6hEmRqCnWlWD0Kdk4KBuEwbGSg9JaFjez0D2HzzRQ
g93Xy7anC39rlFy6cn5VRGNUt/9fVkHhKSxUxzWwlfTNiib205JRF/g//osDY6FOhkfVWZDWpIPH
talX0UXd6vz6vS+Y8qGJ/DjfCOzopVYaMRpjLFYSH1MsBg7AoSqEOHY3nzm/vp24DvPQl35sCcpo
9D1ujumFpSHu8SPQiw9C1RHePDK+dh6R161aEM9c1RScN/1h38vIQTUvx1cVKmKykCRYXTSEIHjM
3koqEpqQYkqZu2TUhnMLgjT2XTkI/0tjZd8PLu4OLMWDqdMkcEo7QuD458ES+9mEvDAkdeaFcqcX
Uuuky+zdg0OrO0fn1+UjzItOoQUXXSXruIQHFeb4rjEOGNQwT4pt00y+bR5/h5ztbP/t6LQVVzBk
ZP6aSWpWLXwG4iIjoaSKF9TkH+ybEdZx+kSqGZmWvNA3vTTNQhiRCD19o+DQ042DYRNw5jly7BRP
JaygYYIQWOSGb2FcoI5HQ1VZhl9Bh6kdj4yBXcQfP5UYBenFizbd4vXMWIyRbiUY50DoqmuDDOPo
Cq5uLGPgyjNcAbVfPCNN6Kgea9ZglF3S66QZt4WzLU+Y3cw7Bz9mMyWtyKbNQrWa6Yo0cuYd81q6
2RaXsmPZIrnTHytwo3g2GtLOHGTT/Efyv7XxcPXbI63HhRAIlfd/fpKOKPhg+ldUFlaWDWeubxAc
X2T62MtpmA2zraTK57theVfwDxQhbCagTx+qHeZgJ3yQ6yg9Ba/xh+qe/PGO8cRP0gfdyknbWc63
vOoAzVYty1xqN9aFMkeiqTsUKdoeaTNOtckkaGGKSgdTrWcJyjS/jmbq+uhThejJj6MsABsUfc+i
U8PMe4qZEdvg9Kkgzqw6oZWg9D16gPJ+jkBPv64E0dfAeLGyQ5rlD4loYPv2dHHehOPORXVU68KH
GqlqehbQmbbwF7fg5dFEcpBRso3sPabbT9yzC7eL1zINP1M9HyRqHLJ37C78N+Lxo/KO6KYKDLyo
qpxYdBlg6yFfsbOweF+hx6syUzqod5Ntkr0kh+kWBg2rLsjrn976lX98ZiOiqWpflBUX9tg6P1zt
Dxba5ki3iSOVpRg1HTIe0Cz8ae7q2sayq+HYiJf5rGS7mfI07LpBNBTfqPqP0Fb3Mc953CIqNTdb
jqk6vOOqM4jcJblEvXoarXZwi0Xx1mQpYNzHalZFFVOO58+MSnJVdEkbygXKnkM3wNCUV3arCEUu
BB3jWFIcpdTHFh9YAR8Ic5+aBhG1yK9120W6qxvFFwnMtqOJdVcZQnKwcXd1babveS9MBwknS0Fg
OmFcGEZXeRs6BzNgF9PJWdSaUL19xgSWCbA7lv9/8s9HHd/gBRRC19TA3xxyYsJgidPOkMgEmtqC
PfQ9+Q/1076csO8G0F4WVwtZEd56QH1VfxCIYkayDP944AeSiKPKLv6fXCkqbyfIPPdiqakyiNmE
6dctcI2VOUz1ylXxfbkp3cFpBEgo88dpoQF5GTTi2AxaWPJZDPJ6T1+g5Ui7IWYKCoOp9CezjpyP
sahtW0GwN4yh+9HZW7cxusMc7kBzGH39WHbvixjkqCMg/aRZ/pW/U/a035Z+y4dR1h1z+CN3zOPj
6SHqD/jVrxtJzF9mJKDd8yu2Q4dTNkhxh8qHsJcGTohmNwfTZYZ5RuqbFLozz1hTRYuUywqs/KDc
qYbXKfjCagnWWIabo0X5qyxHowtkD/giKTROmkwsZdQ0C2M4wa3oHqveX3LZtgsAgGJTJDF2KV/S
b3kgYoaKJ/mjvqt5hMVOUFEMn6oGJ4Qnoi9W0fv1F+2XB4BHv2c83dlf2YRde4dOcIuJNA3ZZnV4
88WNO22+v9OwW7wRaUhbKfVt1HyeY87Vokrx4BNviIg+GjE/WLukMvU80YRYAuhH6rhADqAB+o4t
HzxfeqSAftz35yTCZ6TPh79GM6Ua+OJlhtXnlQkVyqfeqbotXyDLJ5Ro5VNIZJ6GB3Y/9LdHOiZ6
8sQxuy9JPhDjed6mhHAEXFjOjM/Ir1dc908j42xVzIe1PXPZ516wjXHJTvHuEXPbxNI8aiXr9G6s
umvqCnIia0+2orKp10hQCfTUw2xKgka37q4VAX29tJT2GXQGu4ze+9vgGoWoy+6HYz6tOCKR9yek
voBIqEudzaaIyW2p8C11hMeWkbIUm1tofNN9GOIyktJ+L3BpUPB0dCl9NTF4UESn3LfcblO+6073
ksjPiCTUVYTx7r/i/ZzjE5UDfPB6oUo5Ygu4O/qvccVrL1P/zx75qwddpUYeTi5UzzJ0sKOqSxV2
0+O4YJGulqhK7k5ZiPR34z6KtF5+tUycPdCf9woRrm3XH+8F7y0nr2q7IcDysVBvtZhuVgDIzqJN
ycnuLk98OFPiFUx2HK7FyW6c3ugWOHWSSVmp1QiGqLFnGvX1ztAn5W2UZ1UgrIvDq5jwQs6ArhLM
17ndBbt5EOT9gHXxRi9Ir29DqxYYJ2KfC9MR4Chj5FT77C1Ys2gWHjGFf2Wc/inQHjRyQxlrSSYI
paMI/Fo9GwyKTV+IKanXjeHkMM6ds34QldpGpjjprfpf9AEgZVy1cwqczUel+3/u7ZTVFwSXq7O5
Kl5yfwj60UvuVMxFAR7o884+NUQKM/u+33PgQdNtb1UjTLK4qGg70qpNEk0kHIxc2tjHD9t7kp5P
HSkUgF/C25pg5PsRHnNAkLSrxRdvFYtKdMCbJ4Iqq7qyM0QjAXZr/mM2nqRKWFVINO4bhltxlkTq
OgcFb/HxS6818xIMlzAGOfNOXFDUKMlqAirWuWAUENu6NdobxutmJeIHELu7pj68qa5Bnzl8IngX
PA3OZqlfp3nwO8EqrEtXt6RfwoMaiXi7e967otLG3A7iX7DoCyxathM84pBYaicRyjgTpU28VBfQ
gIy6sskQloEel1f6qlu/+pwmSD/bvtoUVfBe5uH9NZE5LQPRccIyvD7fFQ4JpgEUIKUmpn7YQD1/
jtfXIJcvAHwF4MD6ctrMfdtyaXuno9yfSzsIdi0Agcpt8G4tqbDV5u8002+Rbqdxjl49/O+eVU6S
IR+Mcgu6q2vRc31u45eMts+Q1ssczAKNrE35CFhfKu5zekXn0yvtbo+qjSsdSw5Uq0BSbyuMMSsQ
vf2mgFuUU7z6cr8cw/iaQGBmGjbbyOjAR84hbdmB7mJB6JYZr/v9Qa1je8cawNzvZL6V7RuxvAho
iqz4jZTdWGKe0rpqgm1KZam7CDh6zQqM/IwHDLoGzTV3arHuRQFUGjmJkRCfv2wqMLZdfXAOBQEB
AiMJu/NISmOuZK2BcpK9kf39tzp4IS9MukNEnXDM7KFGWjYCqT58QJxDYV+7kv8CnXwvOUQGywNF
VqLZk/rl0WXU4IMjdD+8r2PsjSMZs8MMVhIQoWNIWUJ/3RST5QO1DHUxvJrQYJct2j/fB/wukfr4
dkhGWm72LEkQ0rICvaw9sROjCHOGTy5TbfCUAfe1CBNV8o2xPYky1naMnhs9Kk18ZONIhNsktzcC
H40RhZG8FpjA2oCir7obU0FWWsU5SrM4Wog0R4iUclLfPtzOkJeaVk8b7BKs5MAWjTgMKsHt/E8m
oNAgGZC5KqYvB1FU8KZ5Y2FXdFcc3/NfMg7VkTAQ60p64iS5sBrOhe01+7aV2pHxfRhn32ox1xR8
7IJds/qtZSxuisLBA7hdCmicCoTItBoh5RK6oOeLMIz9s1u4/uG96tREy/F0uoOmpkUn5CNwRirX
nNTQBBxNZcayDCM3I45gidteyWMY0MEG8IuXkdDrmUMlTZN7aSh326GZnh4sOGMWPrG8Tgz5M7my
endz4ALgRrl+wo/E743Q1OLfUh3qW9BrWMTZ0lLwnBP9OPVax20+pnJSLTjDXB0xj/SyL1eO8+wr
mLo7s5yBoqAsBjZK35mSOMNZoyfXxfZQ5YG6GYaWuEIPFONecsY/tFmW5iE46ZMVuPPdexBbvXuH
ppsbFo2jG4vAOVjO1wu8Hs0uEkKPsuub80+/GJl29vBC0UUE50Lnp4PHvoC0PmstNIR2EU/InpW3
/IBRfF2ylAFQP01kK6FuEUUroa6Y8AL0ohIk3wn9fwE4aIm1QAIN5phq9poFolsR7qkJFqtXE9rp
eReCtopAtgjb/PedFKO94mUp7+dfNOaOfjeB0Qgv/pjKOKjkvoJFFZuiziaCG6IfHaN/v3nzdIkt
cJSxDNqk+aWaGlCw8DB7W8/N7AAS7lLkGxNvKWe5b6Gve/ZBeb9pMBPFl0kT6kC04cus0KKDQlcY
7654cHYiCfReQif3wybqEZR/xc4jNUwGT65L8icUhMP65cQceOmkA/a54HgfHExsr8vlgUUaCf+H
Zt+3v1BGGEo76JSg4O5Rt9FztoFcIwlQL0pR640GcCZdQ+AZ55zv5rKEisxmrIuJwNSFNt8NXoqq
d1bMvMJdODqe1LAYU7cquncHcIP6kog1sEnrectxU+DDTN0jvo2CNUTSnMg2CqkHAFNMwgQGRDsg
OwMZQw8x+R7aFGkW4kiG8ByRXy3bu06nCubWmWHzKzZsfLrF7CPa9M19uojOBjpl91hfJ0xf89pr
Uu+WmZs44Fii3P7qi0zqAgV/W+I74xQmJzNK4yksx5GGEffX6PXYMJZex2PnIg1iwVw9tW0eqgAw
Rcd5c1/0bDAy8zIkQGk9fk6FUCW5KsS64MpSrGJ4tZLj9duWMBi3ODfxXbYEs+tWCAXAYh8V0W8f
CzSwemiqwK1cOCyegdhqM3Lk+J3GVWTsWgAP5t01qgOdVFEurJmUFQf436QPevNdkOzoU8n6aCB0
BgQTWcXU/9Z8koPq9Wbs+Ot0nShWmg6T6HeVhWYH6Y9+kIbm1aU0l8W9xinS0ElUZm/npTLFWDUU
ASXiLw04YPqY2tgZ3osBXD8J9pwI7nMgNbNOnxSRvc0JSA3rFsOoNrBKNj1Ra3zXmOBz4YFCuul2
CPI9np4/AFCAUFRfFIJHohW6uHXmjezoOvOM/n2V/SQRVFsl1plUAs2xNS5Jx3W8MM31ZlE/IyrN
J4s3SKl2bqL1SD0+09RpONlBE2kJh1+2pYGKI6VbZixXXpjC1JTi7eIUou6TYm53oUQWonL6t8/W
Bu+Ke9rLsNogAF4aM0YiLrxAt7h7iAiMGr9XGjRZwk75NBFsf61NnTWFwXT+vyyDaEAOIF+dkFs/
6geDK0zyZz/sc10Ll3pXjmXDpvqBftUCLSIrUfULbB7UYchcep7EXqY/TocWNbBQyMCkTYcPv/Vy
yUwKmn+EOZf/b3c8KMJj5x3oJNPqb5uuPoigy+21qgfPGW48Ihj43Qn0uAbrJoXIZGSnw4MJnnlk
61ebNRdaSBSoTAiZlrMUDpaOuedX+ED6078ItYRh/HdVXyg6bJ84mWZyXUiY0T/5r0c8NktFW+MV
QgBqRCtNeA16cEVs3totDYYnw+89BOg0nKhhJmZpvUVUSE3vfyTrhc8MydOpyYYhOQN7R5Rb4l7h
Q/YJZ54/jhqOm/zKtbXbnIuxCTpZDuIvs2IWvrndanoLKDAs/GjK7VQovQ+4GSvEaamlMV81HDJ5
d86SyzSSpnslwtejWy3GqF5BDkKdvgAh4wI/NV9Wiejs8J3QPA1quIo0a65AaaeGB8Eg4RQy3fSD
5ZWFwg4P9C/UVjyC3PxCztBCCk1UAnLk6kK62AN4xDvgkMdy/BtGL4Ri1WGoJttjjt6Ku2AQLz6G
pGHqwGVTU3nTNmKbP0NCbUVKB5GmhigDWpsVumKa0ar2IVhCNh/qc1WqAxUFk1m9kn3Evf0AO9PX
/oOJGcsTePjXjucz9QOMY19ZNKD4fZuX5jFdf+WcnsM8HOXjfEcdKM+cugo3Uem6xl/X9Bonp+5h
/YJ+KzboD9aQQPtOxlszTLn2UT/+XoLd4el07BcpQbPk24wB+MfLnUI2i4Ms59uc2L0moagW5NND
ZI12W4vLSd+pUcYpnI2RO0nTGUWmt2bNuBeDRcq5cafUxb8JZ4LsDy8Hjv+klu3+VTN6lt2BTCQ2
mwdbgoaqM1W1bhuU9WnpKyzKgMt7+FWyc+zR/vtvD8kb/zxKzQFauadHW6evmoQlHTGtV85wpzEf
fr0COqgM8kNUsL0+ZBnj8gBKTMYZ8MpYOiNSLhWilt7I3nGiOUMi8Vveeh0rVZEv+2ctOr79Caf9
Zc99y9IeE3XEuyBg2uvaHOg94EqCNsIaMU1+7LsAbIvkJOUhMPtjpaTkWEHVii8PG07MhZ2V7rqC
k7wT333JcLIdmZHtfnnPCI5ydla+0ZISSkIDmcVzRw8svEEc3TKbX/2UCXKtRr0Dy1515y9VQRcr
EjTMiKSpY7nM/sVW6hR1mBKu3geW15hx5fFZxSM3Q64V+tJrIAWFpW/Ddn4DEvwnDP6vU7833JD2
kvuDT2kAU+IwrnTU/9ApJMEiiAsYc/6CzYjGlB+sgQROwG0X7QWDcoT84SNuCW7/30DyBffE4Gqb
Ej8+osXoyk70OLC3tzuiY/pEg8A49MtDZ9ViyP0E1tv12F+sWTWY7VNgPKcwgczbE5Bhafj+xELL
j4ochvSumLMans+zcKnKOvFWmHf0+gEnlChKdkVCSlhSEYqxDB2JlwLSWLkuF4/n/bpNgh+dfU5K
gsHw8CeUtcIiimZP8nQWQ/VmvKX2plIPi3Z/52XwsVMG6d6EI9tlatAvyTRWm7Ne6sDzZlc/j0h+
gZ7XJrt3HNIi0ISe+u2Y6aqclR3OkpySBa6+TZmnhvPh+JtfhXjtfoiX9RbgjF+yLQritodmVnju
YzENIBBONQIeeyCjHNbSUp+K3wAtJ3+L1pvQOWYOwMUncNWwUQdto2CQ/vGMIjJUz4PVVI+XhS4b
OWIWVHFQzXqmRrRgUTaFMYxqcL3TE0Xm68ZPDdSGpmNXJ0kMLyQLELYFpc6kY2LmYuuGvNxmD5mf
18zR2//NEfxNY19RP2M58TYvNFqDWeYpJV7pMpjLErDBGMrJvczNCIQla21eBLNJ+daLApnf+w5S
VQt0WYVuey4T4BySZQMz0+F6UHeYJzUSzq1n4SXeH8i/HG0yotqBwezVOC1+rVGVYw6Kbv9aXM80
IrsgYAdIkTPMuEhNRiLacQ8tu3h2LcV+Pg3BkbtM+uFIxaCAOP4lUh0M8iUvbsXGUdbwHN2RY8nq
VZ0uYWrrXVhwwl81RNzpNhP45V/5w7TnfhgDpnYJMlA302scjScMZ6/VKcqdlKXlPuooBp1VKBo5
6M0/ouDZn2k1p/SxKAve4wJ7X8Spvpze2SO9TJOtGDrnHgD7sfOjmLGiUfPG6miqGzHmsKC/+qRk
TT5Gj80LkvmG7G5ZaVh2E1oMrwax8tFeKo9KRr2ef56lev2EaaZnXH++QtXe+/G22FFUrhkWIeFv
xFUX7h9cjGPSOD4Na7DIkWq3OviZu7z07pf3kd8Lsqfw0vG2ERLM9BrwA1TDFE/1g74RXVtKR4Uu
CKJlez5A2T4MTvo3DXWDHRfAFxdRqAYiWDySKiufE26eK6CpxuagxuA5YM6eQAsvWxj49Gw+4bAi
L5+XhWkUoI38gOcQRA841z8VXBFYsY2eMK36Bh8p6YNXLCzTuxX+C00q6lcN7u52d9KFi5adSHJB
sYWf8pznX8sifsw5zKnfpnvdMfOSjZOgUOZ6eGvoEhgEg8HSd9Z6u8X+zaS/ZfFRE6fhhraJ13ZO
VoAnYpJcfv40OlsQqK0cBdiv0hoowB/JNALRxpXsDmO2DDUz7je+eexX1loNh8Lw5Hx4f1OHLZko
UZ+12+vV+IytP0WiOAG1AQkhCUCd6Gw0HcObB1n53gnlEnbThKRP95esFmxBOoTEulQ5+ZNGqmf8
q8JRtrLSaQt4Y4jg77FUvsI7QE8OlqSaWRwsC4y2hzqBZLt0/ZaPs6WYX1wKIpjIcmEUIWqQKQtf
EvmIlz22WKFc6R2bz+5/M+SgsG4MaCLEYbw2gnUN0Aeh23o3a2utDhN5oz0NXAiGFjxMPeUSbom9
6zSADkhRL/P4a8Y/yse1KxWvTV+o7UruJ12nOayzOH4VfQOsF7sx67ZFmJotLPEF/tjzwc5ka3We
96KZ3zhYcTemO8BtpmPDoNys9tw9mkAwVe9UFuEFh7SwrT4Y7W3xmksXAdd7KeT8h3oMIjC6WN+r
8Y8oDsrCM843uZSLsulIcxBmJNgz8n5vMMIqzUF0SrNldUOxLL/T/xGwemMQKaZCpT+Im48Hz/DC
u+hH8d51fJ+lDcwLPmf5Hw37E0HiNpNgVN7+EW8w1vVp7VscDm6IMjwKqfTqNfCGG06hUCrhnrYy
HtHK2R62MSIuptuaCnXmAsflwjb4vpQ3fW8AXZy4iEGpk6anPRMduBsi9nfiz2rCObYB+4eoKsB1
w0L9ziq7Wodqazds/DiE92+FW3xyZT1Wj/wSd8WB5ECeJ8aSTPNff7nkEy3/FRi2IF3CJqd+P1Wf
ucuxuqG1YHmSbNOIFZxCywk9Xz6LV2+PyMNqgfqdO47sb1LwkW4tlokdT2e8bjFxxB1mK0HiSgzX
FU1eRTFCisMfERg2zFa8d87BpdtL1jjS1l/wTyVVOiVbbZq7+ebBFzZMe3NO/mwWK8MkaxboPNt9
A4qY1A66R/py/FtJllnj3Pr9CmfXnAeBPlHcEn387S9rOWc9FW9Uy+ZF93RIBnwD/mQVpectDXBH
W890icQl3CBcMaDYUfw8H5fJ1gJejeN6sZa9k9UYwG3YH+8uK0POcEYF/v3asNb9CPcfK6gdubxc
XgVnsvrJDzfHKzJn7vvjLfY2UEr1ghkkofGvMxKS8ARaMNo2d70kZUOeS+igb76kPStB6grtvvbR
LBtAoxACdf+N2JbK1KEI7VwhU6BjEYMtcdVlPXYc7GqNn0Ypt6jnvgz14ZmNl9wKIW81dlI80oA8
0iJW5Hhlqdvsj3QL9GpKOnAmT5674uREbOaS0FZtj+WGIQT8bo/26hiDabhBIyP+73VDBYevsnug
shPObUSHyjztLcgOy5uoZ486UPGSE7KSY6NRdICo/UKNO03PQZSfSflmkaBZCm2BXSLFFOVHLp4E
qbppR5z75zhe41qXMuMY7CaU5Ni1agrJb1NYMrUbK6ZiLA5esyBHAjRgiaBgg7OynZUOwu4eNcB5
0u/2insNBcYM8F1dyOl7WeAGvku2pSBByO/O8rhhjkBa2op29otPAHMtOniAhu4wCKyrkPNHKnyA
QnJD8HtGI2QA4z3Ojzgc7sAA7cqYpi4lJL3uGNJSYgXeH0v7gqgOpWl9V6dFWpjh1GqtiEQgrBMz
wh+W+MZfWh5NItfVGe8e90SBhk4o7WfWVrQmhZHJlzxzdrZmH0p1tLIQQ6oDrkmZlChq+dIaLuWy
FJk1YvpYhrf4j6AIdEz4MWNLIxDfjeWg/U/B7KMhb+XBqBFYmXRbmNmdFWDXSvBdpXItGR7Qq192
PrbXh5gFrkdbz5C5DRrM8eEsy1hNrtLf25kLAGQyNUe1aGlRDW25rKWNItie6JFSy68hS6GhlCTS
59KhB0REFMz8dkjwSYni4vvrZCIl2eWoJ1loHBNxgTJJtjRSOBKb1/9jtKRIqzjCQGfBXYs7wT+O
S8ItuW7mDEOBcAJZ4mdEAqN13L5tCN+0M1RwoZSd0t0U7RqL+se+1Zs6sxFwbNtcfzwqZbKXDY2i
EWvvTpSlHE1S1T7adN6/cEZ/0mP9hz9rC/3r/kl+z0HZ5Dt9MYK9OLEgR+nKaqv+03nr/iMKVrF1
cmTNkFo6Jd3b6A0x7BbVo1RlGPXCqOY8B2kC7PyHoSSQd+dSR0Tnw+EzNw+4RPk0x2AzTjiKO4qP
F5agyJGB7SSbMdB0og1mMxUNqgbujUrleOAB8SZyfqFxxXB3e4fITHp/lq+Lz+fr10zfEB5BEkpr
Rfy4yE7POW8lU0Aoi8HvwDzYVFG+ifGycQbpXjtC9MNek/ArUrGh2bkTMWf+1NKFCJrWdHGii4Jl
o6V8AwPP1uUjtbxXxKShnCMuh3jhph+58Tyd0xnLvLEucyFgOCE7sBM4FIltVa/HnpxkJMuubupn
U9lBP++JuzqUIJbS6oI9BMnxcUzsJo1lGW63ksUrZj3WM/ll1LFf//k+ib6tmg6o+Jk6LDEpzYM4
RVC8V9z2XysJ/tyvenpIl7PM/Q+TCB25YA2OVb80xEmKQH0LXhciXHCBL6shFRdf05814ibpUoDQ
8StXO7nXyTvrNSZgoss5yCwMLdsasDDFC839Tr8JZ900y3mbyI9Q+GQH78dcWG5AdZ7dpO5MSIAI
YYGKdaTJ9Mc38W9sGb2SVYdq3m8FeUplyzDfAvZRi0NYvUAlG7L0kYjRES+XWKxD805ps2W7F2nH
2wSDmZA5zpCNvu5YNjzNbSZ0XBayakaPHflTjM3fC1pEAplEH7hMe4bMyF7q74QAJyE4yVW9SQGN
jCqWHv9cgzL2qC9Ism+gpJbtXXLmIBX96RW2UHTS5IIa5YtL+koa/Kv0jspogLZ+Fj/KsY/7KyKF
NR58EdgqOrc2AR9Lu6VnzoGuMODSW5Rk622uPcdcd9yD0fsHCsb/h3l7ul2fCMaXjavXm2yTDbBI
6dreYd/7u2xa6PiUk7iijiSgKYLLowOAPhHH03XDqVMS+XC7rBKGWyQaJBOx90DhSC51ZqeCH8QM
CWVdiOS8olOfFAFIiLNXSiO2OoxvFJFTp+jh7xLbaKFJz8vOezwY3GN8Y7o8HF6Pi+LxC1v8oiX+
CX5lrjI9uxqBFtVmg4QHFhiDKfuLojLck/bSkZuFyiVi/i6zkLUevmQBIcIgl1nJFGOtFsQEu3cq
+p2gSBxQWMNTMbY1YcWMDz6vaSPV5GG+fwx6UU38VCDJPVcWCELNn3jcoYppCxkEHvHdVKlKGBUa
fyuEXuNKk87/Xh63WW2JLuOW7Ovj0tSlIkqHR0dzXZ/bWFVUTym7gmlk5FAUp7Wqj1VRQiJlRQnu
Dqy6womkp9NULMwiPikuehAOjTCszktKl+tVZwUwXgFd6rfQpxmPER/GmFPG/qJnl9NjE8yMoBnc
31fofmZZOQNwW6MkguquxgCssWwR5VEZSoqyhOXLs2fYIYf8itiZ9waA7pDBdht501fUluGRavl5
ZH/0Ui1Crbi+sIzPVRAblxxJwVQkkKiTEXJT8Wv0tkYf9mqUXWdr8yoHKMIosqSO0ebSNXNQ3fcv
/o9n0w9Y93iBCpKr/7t1hodGesb11L0MGyv9vjFhMhBiYztv1HqSN1rY23KOPTeQpZQXKsT9CID3
ioOwy5R0QPESPwnFISlKa1Z3PZmctCWUnF3vGxO+xY0HpyPUbK3LHUMKQUL09j2clohEfjHsDsoD
/XcQvRasw+RsMVp5fF57zCtPk/22ZuHDUQr/oEtlqPxQSsqjO4wAh1+UcHsRKVXvGlAVpHhOqfW3
CxB2U3cXcMen7IOLF9+hT13lxpGoFdxWfEMMsJITUppO7A/Rsyi+5Z0llMhsFYo1tklc6UYnO20O
GkpazgBT0RKSceU35cob2pPEFw1dBHHfEHPuUlJXiW38JkX3qTxYZf7FAu9/ezvZvyrCLA3B/f6/
hrcnj0rhOVgtIctfAv7N8lL3cwRlZM7DDaFK60JFORbTuYjvBVraM4YWyiUltB8oT7RQ2JQYiLv/
x81SBTHiupHqRoaG5L8GxJLFjUq/dZnYhRZ1exw9/GYKHh0Fj1nTMM9mFwqoEWUHRfvGr9Z6eGHQ
Kq/Yf0akjf27LrCldsQbBAnTxDd4lOuYrdR9nGo7Q6VLHpWLrKlvmXLxGIFKfD0/vle0e4/Ce0+z
LfT+yFgw18C1ljFhnKlrvD2yvqLpkfTOb2HPEwAhmmUMETvlQQxAMD7NQjZWdI/K9MMELKRXCMAb
Ld5uvl/4TYlfv4OJ7D7+zRITnETYFG6WPl+AQkCezWBLgGZkHcntIeCvXRz/1U+QTjhKbOJ3Btfm
EsXB/tQQKZKogYIY3UFPNVonzr98FPQjfIeQwMbgbH0O59CfSf8/ShuKHSKaBGerLNuwsAPBBuwh
rFljeSgJflm4iNqL7Ug9c2ejIhUUEjUqPmMiUCxVwm/LexQeGSiY59WoQaZu01T/ETKcLNjW67hE
yZy8SmMDkYlWOmroee4/KYmP2on9dsG6UmYm+G16lqyCABctnVaqUooYWZ8pf9onJbwEQ/OwOcAG
t1j3hSnGt5V3b2T3KZv/wVh6k5tm9SST8dEmfo4N90l+pdixvzVLSM++pHTxNjohK+oiPJCBWzP4
1axstNj4RBF/yMh1oY2rrNE+S2VRCfGcPxxJHnsV9ChPzaeuRGumBgfxmxvUoETf+n3Y9L/EU32Y
nlcbcwsvdfxuIPUDj1waZBUDP9WjtSWTvjQUNCQ9Yb7WN2Y92DlhSI9e4+95CRg1FGhLvvzoxx1l
5sHphtFhThfmnjwmXUdkP4HNgXgSbhp/ATYBvh6yMp9HWyNa91mXeRCtXUoxc9n6HUe+epKntrn/
ap1+1JZ9lGC5ThmImCpxC2H1ceVGQE5+hF9zpSmDwodTecOLsFgpbso0vxJBRCelwMpYZ0G3z4yi
U9oiv+VjQBZqItxQCE2/PW11ryE+fCUzvms22XNkmQkVY1xlsB0B5Qpfj+XOYCM6PKaBcFqqnFJN
xJatl2ZX0AX/1hZRJOMAxf+R53LjdWcsA1oOMb7/RphyECeeZWkuNjRYr9yWEacei1pvvJRU8H6S
5BGkZAvT3leDAuX3X7yOBm73kjYX21Cu4RQZOeVUFpMNTVqRVxDvOmX5nyuPkE2Vm9nY1eCNA4EC
k+Yt1m4klkhB/XkeJ0mLBdap8JKbgisYf8q0dmwT1daK9yYzHZfYLbluHYusbocjmKkcoNERkdLk
WsO6YZ5f3cAxG1QVWjHXj1Gv+H2rlI2keU1OhZTkQacoAihsKeA893pehKkCYSvJQMoM8voBmGot
0lkeplNejKVCxkhrd0nBpvH8HkuSYA8/BCIpsB+5Mkdin9uuj5OqEoEPYFczt7JlfQ2Yhq6yM54n
EGTN7OgycVBpGvEiQ9XJxm0LmLdroTAElBO+5Md1WNcVttcr4poSj6ubkVmr82EQ8suYgJlNJuuI
kvcHx6ZW02BRn+c4qt25YTLE+NX4E8lkw0FlkKnubrPKKAWyJVwiEx+zxZzXrZZGCUALffDk9yhn
CeQvZiUEcY8DGAcl8sRC7RuojB7GYojq6qgSeKaEwQGZt6S4cAWZWqYpu9dJb6m3VXgbc/QqC7wu
ryMIvLa5TsQrDAAJxYbPm2Ap9HGLgXnhFmZaPwdvWYH8SlayT2puw11ddvfEJJtNxHIGMcVbuQ5L
l0TTa5zQTc7Zpfml2NHtUr4a/YWY2Wfki5AeT25RKGKe5GmPikZh+xU2lvHR3pvLUobTSJwH4JB5
LfLO1glGQyHQUxkvtS4Zt9cuvVA33l+0H23yJvK5rKMFUF+XCibcKDHU00uErh1jkcZXvJAV3DrO
ibdUNzMP/84MKK7i9Y0hVAboRKK5ft/nPHZ5VKG6mC9ZoDPJZrvUoUXaSu8s1iddmtfp6qBvRgjI
kHWR3F2X4yCAZ+YrfaXApsmbKUHvUXz7F6Pqw6DkW3jIamYwh75RthMkIvY7W7RfOksNchl4HEY3
5DaC42f6Do/bY7foCBptHn8vs87TtcSxQbL549ZwWinvz1mY6Z2eweJ6Zwoo2InIDizU3VELWH/h
hJwjaxCSJvMFvGgjHXKmW76RmEK7D19suQ3X68Q+Tbui1vcEYNKEq9rdx37qyHp2W8dM3d2KHR8k
yq4YpTtuL6w33eUt+7L3KbF5k/SuD38hswLtQxgKfQdz+gtiMlMrVB39O1I46Dc7gR0aURjIQOTO
NIn+menBAKVGhsKRv/D4Cmv54NJKRMhVVbqWs7/THZnFeweuoBqpHxd7Xd4xIHA5vgzMZkg6ydjU
Mqmd5JQONCBqbVoU3UjSn27eZ7W11Kq21ezyU+aJ0EQTemJWVdVIgkPmhtzHKhqXY/fGzcOnCVuW
IvqOZFpuf8x5wsW1o92cY7nle3fMsy4iNlKbWrc2ZLbFiHLYRKkethiEAkA4QaGcdNa6Z04/RGTz
YHl6J7RZqvErJYR3ArA0uxEoKzRuX5ibCBPyB2YK3r1v3hZtrsvjGXquRRGL/R5LKdmByUpYB772
9hMfInht9LR6A63Ru9qDWxUARHGTkRvtyhLL7NctNIVePuvLeOLkM6PgDv6v4jjNZx8jVpEUM0q6
QHYWxR+CKfzrdFAuZdyIS71Pu+4swz0IKMPbA4gsb94vm3eSuPXwxhViVDw22GeOGRmajkXnJHpl
8WMPwQAkBolIGzLsmV2d5Z1ng9ARn4kRbheHfvKSRnLtGkKCrCrOUADY+OTPMrrTa92FDbaNinti
AVF9Pg+limxxoBfp9e34qgIn33FQBtme/u0l0gftwv7MVgKzyFLoE5eer+7dXcGjKbyxTm7cU+Kq
FBqMpMeMU722tJ/fWmrpun/r2jfd57Mt7gWmdppV5xvdUcicroOvgqOXPqbKxkxVqJZSI0yhyTzY
pTbCU0hQzmJZVx7ZpqEEmf9DnzrSWukcvadnow2jZmeWOICV1yo5C9sZPwe34oan+GspKqwjT/Ze
cw+98LigWVeVBkCNZZN170xRFCX/pSSqzwpIN0tU6prbAQ5aPpcOXWSgNiXds34MDzW7nkG8+7SY
Q6SNfmggz5Rzfn2krCDBiczNxFTAevKk2e+PRz2Y5+oBqfj3xJrWNz/EaROext5xqEYZaxGJbhb5
jtI62XU4DxjYTQeZ/joLxF+d8OaCgvJsq1jEQPB8ia5xFdNfRb8vIa8/kwMnroIRQGG3yJFkCcz7
VAbPf/FAYxA9p0fRsMION8K6E+7eQVLitjlctqHbUs2sdF+HF8gjtfmbE8/nM7PlqAbdxfA2aa6k
+GX9QwzQV760T1KZQ1aJ+NPoNxfvzzi6mRtDYqOM5pDU76AoCSwtzrBMh5WSU7bz9UjxJQ3L3inc
jO3ZKlfcRcEEYdE9ZYFx1d+E4eaeTd9R6QDFKgmvZt++RiR8hjqhhbAWWyZJ6VhA+Ypc0wOKODE7
wuljb6Zh3h4RoU4o+m626k8Lo9sovh6ow8vcgBoRKv2nh1ZR72LVh3CEJf7rH+GheOUx+pgLgpmm
oaDhinhF28pEfhkFrn3UYWXX6X4/g+LsHkN9pghU2BaKw0UZwZMF7AV6qMoSosOKjJC3J5YzBMz2
rNpGdWTK0EvREdiidOltD4vugQUxLLDnhr6wwXtQ38f/XIYbQUIr0Eo9qlBLmRfOeWS8Ep3dAhkx
JbsT9rT2BalQdXJFYybadoibpj753LbOKFfZpx+J8Xzn1gn5VPL+qDWHq2X/6BBfeTUxxOgwjAf3
drkCniQthj8ScS4s2ZUKFl9PVP9+OEdrRXBSf3HcmTIA/oNVCdN9ikauJYwDTF8e4+Eti/cnz9Qa
LciUWv/VhO5auQCaBYY8XUlwBJP14eAeac8oAIvsEFTpPh7S90MTtxhDom9jQPwqWbGYvgZgO6Mj
jU60jUefNl27UpkkTJGZWP0l16zS+le0czLjecKGmiR5zlxS/MUBNF2Ub3eITKkMqgtjn7McJ/Jr
r5KiJrR4iQtk69BbeHasRLL4IhdprVRYcNjhIaP5kTVBKRgIHb85rQP+f8pfqMlc8+T/ghKkrTAP
fPxShES8Xo+wEnIDU2lFuaooh8GUIjyu1BnowiVTMFhtdic/Zr5wd/1QCLZJ9EJwi1WGP3hvmWTx
1UsCuGidWSxJxGt4SEZpHx7tpzhalyCMFtETz1g6LbKUP+u/6mkkaJqVUtmIKlxvJq6DOgCIiqEW
55qGVDQojlo68EId1mnlngPgbgPPebU2AJZnk8T5HlvnTdIGV7rTAXxWO81wio9dLsTr3/Td1nWN
M8juANp68EtlwHFgwuqWAFFh8enY8JhhfsRyj+VvPn91fvZglw+wUf72pe+L9AOdfv2Ynzm57aew
LvE/ndGS3MMaR8wNbHw3tn8RjyjBhswUSryVjYqewAwRBIGPD7l2Wqk+QeBAgTdgLPmybBVZ4oyk
MaHHcaOg1BlcMDCkrXQvRnHRaEqzISyPTR7YgCf7be1TFmc0I0XVeJGhew55XWC6SJtixjmwaaqq
50ZkN+OVPKDKX2r+u/sctG9Za0nbv3ljyItB9edoIxcVOC4K87vmZOVfXagzAZunLyGnES/RY2fD
SgZNjLp2UR69SyO3cp8BAsj7xKb2aKBxJDuykU6NDTcpWQb2pQm1tMxJ+iIJLhFHc0Ax84mqaCcS
YuVug+IrxBVangI/foVKmQ3FsttU4dFGFGzepqJic1KOkY0wxFznXkLyeydnMbxBoNb/HASyVP9k
zSqzw6pqGNdoNhA/Y7W8hsbuDax5DcAD2I8VHyjpREIyL3hrChdvSMya22Y2DP5l/ez/67dM++gP
xTfhqqyjcYwS+0uKSLSKhG0p8kfIO5ijlYHDC2fUvWSNTD2PDdVVSy9LH6BrqUaFJEmTisdCcsGh
kjs4aHEJkNqmYIdEx8+hFUccD20ZOzKhkBKkFuo17xDSGoa0iHLDSo9M8Y+9Rpu7D/k3viPaQ+cr
4razkXTZGasLUsXZooatIgM4vBK/ILI1bnDdkGTMlIpZXf6niCvXcOxhsGmd6HWdjfRyAH8VCihr
U7U1ahuZZRS3prFkoTXrIDB3j8FjUOcAS6NkUlJowAJl6IUZP77of79bpMru6732oX2bxLUX1Mwj
5ml7zMk1k2Q2EjC1zBzFi6lFRwMtxUmjx/jT3C7vXhD/6f7ujCMliuXjTCkoqjo20NBLG07ax/l4
OmN1geMAMNwwCDMt8vsB3MzDnhKbmuDysvdTVoj+vqd6j5qVot1Wm6PS3tZwuqI1wzMJ7irF4sDQ
g7PVcahgk9+A/GYbzLCAfAfV8EDeSCxf+CSgZnYMTvEhGNsAxnOH2jXKlVv5QecltVvNc6GVj4Uh
a4iLt4hfAiI5ZBW25ZWXFz6pYjsJZ/pl21j4F1u0tUjD2j+48p15hsYXWe3glYlBXW7gCfXRrx6w
fPqQF2ZAdyg9108ST9f7MjwuRV/cGVssMt+0KwwvQ3boBFHV2KnTpB0o+N7PPOqe9fynnhGKjjo0
Ia2daccg/lct8t7e17HZpOtX+4zieTGA0DufLwjIDWFO4EGCQaCsD6HnuOMPPcUBSRVdpASvkvaC
sVbPfLjkXIM2d52YV/O2Y/v+X5942CHhRPV/eJtMtOzN2qBNdeHy0KeMJx+5ZDOKFgL7r5DrIj6X
sNBSsVvcn7LpUm+LQOeQObsIEzAhxFwTY34HyPoTijEg0O5zAhcnGx38/Ii0pa7GVQg6S6t3zDJw
e4UJKJAPI382XN1F+QsX4JdtbQhyxNDK2jEP18RlV16oNQvgy/6a0RgVa6FRLUVOVPsDF5bVBPBu
1/54y/9hw783ce45bXQwq+YxmG00hu9ppV8eJXPfEyocVkCJ6auwiLZImNXO0NyTbp4mxEGoCJW6
v6gccc7aGK0mHykuBEjd/f6Jei2Z6MlF/yn8fCQsOmV4duW/KCr3OrNkWT1tIFJabxbHovDGQh8p
BjmHkm6Z/Z5Al71DL+ygjJkKALk2C4g11jKTHmbYALQSZaXt9frkw7I7gps1Bew7WYZpXoCeIhfe
FUx4JlxAit3mSwIrff/8Du0Ep4KP8KFcmH/aHUrGLjrUlcg1x3hj8yFYRTuOY0Erf0DCkLkvyLKe
DAxGimCOfGsPPTCEiDXPWG0zDbZWMPYrk9bu+2KxWwk5Mr7kDalEQ+cAsGmmrq5lDfVl5AV8at73
5xxo0Yr8Sq5AuDt+m59bUz3Tk75dh7Yi05uRUM8T5JCAXwjJivHqGoaf/bA3K+mhKb0Qrr3jMJer
UAKGDaSMLHzWEsCAE4de8TbA32Yh7Dncg4s6ufvkAUEJ4G4GetL2v+nHSxwkuZB+XhW5uDVlelFa
6zBp8I6yjBqQvAddjpQIYyhLWWWeR7wG3wQakkpyGVNcomy/WEew+RuSp8WihKK+Rj5Y7BUGs18T
nLqAFrY2aoeEYkyBm+FMQn8xOBKihL62aENKENuKggOi44OzqJnA8JE+ls/dsQLLKoPpRVfqgRPQ
+UcC/NgTGRXE5mh2McOOqTr0Q5a9BnGiI/bsUagVA+D1MuRwaXDUNxZU6lZMd/brsShpKEd5YIHH
109yWK4U03NkiV2Jf5d31Gqap7q32X+k93jY8Ne9jgc9Ze5og50w43A8F5SZf9MM2mpGvuZQwsuX
1+oDag0Ir8LF1CNpbUNaJN61QcKxp0/OLQeklhsAENjtJuBXhzY+85BoP2ZfqqlW6Qgn1gay/6vh
OZwvSItjR+d7lrN1jTh86Likaj2Ddo9W0FKl8XKz0HBIH0+dK8Y1QNs5kUHWypHjUUf8cNK2jvBu
4b0wUPXafju8l/k66CB1yUm+qUUNZ7hoz3o9SQbvbx4jtTkfhVsETyrEd3x0jowQvL/c1hO8QDWX
RUaIgNQpRCo+/IHNFzclrFCJaQctwy/jnTP3xopw4jdeXasp4Tozs+ZLT9hqGDEQqyyxpYNbTbY+
mJYY/L07O6MmdlrPYX83ICc2SkTS+lF+hhzNwbrjDIMogWdgM1JwVv37KIoyLqq1rHY0sr+cx1GC
P+c5E4fVohAicnoPbb6vkQ1eSm1Z8R30e39hsyuRXzn07d0XszBUDgGX43ubT8MRro20+0p73Wcy
5zkNyptsjNrIRV2/mQsQT6PV9E1M15gKBYKhRM67WtgUoc47CmrQCng53EjoKEDhdUC04QItPkbm
QfI3z5karadw39nHSQb4p2UQleuiL6+o/yYQftJB6efIhIYzDxemEtJIcraREilnkzgTH/6wnb5k
oIIb8ryEBMeQ9Euv49hH/TNtVleKMixqO7QJ5sYLTMY7rnpyMdLkOWK5tGW3WaMAqS1frDprU26z
bwNUlmYnOXM/P1dRiZ8x0SqtJbvi73jfVgc/W9R7OAD9n4ZwCzWba2mEPgTB2VSbhuzeLlcBp1h3
uQNNAq6U4tULe4qQWzsKdgIyGk/THjUGi74Zm/cYArA+p0odVctVJP45CMP+agf/fEk7XRP22GUG
RcQ2t+VFupaLpcb1mLR/V2acPgEEWuYhrbmrHVd+G8BIuOjeux10bOfL8Bo1KDFdS9XTXWCx0oLy
dunIn+q2wgW7Bro9NwpJbFBfUqyomz6VJbt/xFE5b3bn2Scd8PWJi0yrQR2pyQtpNvPpKsmhzshS
mdE53LRpkjqxw9MP1XpTSWHkZswEd7P6jQL73wzyo6WdJcwxKumtBof8D8SbM1WmfPxi9afGM2Jk
VO6pXImg8p3qiSbYhOB2hUhRKzeQgF/0M0Y9DDgVK9a1wpE3qZ7vCvoMRmWEu4wcEki9kJkb66xc
VKkD8p5M4LbXUtVCOuR2jOgbAvb6frSBG7BeuE/AlGzAvPod169vwakXUBQDTXFDf1Kkj+kdQ0jN
h0jan6CDupDNMEpb/4H7M2L1kSzLhl9REJmsRRtRvOvaB1hYoRV+N3R2GIYE42AfyX1/Pu+vlASG
DXQrduRZwtwDASw1WBdnjvovAvKk9umOUBdFd/aLnzc9cqmqtw+y5nZuXtifL/OaSpi22upClWdy
SP1BgGfkyY7ccfOX8iy0fweOCVFSIFqEkCMD0XPb1N7kSuQ5uFtms5zTTznG/nTzuelEu1xcVuNN
lp9XDsvC/rAeWXfkgUP7nzeVH3Pq9sfvnN8bZkYu7Gwb094Mkp1yarVeKL3o0g1PR1tY0qBI8SEY
P4Yp7fXOttRL5HZO+JHcC3jM0sDjBuXN1X5qsRTxoLhLzhjIrce27GyD5nrJeQa/4qHaf8OhUjJY
4ubsgg0MSxa/xHZqHysapajAPPkE/4WpmqGSC5h4AzJiTP0TP9JVmjVE3V4iQgHmpLFMNQzLeJG1
VsstfuGCbNGuK4VpZ/NumqhYqQH23SDYb59sVIfkjasrY9wLBrkrW2Ny9WxwT4ApRQoO1r09T0v/
vuRE8Cpmmh0nhTy7OPWgW1BlFo50g4m0FDD4LuxTFiNjUi+frNAcmQxgDZDjfWmrq8UumNlLvuOc
9VwAsLo3v0XA9JpM6QPKHXS0edDQeYvDJu7JQww1K1AfHOvQXag6QmK6cK4txKNxmxHJSB8wl+vJ
dAgCkSy04whfylT9949WfZ18QufOMMNwTv07KH5wmi+cSuTXXgLq1/WZxFs+x2VdRPhGVJc7YFZ3
TIZ7kv5N12ot0/RNHj81E4hRnD+HZJSQ0y5iFIvQLvONP8Jff1e+CACzGqn4oj6I+uJuONbT99f0
i9GUuTOB3nvol5HqcSGl6Y3Xy4Y2xvzEETJ2sE8+SeIIuy4BjuKg+Xg1vpnjW9l4JsUYk70AfIYX
C1E4wk/ZKrmqTaHPIVvY33yuuh/wJFkxvoACUvU3UeXLzZ+4p/P+p99xSK1dNHb/dUW8wt7XCdCW
D5UcsOnl1FBNFIZDcskPbCGdvaUiQ0NRnL53h0DK/hplKCLYJQ1Kcd3HHMnlU4GX1BFSkde4kS7N
32LzVgmLqXu/NtRBXi2/dMpD1XKjWFhOqf/chXoC0hpmkL8CREyrtEOh7VrmA+yFH7IMcoLpGt/4
qO8x/+Rvuvw/8wgxEh//WIxKSz4kH2cZsww+65cdqoEzMoEUBIWn48gZJ53xDlghX9uMiZ8ohJke
gpqKnKTw1+EMFIPmNXbMbAUPLh3/NBjOjL5vcEOwrwx+6cP0zHneqT0hBQMtzpwEAEHH/zGWppAT
zU3ARGPPw6MP+A1p3Vb0YzhrKViI88UsWFW2LxF8QQ9Ti9TQ0ZxOt6mQO6myenoF9eXyrscW7gwq
p20SfgyskM5dELuIBy+wpOMg8+4nRbamJgkIFLB0EaLIZno+q8mjhP8VXMkORRZbxTperHEHQ8wH
JLhQDf3tRwc54tjUBZGixEWwstdJtFu8at8C1Pl4Oe4m+40tpfSG/JMueKynMTacrDMxTzN1RnaM
SS+mUVb5VoWV2ycS5vRsSnJ+x8gvjZqJAAXwDyT4TBQgBaXTw/ujYyfwZzfk6DmXdhbCMqyUtob9
3MpqHJAvPehJD7JJbji8s9/NNZprtXowJJQdM7gU8S4/3UCYmhflXOoDMVRmBJIKI7M1T1bJ/INa
Kj1bGOL9c1MQBsL91stCbAy3KUpq57bAbnFu4UKTxlyLzeFu/4NUR3uVgqqplRe/MnO7+87WfV1V
hpbB/5P6Up7xIdyKs9TbMzqryYBBrBEjJpnHj31PvZy/fr4/Hm0cHEEWR7qHnsasmg4Ta9pMBZzd
q0T1lE8ko8qn8INPIfzL6DNxa0qSL7UwCl+AvackaAzJMKCvr6bhRWHRFK+LDCUw2265+ZS8saMY
K6VQ9RgFmx3IZvnloWSXVb7WlzkbQfgV8CNAygH2h60awaOaj4ZswX9Y6k10RwMyliwKWF+rla8h
SHZn3HxOIR+zI6AGKr0bylkeVIBGnrcjCKYw7+Pfc2je8Y3GhrLwZTSIE+0pUMP0d+Ip4MIu+zI7
fa0aou7K4+dPhqi/l3/dqFEydbuqQeRL+UVfqCr8N7MJG8FeD3mMy02pdea4++59wI93FPdk5gzF
WGna8nXkJu7UqRU0uYdmiqc9h8/Y28AhXNxchlvinTT83PKeSGcfUha0TeZLpAc/1uB9anvkQzcy
Y4DQ4CYsFGsB38eWttMWR0G1vbx+3kNZsGo0DWzIxDRkdltF8rMNN0p/GWAYKj8VBLFhWhXrRp+C
YLyfX9uqwWWiulU/gxTIMkmMzR/q78uUttw6pI+v2n8126qC1RTrJ9e0PKNZzVAtsigoIl6VUPq7
RduQHpsA/AKaVn7ME6Ieak/hJR0/ckjh3vHHUyjEUH2+wlX3aNOy6k2rgBO46Cx+NPDmIZC3GfA1
IXJ8bqh9d2R00sleOw9t0rpjBa5s9mkbIqm+s2UeAnJQiLcgXWm9vT6iE9ESxbpfm/JdDewJmHcX
tw6GV5qmSXtXB8OWhofU5Rnjtd/9iMQkM9Jbae2iPNi5lELG6zZK/pm1bL+3qCXDgjcJ05YtEExY
FUllh1FYDl3FqI5zFKSVaGpbV5HFYS0jFjqub478Nag8+V/Gv12T7NfDalDYUlyZIqQRJgpAMcet
nj1ArKmmD5HdqRKf/iMR/xjB8V4as6uxEWd0KJ8jXPYwgq3rbA0UCI5iCC9bFXWeQVsFfyQ7dna2
uDjpEVvVa4B2e9FzQOYH3QxKve0GM6Gri5pCbZ2A8RKWhAG7d0MSpvQJh736PIJ40HhrZLEsrV56
BMy6btG/+Pjm4Ff/okTl2Y9TVzrJ+mZp2PHmZf3jvxYMNEvGx/4i2oDErRKHSBHALmw0tEPSizBB
rhsYSmcG2z8v/+5XqLJjNHaqRPnK/iGZrNg7Pk6csrNJSaK6c2pKpeeJVF85zNLHCIw/ctGtFpEQ
4oel/zRdAKoNo6QPEKffxctPSHc6Vz9ZisY4VmX8DEsUpJjoTjN26Gu5pp8ur5g+FuseOZ7vittQ
qUFu+I8JWaSjUvWT1ru6yD+thFoo4dWRqVIOG5AvTWwF/wCnH5EaT6Rc7DUABoHsXIyBbYXma744
iI2BZZRif2Q6oIb3MTnfpuHUyk2fL+4MdP0AXePZwpF6EdAfcvrNFwrqVuccbmzUqBW6DRa1qqTY
mvuyJaIzVno1rj4Q/lKOWNNE4JpDtiiEMupjwKvJaEjiKQqh0K8KuKW73KcABjxf+dCUi02icB9Z
EodspKFfPLS+zbjeHWMiE8rohH24/lkfNVIlvec/JAbwsCxhSN7in27MTTiSYI4IDkxaBlCQr9s2
8EtuNABQy1zePWJpxX+kT2R/19myoa38rXNgk9P3TCnggn9FxN1aCsPku9M3abm5h5+QdifZlKwL
sv/bD56Tc6XKOW//ltubO5x88h3BuZI6r2O8iE+LYOhXlHw/5YFCiclDFAxdBXB484cFu0/ucRDX
4HeYQPTmuz9j6Oku7ZD3RCzzYJGM350aFsKr8J5Zuc1np1a/eTC8uBKctZMp6TQCicReTMYxQMu/
E/4fphfHiOfZIoHuCmpW4/lwLbGYJyIU5X5BiLEJECKWs8FpxyXKrhX3HmC/ph4SvqVGbOwy8enA
7yHdrrzjSchsW7golDqyTf5jWdNe6bgwDRfRVbbHOQIEElccVZEK8HDdv7b1t5ZESbRo8plvATyW
qHuhNx5IeUFW44/AbbVwkI9uDyvqkQH+oCR5bFwjvhh4Cbl9kwGu50USYCkdX8EEuCLOVTE4zEBH
eU+CbLS8JbTqCwQ0ncF3qrP5EVpi+pVSNR3Q3jcsGA2ALyq036FzrLFLLLizrM1pELyNNJc/L5Ld
QB1O4Q+mU3PmO1Lf6aBMrMqv6O/7dscc3WXUhpQb0SU6Qray/oTqKzDOnHGwVRO0I2zpBVMQYezb
AVBvyZKJ7SSPbhX7zTXDBo0XrkwJxUZAzYZ5pB387bQFgdcuhhRLQlNu8WfYILLTfExyuLznWnaZ
TTUO6+4gUy0IrvTnjWXwZOZBhJ1+R4jlUwipthhdBEwFguFaeF4JRszYkiNujUlChl4psl7Kbw5L
e9EuwVteYXAzQS3jVAubIDboOq9jqknP8pO9mth6X6Cc83zWjimXS/+Ot3bxaN5IHtX/TczVvkfN
VUALdtAdHYDki02teWA7ivFrLMPz6dzOiO3+pq275Yf5e1CEYTfVr/k2/UbQzcNSNDdm3VJ8Cq3j
kVfhch9WBM50VzgeuId6MNX7/JMobVhygXMKs2VS1FH+sYcp/Uo/JVpy6iEf06biwFb4dUYMJmV0
12X2z6HfB/7YjNb7dF3qR8bXKc5CQZtrwCNUVIYgIFooTCxDZ1nGJH9EObFdfbpZwLFtxfD/T+4h
wG/oDso2UrAAr1gCflBEcGx5NRfIA00Z8K1rg7c+TOqMspeSZOj711dtD3re//9Yh/amHtxfyRYu
nOx3wsQ6ABBshErH0FnhCW4AtBWG9nDvqv6w8dKZwIIFyCbJXvjuOaostJ7+ydc6Ts6jZ93S+n9e
gCnjFiLDamoaGODqPoucSr1UnYHOKiRovuo4hXEPYnqA1BO62dx7cuk+OcsaV0hDLzDgspuwDBPZ
n6XoHQovVYj/dM/fyMEl5xbBptw4tu7/iz0NuPHpzYorOm7XkYVNh8TbtWPDbvDMaLEZGDOu99wp
nSEvdFHQNDjhObrqTopft3roPFko9IwoEUMHFIdY6bml0nDTlaOzatdqWO1/LNs7RM4l8xe6+JQ4
hKQriVDryqKRhv8yrhdKRr9zTeW1tVHFsUL1SAaEbUXlk2385UDDd/tMKSKbszS57BcTNgrcp31+
SPZmubnO01ty1LHwDHs/dZFB8a+SdYFGJ9Kyc43BPFK5IkfkLXdUGDJw9M64MKW2/NPEja90WyGa
/FhT4Mx6hS/hYoa+slVAWYOUicUlmyRNy5wHySk+OUO6GYv6JrwXkRH3C/8f0tolHj2dSu9PHeWL
FTji5jEZX4AWdkWrcK0Qq2GLLZYki1f8fioumP+o5o3wqUkBLpyRnFcWwknsZvTMdz3EqTZT7F49
wA2jjuKSryx3+1l6YxgNDhEbiL/UyyuoWJNLp2nEW9/sm6x+kLyewQ/lNlHOy9ru9TgJBtwEKDIU
RQfDUvI+9vO+jTZlEz1QQiHnPriTSv8Vt2APlNKZmFZdb/dGjVmBStTxuF/Cm4UyR+GCNM5F8URX
QWGh07gfpMlpSpQTjNzWn/acxAqH1YB9VYNMu8vCJ2K5DC+0VgQwJBu2EbLdrIqaMxz/6PWZ//x/
wqiayhjrYfeDGeH4NzwBBUIKzo5gDPeJNEY8rZ2Z24iH4ENhrEtX300tpJDmpRnlJVbvCq0gwHCP
N3OGQ32HB9YUXBqAES9Ljf+GRxko+yCG+ySb99tUzcqHcmuepi+/U7LclktiNYOdSbUVj+TBDWay
TtKGMUueQEf3ltqEbTGuZ5XfVs/1fzNkgRyemG16BhuKJUBn1YCj33qDzBVE0AL4eAqz1ccaaoLg
FrXY1E9ob3k2DIGNZXGXZ6C2S312ymbPUWj4KJYeJNFkN3/AxRLvcPRK0rIc3MPQa7XKgciC+hIs
pD5xmNaVAZSPH+OzZXEm5HcdhX4mstgTqsjJQc6Vt5/FJzOugip3ORuiyY2XcoC7LEX9K2Ujh5Oj
rx6DPmqAK6Mvxz1sxI/2k/xdGWRRJoGkmLgduzy4Ckb5jfagAfkDmDRpou+G9fuXpnGbi2mxpUel
ZZ5gRXqa95tGZnKGIpf0o4tU5gH8zDDmzpBQ0wIg1OGITQWrAfLygitfGvEjOtBXchqzfNvy7VxQ
X7tdyp2HRT9v/5JVgVX0rxFo7tXveBPWMiUpCE5PC+cvZp4kxiLfzenPVLN+LKiXyoGDKhAOt16u
HwuwNdSMD7ynWe39l86hN9uLMwU6DFG9WBXHKvbLPPuPzBY1KZQfmVlWtJv8K4+NuG6Tanhtyz18
5MJ2h4xJ7T2rXYsGIyP52yBo3s1/QVceS/fvA7nje6QUgm07idKDDzerZJysbIpRt4tMCa5r35W+
/c1y7UTazi1UNJ2yOr9BktBPJr7s8XrF2CuMCLy5bOU6xbQvmlc7BzmZzuPSu+lSY6MMA1Pvjx4j
LCUAXyBMC08H5uCVRpaoLpOK/MDUPUArmzaxBigKBIDu9tKJsuraDwWPoIsNpIstbRVYg2TV9JYV
uORXOUYrzhG6tz+PnY505T9eflO5bnq9Z6w3sNC7FzB6u5bw/YtKOVV6dm0erWSTRo6DvU725zXM
n8il5PIMOCg/e0knurXCHYCxCiwNkFg2HEsarz1PA6xJA1qV456C36cz3RppUmxr7wxygDAYliUK
v6BsPr1tHP0SbuF7Vw1r46Eva+73lbhX+AMyeTxsNPto/gvO1OC9YxWaFEN7PgWNHu1mOshcVz98
XoU2cZSnezsCWM7r+3q7ho8s/+QbzM3UoFPf66FryUci2zPv33aMbjabIF1c4SsPvHg5iCVdm7V6
dQRoYI3k+iUljc5YrulYSNpZa74FjVsJZXQ7NLVwyHb4bvJS2Rn3VelOWRsju6CxHo9LaSCHAnIr
0HiKlpwo8VTYevISw+ZB3LOj38ihFCiqAIgzaZ0SdtHMU46cQpqTb7b1NjO7q0G4nOghaS3xCbV/
7kNWl1wyGR+sYQni/K/expac1BPjOq+BIS6AoETaRjQI/+yKhBs6xDI2AtvYCad1z/36KL0MDIxY
HYeRuo1rD88P8SccZWvhI5NGcdgituOxZ1pJQla32faHdJvUhAJXGS6XV11WaxEinBxkdAlsZMDM
1sCsi8CFw554TEBTG2FmPRuOkbe6/E8rAzWA9iG/WK1I+5A10x1kSoHcrKzMNkB7ZDvHofVZpgUb
t9hnusni46nQaQb705CYq+85FjrzXs8xJZOf+rpuJ1e9Sv+1z9500042LYCIkH8nj1ekTczZzR51
0Oi0OVmD+e0H0SzgDeMNfyNM8IFc0UhccpkwcvVK6SVY7SbbbVW70rhwGa0gnj+Tval5IBx0vMG6
9RDbbZiyzxpMv2HErAYUbGSvE7hVO0qFRg2gz64H8HazxPPXyBFAP182VZlIY5lUcnfrikgJqtfE
EDX56jV/1wG5fc7jnKXAgoLyQGD6Wi6Qvil1nvFoxmKzcEptt9beqw/tXq5Kk1f1UzGJUKP/F7pC
On4X308FHpOiz/N6SsR9vv8paBSWrjHLz5tzUevbhO9ZOs8jnPFXJu2ejp2Y8ie8PRQAZXyYE/M3
rnrjXzNVmAC9RyNlUns8W5U+B2g3pyC/EnnpGZvQ1NgqZhdTr5gfPT+qUVBqQnxv97yMikeRQkpx
zu1DYqkjS4YSFiiwqZfYCSU8CWgrzBb9TFIJgQDyemKLMfZdTiyE+VbufENnKbmIfTtTIFMoCw97
KoxTFV5RJgcWpb2wnsw29mtcbqj3CE2HScK4NFNeSxucvJAXKr5s+EfxrnSw8SSmCIklRz7v1TXH
KFHg6MT+UpPO/lz627bK0shiE0j13T9iMdKcOCoYWnf3KweB5YYT8pwC96tbc6lC38hNNvlykJyh
Ud8HNYDGWWWJibCLG7Ve8BK7kcqyQ4hkXsqkxuBd1rcCfBHqIV7V9bI0ctOr+eMNmNFA/AjnWQx7
6Tf5mYsle8+qzB/yyMrkx4sRHL7oaYD1m7q7lYGTc7PXQGd89lNCBF1eThFV5qzeWpKEi4rUd11Y
dxupEBJZWrm5R4rrb87ZaLedzN37pSczkYOiYoSNFW/fO3QHh9Cp35Az7FhgEBi5uTrpdx+lhOBM
yzxYW/m2ODlAvU4ML+4RHvL/VZCK2NCJu/lZTK4X5P1CSIS1esS4hOq+yu374ziN64DWSxg9iGnC
StzTjkTtEUy62Zftpv/AcH6Cqx3ymwQoEHLnqBsXR5iHABMonpA+MAyZ8h3B707SBSDVyhThXs69
NTZtKYj9FqAU+FXQjv75TeYUntCugYj9CVIz8KqGk19yzPkB4CL7OcdZnUqhlEWffuNv80L7mRnp
t1Fiqfd+nkBVK3ScGz+oobDrJOMfz32jwCEMG4EbIAqihdcoQ0x3hRhghgS94QX8cvhv0H2ERZbl
rSMkLTcw4aSB84w696REKd9rIsYxKqfq/kMGlMXxY4iOPMdCfgBiEOp32xzpgnxOhQ+gkcNyNNT3
s64rApSZiIVM5ZwIZoFRC3FZWZqVqgFFnc/bRQSdNC4G0MiLrVSkJ2AjnQdagtR2oRRRAomo55L7
TPV0JdSYvi1Qf+BFOF9z9rGZlPCxLB7ZcOLtNB3/J3re/6J1u17pA/lq9RInaz2F5S0+QyXW3uv0
rkyzVqqhGXaYnAtPn1X5GHnwm08APEKar4rYZNTV7UdmwfqIYpgHVpiiY/A4iGaXsgXInSBniRzF
UfWMzhOq7UESklKKMF1PEw0ZhHbWRJ9Ba7z4YAuXC6SNgVREU3wbB+Hj0OhIMRlsE042qpARAe40
RVPqncL2ELLxDXXWAxUfacwiTJ8ETeGZ4P7QnzJ5mtWiLgFcfKvuKt7vSdajIOa67SFGRH/wtquy
lQ1j1yGwo3NomJ25PjRMxio/UIIWEOWW2km/rXmn/Hi3/TLZ4SkWFVRvtVR/2+Svu7RwxsOS5+AA
4G46S7Q/+gJLWjCXGc4ly/i9ix5iZyE7njM4NHYx+Qj/jCcL/qBKUc2mb5vZJg0jCjBiRfhLKT58
MOGsswTgvcXQbieAuV5HROlsVfAQ1/L7hjcKOoo1qQWuLiDU9NpluHwQO/MKD/40oFjV6GeEIWwz
8PiDjSr/+keyyz9E5oKadrdauU/9lQqdmcpu4DiguwrYQi8AmgONooZnUUMxNq3ebBOYNDOtfhVx
YQsueSJCyevikJNfLCd33I+B7cgELGO8NxVWCYRJqYzMkiV7EqOcNY+zpgP9mxVEYbMOGZHLpnEw
7ic6/lsaKZfjUMLPNa4dab1KOVP8eVulEyhVg5ttZwzmoAo/eS1BJ+wwvXFtBQMWJEff/+LEDxsF
1my1LJOXZSAc28sXFM/O01veWTq5uUdl4Ti9wYvdi+PFuowQbzbK/h+SemspFzQhDk1xNt0qwglE
YQtRxD70jhplQpzw/NjoGLUW//7t6UTjc87wImvFA/T1IpRHd1ovzf7KfxGj46smKK9tQ+8TJYBt
wRT9ryvhHlw8q5fedc/JbVsNTvK00Eo/ATNbZLIToN6j8IGMbNqS2Md9W3+P8cS9ruKsKt0NJG8O
SVEZQUASQwBbx0dU4XH09b+S5BLhoj0CbOBqhAjolJ+mPbDEiTLohndoByx0AFI2hzrSjqnZl8k7
UGvbn0tVR3Ff83cjfiyQ4xqGDxBo7wS8F8NcsBTurHahI+y/uAsPC//klaD8beNhf9EdWuBDJzk/
LzlCTPpsW3Liy99+lnh1iU7TIc8I5KWuR18Po+j8VaK0IgBD/wzFqsrNfNxDMeLprXf67kE+pJyL
CkCV3JX4KDtc0LHHYj3/YSt4KwpS02bFaENxUu0PBBKOp+77Z+Br1aNGCmTl9jNL1Gb19WtV9MNV
kUqcikMDRHTnkSkjm4LkqfAgg5Mwyi3AIFQT3Opw1dNZFcFHzoWprP2sb4xnH96d3PS6YuLVtBJ6
98F8Im7qSaRKdOP7tZ2X2Z79hgFOgqNQVWUu1OM6xR88xYa6o30n7EWovAIxRXKByIdxGt2LuAKs
AMVWppE8okdy9mohZxMJBFNZ/uyeCqqVwvpPB5EkLlUe7hS8ltfi+Qx96lw89GqFO7yboO/X0vpN
SstICxawLKyrQe2VhEh6/Gwez/6Tq75da2VyL840xsfdyJxMLi1zG2TnmD7jLf6BlUuxwtOPCS+m
2NvzFXCGdNMKh/+g27dQpyNlYS4TLktrvuOrvTYhPD08df8cM+zS0CjjJ1/FVRgBlJqgc+ROly0l
qyinBYnVnKsQl+emZR3w7kvMktKzxr5cGdrDTZz89bTfwoPFlSuoVuqkVo5XSFycsqgRgIQBsdYk
inlG7Y4iRBMItiAbEJq3Atm3gKJR+I0djL8+xaI+md5uG2CjmYwijmcPbnrDjIoScDX6sGulwWHm
aD0goQjidc+8YGYIM0lmznSEt6/jvO7XsdhxgwH/4E5VebrFVBaXsGuPfAzTIXhJvtD1wFqTXMfE
1yoQqEa0Yb/xBEEE4EQElLaAtCwBX+KObPhN8D79019jgRmDGAro6X1pJU7VSl3yln6unsfRLq2w
7fUd50YV/mMK4ouZZOpiMexBFvZRr2rxCzocowAqtPyBAE9+UkkiRQavolhrN5G4BsipiL9mkPvH
TR6NVnDBZiRlniQwZrU7+A3XNoxhKsfqedlzLdtJPr3NIzFOc+cLU9bTxroJcmW64bjnEuGHp5CA
yw7b9F0PtWeTBpN1z2d9JXQyB1PcQXAvWudngSSqDEmFIO/b1n7ry9SxRD4wSnYuddSB/5XnPhrw
IkTUN0Gk3hxJEChjamyPtnqwPO5T3U62dmiA6b/tiOzC5sTJrJS/LmRSITmec/5lZxZnJPHuFeIp
6vT4RxBF2x4RwWujS87HVnuQDJvslMOwmT+uicEQnb5L3fhlsbEa5fenIkyG8h4zZC+lnguL09uz
w7RSmR3l04zWTtwGHiKjsrcbiEUwOyetf1T9p39eN5W2nbxo4yB+HfHM23Jvm4G+rSc/d4L8ypkH
8d27Z9XnfxFM0NPUw2L8x/RMeXiBf1c/sUZs9tUfMBXMAXNw4AMZfnZ4Zw21kBBrVMtNWg1aRpIf
eEHY3tkSqSnmi1LItFUObyQ2PZW/ESVS418liNMwnK8RLk2DWpcE5sOEEpP7LL/gmkBHNzaQ7Xar
955uAsNFb21vjf6wtWMaL2zJWPE6raM99NG0Jx2Ryw3d0lZSc/vimQra7zoLj0MnYnVtuQetSACh
ClrUV6SXr8bjtfEHGt6p+Zvk+F+Bbd6pqdP0y0ksIv1102TEC6wuHyko6Sm5fFFYoAAkfJxJpmxs
q5TAk+0HWHJ9WFuJTngYY4CmGrCC0P/f0IrB/zcCCvDXnHDzvVYO9dR+tIw15pBQfVDhM7/or4Mc
vHt8SvZoaVfB2lDjsn5cr7meerZRzF/CFTTPzF5bPDBySzLlKgCmHk2nYTGqNbyXYWBQYcduoVyG
laSFmq6x799984KPF9RMVHy9Ru8ce1UiusvluSy/PJLYe/p7hPiClDeWqqKjhfh43AgKbaeUeGbX
unIBUoCJ1cKVkF9SZfFssyEwU2On+Y6qfeRhqv7limhf5Hk8hsB6XI0Oy6YR4rKLpLfHTCmv+LQi
eGKqvlwYnlBp/hxyS+mSIKYN8bfSjay8OQVJLc1F38bX4j10Dydr/0eu/tZTmMo6YBRPBHvIJgs0
fHehm6wdiKSGLPoDLSGAxafkAX4F0OL3de706TumI3Rx7wnJcjSje68DIvd/BuLRjaApLIxVRh9F
KkTw+4cIAxusXNCguf5KQfeImcOwNdv+3yC8yKzTLp9V19wgpX9gKn8534y7zKfZ3m/gK/Re6Scu
8mp8GzpJPMMk5UVP+aCb2VffpmbDYN4M3aG0JSVooBuCPT3iCWYA88b/kcygeUU2oJJ9Ush1SJQx
+rkz8QumUypNYFxNGMwfzHleIatHKZr0wQTabZTSEL29AkESWww7i8dHreBk1Jmhj2Yid/eCEqJo
Kz7SmaCEM6Khd85eaeAz0prI4zsKMrTTmYV/Ql8cCtugR+FhlzyU80jvYng6SaZxkP9qKnSJNbxZ
ycSFRsDbKkHrzd3QyK4g7sg77zWoOGC6eShDfMVPX3SnweDHViowH/pTE1a60qE5DQyGyJzWEfjK
5o02O8QzE7/gAf3++a8pJDnEmk75hgr8miDdLGk+uG5gpJfOvN4+Pktza5HD+Xyo24uZftC+Pk35
DSEoDFRuQEatCSIK8ec0D2JI5nz0kdrjadbl0Kb1pCExZT/9YiZbZ50HzLhkv2Ge64Nn5RHKdCtb
TJzyi4WbHNUlUhS/RqsLsuXOGHzSEld5d4lOYOmCdZZN+r+6fXiZKbZaVEaoMHVuEQIOH8v65k0f
klwJjmph6pyi/BA3Hy8qstRRifYeprz1+boPH8bcV+A/cn4bqElPOIeP5s/AmYer5w1A347gosOd
HCDgJJQFzxEGizP7NcATrOEJMW+BLfNmIIBS4WhEPcsYhKNfn74O/QeD+oIkTB5Y1zB9sSB9nWb6
oCOyJ3F6gFKrVoLS66UJXcJ5rvS+nXb3uqyWnnAxxaLjm81rXF74TgE0o8phe9DYs0yXmoPyNZc3
mRnyIh51EeDtfcacX5sz6RbH1DPOFD8DMorJTkyIeo9JNL/vsvT+M3FuSrFXqztDPSDlrFjihbYu
/mRiaH1dtEahG1LOr8Kln5TGKX+ExHJlOAOyju26frFX+Q1pXM3q4DgM2U7EBUW5AeOIi8DIVlwO
ar1Y9yruTjmiu8ca+odwd0XtxzAisuY/oDbcNOgyXqOTc5tqkxLfxedEUO6qsai1B/BbTlPWCkak
WgE15Dr0++LZmr9dsYIF8aXj5ADeMONxVcY6oiI925sQov3M6tATbjuV+v3xHVerVWr4N7L9gyTN
0tW8o6TMxiY9AIFSq5JtIE+li2aTE7623YvovlpjsiHKlrStyDnQLDtLi0UnSLyRQRswG3VDBkI9
KYRSQCLppdPTOZQmv+0JmrkN2ER/vEQDg8uPB1Q4SyoQ1s5TEhGJEyAMUXSID/PvG1j540tcbaC8
oDJHS24+3HEFJSUXcqfSzrc7VmeY+d/HRLj0YTu1x+2qBf7A1CaiOMdEkRBjMxZ09mAIhzE2Aznk
yXUZ19SEp4bJdZPuWceEbciyQDiU61YZzPFZ5YMQe9FioYw8UR1Od5rDf9FVdB1x7BQQiYAWQ5ob
FPv98jr62XkL9kUr59eNo80CCxxw/PUU4aaIYU2mr0fmnPUrfgiIOAvQfSSzR4dbD3d1G1G/zNbN
W7xPun/Winfjwm7RkZvN0ntPKaZ4nu+dufW9gqCj0f5IQy4z32Ojir2YpteuMqUxXl5Es9aXL8aE
/9UiFqZxGR8EGlPdQRt1eLnJUPe3fTnyf53xLmV/1x+WyQgl06I9eAe5l6wXrHqTV7TuvfkobEfn
yRvw4yMggj73WszbhclnxWHF6tXRgvb0mVxbX/r/K/qxN9Vykq3U+0/avxp+9S0DDjtRt8utmxEW
q4gOlQYxVj4Sj25VqHgg1gR2p7lIDs1I/6Yn3osUYNd9UeRrejJstxkKBiJTjSv9cwTAhTk3F44y
w71RpCEx85SxkoRwcm671awzSBakVsEtUh2HPNdAku4L7P0EWgKAz7JTAMxq0OOXBEm+nCbXJ6ov
tCnlnxAfSFZxh5r9kNjAch84mNHEfVeAo62JgtJZBBjuytiHkzY+Jtk7HMGLoKyqRlXM76Ys/aSG
B6BRIfbvEakEutuThDPOm351ymf4YdEpHfd4isNrWtTEvXT/e1+x6AiwLLiFdIewpzgUauB3FEI/
Tax7xBjbOR0/F2XH+BlMwJSBymqA0ZWEOaMl8ms6fK1SQL1FYzu2hxChjY/OQTh6afq+PIuLz99V
lhz9b321tWcAWgvlNIVn6jjGalHOMKxo8Eldq9F1mRjayvnjbdaFh8xYdR2fHImLVL35RvBdXmsU
VUSbNsN2zeBEiyuIETVPpq0N3ZH/s6fFERaGmC4YuRmlzNO76AZGnBWYn9fs9pAleJzmdUPdSoZ1
Bt2HeVvrLDueryt8yTJH+ZRvAS8QrbMy3WVql5Kbn1jVIdb5QAlajOp8D192tTj7Q2CHiTcyBJI3
9fmjGgiKfJEvGsx/fCIAoVHknke7OSYECCDMvj0HLJC/hS0BRchesN06HkC+dYDqYEVXTM4ZZIDR
mKmpnP3V6eL88JnOCzqzGZepzvQ8lSL44He1gxVdtNWNiDxE5TUVS/0DjyDmxYRfVnhP2t1tmDjJ
hPPRdtgFnkr6HAmNgAhXWfsJ4Daw85Ml0xYkRdbfeXvvNnr0Wc+xWuzhYHOxdGzgl/T9hEqNNS4u
bG85YIBxAJETmVRBrbWI6BqGB4poLQqQRFcrWotwsI8a4HVwTRk6i9gtcftLM7heSPFr22NYsg73
rywRV07IRnX7k4BrugknKpntYrsnMEi305loCO07gAkBTLDzIuypdxbzUk4csDBqNvBDbw/mpgNj
FeegTzjYWzItUWj+YVmljylXrngZgOoTALkjWf52IupIJXvKOF5wpkDGp5Z8J5JB/PMIloLEHTM0
Wk9K4uLMFS+daIQ9oadysYLDbZoOU2BiYIeTqCN7kyOmChmdRe9T4ChJ96wbTABqULIG6Ip96jjQ
U1dbPkMmqldoRhx5ht6KGoN/3fm+uvC/BQhZwCkmuc+TGyNUJFx973Pk77CYyKyNH5PY2Vo78Fa5
9Kp0fkB103ha/cbMuUTFA5lwC/boxina/lrsNqbCx+xqPyCCMOJ8JpMAJqJM6gFuHifkKdTVBRPG
FnVynwL6hXDLeOYU+XEhLUQYFYXkjqBV87o08vxVPwsRViS+n4qEW+ysP8uJEs3umrEkDukFQhtl
dDjttMa//U66MDxl/l7J6fKn0HK878XGLBWgHEUnOaWLJ73kTN8a27kMHOJMyWwqkxHUn5PGtBPH
Mqy0JyXpvD5YrFM3Pe3NJ71fW/HhOwIXfTLAxrxPjtQGJw4tloWHle0N5Z04KbDt7eL9BkEPCjGV
boLIHTUdtBg3jTbAa+lw+JCQBb7U82OUyZUsvBTylqfdhyilAWCEGoNfI8HJ0bPOTgsHgx4wqe9x
skn4SYvL7SWm1qc0TfdVjJi8+r59NFBcyG3qk/zLPhV9yebBeWPAmU7e5uj/b0EXrWHMy+I4N1h6
4P60CmzL2V26nLQj1YNkkSywF0UuaqmT4IX2MjQjuXkbbyLlO9veFhPua7l6yPhjxyp2vwYWozCR
QN1CgO5GT1h62Nv7yXILzkzSIgGmauEilJtcEebjx+4Klg09J1v/dbumru+M6iyVLz1RlSU+aQHj
ncxeASPJeeIoNlsnLDBO+OH5TlooJtcTIroHSNfEgALaXU0NE5PUUgD3X/4fKCcKSJGtUZnKWmCO
qDN79RC/pg4Fnv+TVCiFG1swDVTjDR+HPwuGwU8IAAp4tHHstQyJSoh81oELZVbll/TnExUCxDq8
gWbjeV5gbcNeDcM1PcCe41VT9qimj3eqVec5NKMlvM2DgANnPXJdnERTTOd8F9vHkwxBkmX0Tfbi
ON8SymR1WKL6FWyOWXxW46uQAY0L5hiBt6zULz6F1CLhpv2rrrZTC27C8HKVkoM+Is3g+8qanFut
1UwYLj0v+Mc3rALHDb/d2GP58RBVUCWcs9AfCqClPdOSKMgjFY+fJLo150z4cmcQ4hHNSCPGcnOa
1mnhsVrgfNqMTUA5mPqsdgp49xT33phBowhE0hIMEuF6tQ4IvBrmL463hMaDhpRrcvHSbOgNM7OT
k3XM96Mpt3UMRCxYZE4la1g341lAoQ42+5My+RMuQe7ExVLY80RJ5gT4TAkW/1N+mBmLEkgx6ah4
r4S/LGNCr3JiJPSIqBCqwoU0aN8eT1W40kBH36RCzmaRB+z8rW/R/5+YIYws+G7BuAjyYRO26A+U
LQiL7SbNu3zUtJyQchiEzYhJedysAU6H9HxnlirWb/xgYEHB5QRYvOpDh55+CaBBoQ7wHDhAqKCt
aomPn3mS22IYHa/3xYE+Z0s5tOxM/FVRUm0jHKW2JXlxtor5+Iw3WLrSvMPYAUrI//8DHlSHWHtp
9e8TrXJ1SrY7TAvkoZlLBbOewoSCQQHiyhL+9jDXSDi0H8bvKTQFsPMGrmsvAAhNldeSn4yHjoND
LL18ssdUN7/f9gBP5cKAbQnNNg4foFIrPQRSWP/w8v9+1E2cog7hIRho5OQuvq70UfYCyZV1q6mp
nBUwZdMfDzknPx1Zx3D8AP0wIRuIX5fmTb1ob45bzpKc45cAAy/oNErjm7hilR4J5ytJ4I8C22jU
PpY6Ghro4wZgxqf0c+54MyOqZ40Ru2rM2+WADxWulcDKFP2O7Pm+oDYNrekA9NM8QgYoYE/Dtjsr
fq0i/9kyou73o0GL2VS/66xws/rqtZagQRVZjCd7FFd0d4knowM6dkOFX5wQP9gV75ffH2IOjqKi
PgLN1lFWLbolrWyoaK4Wq7FcOLiOZi8+Sq39n3c4zG4/JABvTtKSBLvBrDBZihyaWtzDTtg1dT5K
LLLboibmbBLqd9fGKLa3Qm8wh/Cne0CQO7l/UFyvuufU5ZI/QtnoWYLFEqmgzwp7GI6xtxPupAt8
QD7Z0BPWMF31K5c3rCScN+SGadfXYPDhDe5Q32JXMwJyDnc73ZQQhd9xtidaZyPTUVRXSpDpDiGa
lq4LJDGuJKSh9Cqb11/H7dTkkYOR5nyzvNj1JkNyv1i2GND3nsWAhIjK0VkeprTmsv+q5zZr86we
GolzxGLcxPRA+/GY+nf3qMESHUAFc08LFPyBadwxNP6lPNzWwrN2O9YRvOmU7bzyfiPQIen5wW7S
PUnn+TX1bJypmOPWsPuqoBR48+E9uWyFEaTR7he4HFkkhL20UknmxhRzy6GOhge8dNL8vhsIlyTO
akgJt0RdYuY8ewm69174bCzsyLTHj/eFcUF/uViYT0xmMctJXOLumouotHNOKqSOdvSOvH9YIkZA
2tF/KQODftkkORKNfv7i4o5voT2g0Ym4I3/0ohgBU4NHaZOOc94gNN2dqBDOPGDInf1xvvTh3nw9
GChQ7sJDkKdZrjt61TYID67BWyu/l1M4Eh8iHYMFXbbu0yuEIV/mJq0T6kkpSGBf79B4vQySnZ/a
WGcRciwRTNMWA4bh21jaYKbrl+TY6jr3zcPEb8bOKte+mc4l+MLxfFJu5PwzPc+ONrG2JT2w8QcL
QCAmaDleh4Pv5Od7ySal1+2XqlJXKvsOFR2m1+P+FCvJWT/wSEAhOFO9le5tV3mqJmCjUPCaZ4NI
5Ll3UodpDUP7QWR+5iQxhMvoNqeDTXZ4CpTEPBxp/uDkqsOFH/4Huuz7cvONSUzj0X2brYYdvZtN
kMd9c5tbGcpgvfboDEzMzHx5S/MN0Q5IwVhIYI3/RpL/pS27QW5OWW8sFdAWA/qS+NSjNr7N4toB
DljHeOrfrC0Z1wGjgtbT7mkLNSEHjJBVBlLD55HDXIneRPoWsaSlnbRTtx1yGiqA1V3NG0LSO0Zc
5UWeG3i2DLUVyZBSM/9hO4RJPZGcmFuWa2zMT+ZUH/MBKpAAUHmLaC16mVfidVjN6jVGIUyalIaV
B2KHbVyKrDC5YvTXwPmCpkOmWhbC8/RT+k40Y+lhxD90fcF3Oy+PI/lpZASe3rbi6yH9pOR7INRu
Y/9ZyvZeunWBEMPLnFxyEQhLrPyzZ+d89V8A1Ocuh62C/LMYYjLmtoEJ/Xly4W2qLGoC1dekGb86
tPcOJzbK9CsClManaFjX1YpJvall4JTq4iz+Fo679PF1/m0Ip3WKCi7b3H2WY5d79yG1Wfpzy7RG
EB55QqLj+Ai0ZR6So4L8UkGZWxkLzPCPon9JL3nG2ybR27mXpSu2pFuC/LVZ7fya6adMfIU6IFTT
sXba8lB9+/FXaLAWzmvpsl0BdjD/oZ/SkMLGBenRFEFzR0ka3xje40O6i28zTA9Iv8Fqdm+VFzZv
Xakz1lHZtBvCbjF4DgQ5X5rzRP8PaVJoIISpGB4euqJIokPPstXOk7kMg/niSu4fWQvFtl5MAXcB
m60qgeX4Bcwdi4tSzTzIPgjDlEVSp8OMrDL1OERaSR+YAah1jLJqqlx7etKlB1QY2NoW6XD64eKk
sYPhvMMwrEE6MW5NuBK2Exf/kt3gXSvRPy2+Bumyi2hNZZrrvaIZG2IHM1ejh+yL2xKkj/F0QdTM
BMRL8AB8BDtbe/rwQKuIFNXgK1NrLCuNpxZ4JT7xJnUZBKly4LWW5gtbYNcot7n22Pk5MFZnZI4x
QpzmBfmjcSuYdUFL+COWBNXU76GuOa8jb+d9dFmBrgsUjDwpj9uFON8W+da1Yk4jIkLtB8rNUItn
MnZxseJx+GQ1O3apmbmUpC01dZ5s1zz/Oo3TyUC2tIfaAciUL53OtjwLm3xTgRRPnSlgDpBvJ5r9
TariIaUBWE26YABRo2uSeWQbM7PJRGRH9/6JwIeK0mZEjYeoQ4Y4GzMAGUFOoP3PsIT57WPq9GHW
EtY7Ypz+anqmjztBU8fw7MJPRZMwOUT/ECau0SudUpct1EO+LLqzgK85xRtM2ESgRJrxol4vKIFk
IutpTRElu6/fnfz2W9AtFcXZf2Q7eP64AGzJaaF2M1PDaEYt4OanWtk9VVme+jAwcm0q2+C6C6aC
AHCwpeZ82ADOr6M9m+pA0dErGlgtv4jkIZTw1TgKIYOZ9eAxBPmEqhUkpw4SdKdy289qedOlw9bh
NtqLxEsDugurQ6DdgS/b8KifTf6w1UVV5hL+WfuAmmxIjqTa5QdRNYcfUSiyQAgUH72r95hiFNL9
EBtIhed6IgvLUHFct1KrlNavU7Zs1+Eo4ksJC0njtmvwvEZUiN99Uxy9+dKwDRCfTtMBXAt6++jr
UNG96DSTPIy+SmCprBB2s5lURbLYgtr3TmeAdlMai6eB7qPppIlvE6mgL9bib0OEDbyJBg5O0j/I
CrtuGTx/UDMU7/S7MjfKs8X4l/gWEu1oPFZqX2FUh6JZ7JSLWaT3XMVwPjh7+IqhM5m00NM7lpsi
Ww+CUPcIxXixKIG6NotbfmMa3jSD76Y04uS5arLsML6vWbVXyleCvXK6RUGokWOR1VqBrCmh24SA
uXydXV/t/D/Cm/P02CRpJ1kirbBXGIfyL/XUkr0+DCbjUdmul5uUDiwp5EdL2Ke2h5xKh2SsTyHk
Mc/O3YUI2B5aAa/37zV2LLo1x9E1s9eydpVbJGmON4YgxHjbzhlRvek6hskbd8ZNxRsKw9bECH0I
qASn9zSwOn217D9rFbr3eHY8CCQ2G5oss8V/pZElQh1tvY9q9pZ8Pru6bvHFwK2EFhkE5MQvdFoR
qpj6oAX4Oh7q/uPrnMpq+iuJ6h13fmK1hfW03VsNvebBvIu0SXZaSyV6kgdt299dB3FXLTG3fMtY
4Jo4nwGetMEduAqqfXpOXDuKi/LPTnFEL/4fdJFFHKRZf6TiIfBQKaPcHq34B2DmsjECjMScSK4c
aUdGj6ZbTFNKFjW989tWSj8rw7jUvvFm1jF7Xk5gG90h7zkBewCaotKLZ+Wmi+2cb5SYNqUaQTiw
LjANjRgIblmVZaeQf/iKBb4xH6SCGaQBPKFEku0HtF3Vi9h9BxCGJYwKrB6H2kIbEfxSvU6Bug3D
UVaCMVktsFeSbe9kCUA3o55jbU8NlsbJ7OUEi7sQ+41u0sXOneoGmrXSzOltMcZgtYy3ufvpj66z
b6VlErV+lCoWVX4F62A2gfmn0NPH0oTnb+wEVpbzwZQJ4hk0Yn8HkgLJ82N2NmoOZq+iXAXgwaR2
Ne67m45LgQOgYU9wjAeaLV0xhVDqSitMAk5CMOw8eCpb7YoisX9/OPRGf0p3HG/+Teh3cPt+3Fzg
hLg+l467UTvbeI9mQVoQqZBlXpNkGZgs40Up0FdVEGI9VWK0mn4TFZkU4Gta5+wHWnbfNafHij+k
VV66J20cBx8WUAH2V5tqAOQQuX+Cwy22HDvhlnCN5onXQgJcCOsToUtIOznyePT6nrRYNOC2rp5C
k+0gRPdd7oCz+bOtKhwjoWIhgv8fFKCrALeNFF7EOAuVI/pDpaWgyfWDvD/ltAbXN86Y3x7EuLz0
TkZb1w16LDeWLw1VQmhRbdF31z1dROxyBZXtlY8ujW/yw5iYcqq1bhQHeqC7S1z9LcxjZ9bHh7+U
lq61UxOakNQ65jEV/dwK6LfzHzJM5Rb02n9f5EFcByDZ4BWXrBm+uQRGUl6i5o995mMX0PYxqrWp
VhK6jUlb8bbU5gHojTDdfkBnCD0f9dIoPDJWan2q35/hO57Mn1P/aq3eCX5Br6x+3Zc/aZgT2B/R
vS3dC23FHXJW7ft8z80/EmZGC1ZjMdRRTBwOQ+QH2e9a67OwZ9C5TCOV43f/JKsdVbXI3bt4vzyf
I4zHakPE2imF94R12sUFQYZOFtTcMgovSMjDvnGZEmFXUD0KApJAOHFJKPYRtxF5k4l+/fjcICHs
hhwb3izNJ+06WfbqsnPdnIVlxkf+zxiZBWHuo36cdvcWrMtfj1HJWJDiBj4NBtfWgp/6zLJ3egr/
B4R7Vsvzzw+rgDCGm8uKd5D/PlDjEwbl2H92eYJTgvw6/odkb0x7IYACj0HLmP4lGYdBR8mHM51j
8jw6IGkNb/Izgx/zXLuF2JvDORWAgPvaUJ4mBA0Wrz/RQifIarssIVac5IPKy9e58D8kQcHmb1QX
hJlcwf2soi5jYHevutMHdCIymLtJLRI+JgJyjCoWW4+F4LNQjKQJwyM0fSrMo8+zu22daz4seyqB
hT1Cs1KbiWDSSpj1n2M/Dz6AhUIXO3+fr6uyzsEGLI+shSNZhJnz6EEZCmeEUmZBiWNZByui+NIy
oLNPpjsQExZm+QT3t3Q3eShWbJb1GneeWf6+2DDsfvo2IhuvSKZzW4H3beK28dJ+mdP/AZM4hado
5BPqktIR2J6xYFQssrJtC4VM93ZY/80oHNNL5SfOP7jmtJwh+EXGrr6ADQxIdYZ5zM/lLKuPOjI0
q/P47C6d9RdbkAzXxiTExygP6wEBydiLimPLLoUFkxMVK9RXTigQn7NZgASmTyHwsVmYVRYn5zu0
zJSN4ycpyb0y+Wn2DJPWPClfMLjsMOAa+7UcHbxIXt2QzNwlePX/tGN5dtQ8lqH0GRW6ponQro1P
4VavtMkpRI3wj03DR4YBK7IZuAwrtp7wbjKWPcZxjMQHYYvyuLUYeL772SZo6w3wAZBTNv6CI7f0
Y62fKmDHHZg9I0cd4/tyxSfzwUbMjtuwMXpf+vJvQZwPtJIOHpW4qP56OUECesxZEPIzIMTSoHFt
EGspe/2cTRwJ4PP1jzR84KJ7XutfsNBSHVLPkm/ZfYhjafrcJyilMzwU7ef2qAdgLbHZipku5MHJ
jaBWkcfqFP9ywl5aqYtY00KUoGB6Y4QfD0oASX0kGTxauqFTABmN3xQ+pNeZJdoVn8i5YmXOozG4
XFEijMqzSuBV+GYWodrJBxDHquPR6V8wLncCwau7TomEmHJbdpJ2QGjltPSiK5IiAX5HMG+jimga
uCdWcp7heidVVDP7g3OcClzX915+rfbiacbdexv/t03TrKq0vX1n8cuD2vMEAGhEh/LyRXJ0SUhC
Q0oK9GNbhgw0Y2sm1hcyiGQ1PEk9VMQcx16ajUbjXgUp0/42OAPV7/OfBY58zbC0fRa2Fq8xddeW
9iNmCEP+55WCQRfbn1Sv0GUXOw6jKpzPEkoFe5n7iYhEmE3SFPcVn2thlnjkTRsoxIYrNcLfhMY/
A18nxtCi5bzjl+do68QYuRCg0TsnhoQVz3tp9NuMaKHnTkiX7ttGfi2fbsLXC0mNopKe9bB3OwhB
dR5kAKaoVKWJVtyZ6H6xHW/ODHe71SXjP68Q6lsb8qWEGtfa0UjS6WDdDwoJTw+6Bc5dj+eqoXMi
qP+Z+GOaAarrjqhdSWbkhg1YiuEhdnQYC5qHkGetRafE+kRPLcl6celheCg1IhR7iRpeNEx7HFvu
fOCP8cXv3kkgCSdbFT4wS8/fdlBeDQkIuOJloE7TRxXdmGH1lUbuW9Af4VNwlHAtmIhn2ey/Vktt
xdlCZfPkWe57kTYJibBd0TwO4GZXcylcsEbRsPCbmYJTHJP+qzuc1rES0s8db51VhQzYGkhXbsdn
XDTVKVir5NMoO94pro4tWLE2HPAIMLyWxNc//aVQP1yvEjBPDo0LysTVrWgMlGgiXHRyLw3N9GsJ
pQ5u1ni/jolf+4QlUpNPwmB5zYEjjq9N8OfuAwzHDX7Zz9N0YiGA1+An0HTcraZBGEorBBZy5Qk6
zQz3lRQufKYo/eSdAWwTx+O4MrBUv9nO63GvF4c6TxA41VZ0RI6uVemy9u2t+6+Lz7k04JIl1Rnp
6QnA3wRjIUnDiVcYHI5m9xeZHxdH7rSXYX46kCRTVzwRKrwrnMkdJfb/PzMWDQvu3iHknV1XMXx+
LvVuiE7YElCrO66cAYXB9nSQCrbZ0eiYK9F2RxQUCdKvGzv7TUPsCEl5v9z7KY+377wG/lqMwwlR
jsjdhaMbZdDipMqxs1guR27V3mdzSQ1rsql6ebHiN71yuLdcNjaD6q3MUdU9/gGnlRPRmwFHWjVP
VZ2zM6ACvqzTzS+ni+B8iLeVfu6cJNn/D/OnAWgLYVUeq1IL6WUOQ1gcteeNBHj9kdqDKZ9TxhUT
o66vOhjEhKKGD7jjyiRVk8iK+lFCn/kiGuCN9GiDWSkpTGpm0UuSPAro0fo65FEYKmL3sfqiweVg
Cyy2P69o7LErEuAuUflSdaH9a0xnoX3KcHuaadVq6bWVXA9XMC5Xfa9S6k8FXI3QNeQKa/++wCJA
g8degZv/N+AsvweBG7u6WxZCJkJTdJwy+h2Bj4nvISWr4E5TEtOz+BPU/DrYAp1XYHk8dfBlC22z
8t8XOPfx9zTLrW8F27cIJUD3rr2h3IycldVPAd5QPOp0BuGqAsp1NLlHReu3MJQamjZznxNVcV2w
wkf9FjhkOR35m1CrzcwEZvMybYXaguMRkZu64hk3rnFS+J/DWTU+HYTtv2ZDXeoeaOlMsLysertX
CFGOFqrJ0glFyqvPY/lhTo7bcDELAxiEDf/nmeOWn3u6mHI5gQn47Frtj1gqUXd8ugj9Or09veq5
2ucMTT+MBaNaCxHwLLR8mE1kTBz5afxEtUSQg/DHGdefTEUpWJMju2V3ptbzopLfiRSRmxvd6bYQ
mHV/zpgJc0hTufC2yutQHhnavAMd4P1/FqxHLLT4bnNCc+4OiYTNhB/wkIJDk2GRi46Qey80yj7S
oScJURPIV8w5oSKReox9ZCPNDyPkKoy6gKnZ9Q4QKZ4GEnx23yYNQkzHi6ENEVjqDPSXta28Vub1
29nTP+t7ZTMYvsokL9iBF/BkE5ZxuY2djGjuXSOyT6AmhZU4vbXselF0HEwFLBaj8C8+2m+4WLmW
U2S9n4Twf/4A+uIlwdKmqtZNaC7kbVHlDK37qalswp5oIu+7hGp9wRWREFosymPRodmzQlj50/yr
84TBOqPfbcyFc1sqcREZzHT9GZ8i7+/MFOlpK1iY+IQWws2JHo1C8ZDgxk0+cAP6QQX1NXlv93N+
0e4Uj4ejyyquUS204F+QrXSUrTE+RvuoSXQTji871zh/JXg9Ng6XV17J5Jn7mlBN193SzsCIPdck
PIHAtTatwoC253SvZ/BFVVmrZvhx5YuMhv5Oa+mCXyvz+w3h7KuAl0UHd+pWbgGICjatN1E5jqE3
uJx7moPR9+WU7pTRz8jsfcdZINPSV26mhu0TSPkregadt3wCVdzUGRq9cBdAL8IJ95LbwmrzxVxw
BodzPK7bAv16v64g7LSkZ5nNZTPs8/NgzVzdcnZUTjfXmOosdHwQqGqrnpwp/jI/EDXEcXfDGKd7
Qnp+i8kRD8I2wo13qTTpeAkjjnr6hpfZLLQG7mi2QN61AxQnn2UrS/zhlWvSYIgvyLN1z+oTjhby
bUB0JX5YHaT2yNDMpm83/ETUa8JmdOYd1ccsRDAJn7E2Umexp6n4wVKNb3jPj0NDsanz3otfC2MM
HJRnQbiMxj0tzuZQUGEvr9Qsj8hmr5zI8Lg0kHAPhvTxPw9BIg4VmyJAmq8bf8eFbciD5QSmOXzI
T8uaowo/B2JSx93thszAeVyDHcye73+14BEVtXeJ3CWDJe7DIX7YwXiUL3qqCQlDUFp0m6pdtPNn
zt51BzGv+aOr6Sbyw0K7G2n4LFtz1b61trep3NjEDDHqrrIGov+yBH5O+GmNaT9m24tkeaGDfGMd
fAW87RcoSvK6rVkS1HutRn4Rs87kyJ/mNb8RJtafa8vTQNcWrae0DQxJGNUXzoeyeVsgYh+TjAd6
AK4L0e5yV6d9jQslZoOeU2IcWAgesCMFlqvvvJ0ZPmuhJLWrMAYXQHoJo2K+Tt2oRlGYlojNSJEw
gtJgpgp3+aWldfU/qWbh6qbA5bPnhCFuRFPfQfQ+22STvwci9EscgbOfCPjZ6ESQFZ+gQ1D3mG5R
KUvrO4yjm/VkrcCKnnoTtcGEUOKxgsu4B8dmZmo+u3CL3TqTGbI/hKwOJYKV1eCcy1GaxyRP6CA/
xwSnKdppnUJKxhM4jMju5KGONrTlZk8i/VCUBO7mYs+e7RQNSJ8a8PJaXM84VM86N6ibDON0Jtez
iLw662kw2wIiox+lqq9owhO6LHkIEdHRBssoziidWrsWAPxMOKOEFzCiqM2EBFpdQextprJOSp3J
szcb5HdXDiIAzdY3FaMJfJqOs/fKHBrujcts1SBKXL52M7Q2NklPC/d8rBIw+rW+zwwmC3Nukbuk
V8Rz6FLj5oTC6MuwsmBjUGBMgTdX4OYHSd43wvdujeC7CrijlEwUkxy9HPGjvX7uL2BBtbpgiCNf
/PDR0KscDKFnFBTya2qT2m0xAlkpLxeDqj40v4VaRSQ3B+RrOygrcrEiQyyy8a5Asa3ETIcsqBen
AfoVDq/7Hrzgg372di1d2M9XaeEF7DrABo/FWqBo+sW+kJPBWKx6+QDoeKjscoR5uxrrQfLUm+Bn
uW2jpyj6LTFPJikYhH/e760Z5RfAkXQtui+8xy0HbxGaEfUVhBNZsQgqjq5GTRgkXBw6sKUWkcnn
PcXs+3/IuCM2NOg8S3u17VsQFvmLXX64aKNi3t7pvr9P8ygYStubLSrYeeYzCbkBSDlyW71MwpBR
lP+zKSIEP4GzXvDvZLDaJ7FEIbZxCxuV44NzJUuf49o++AOaL0XUiEuB+4glzIy+HvLONUTBJuha
N+bicswdji2T7nmbJyjGir2RtAWlM/4zNvGrpjyN+47bDU4zv284pODdQuk3sssnW8ZmOMMHaQqJ
bKB1T9ytAC1PjTbVaqw+htrCeHYsVOUqU4zFuC9bNmHZQTSl46lRWN0XGmmW198/tsViM9Gpzypj
aG8a2EJT6/H62l6O2t+s7WqRh2/TXhl2AQU4c3JbhFnNVpVUpri9lCiiXZUnZPpPHcB09uVn293F
TqxTeLLuoE/Ob7oFeecYQ9aqTlmcF2XZDLy9m/hucpCYNpnaNB7BHQFYlI4AxzAvLDvEeNpkqDZH
PsANpDxARNDWavNjEVSzrdTwoUymFSPUepG/xsOOx1NyOMqLn+W4Lr+aomJvVd2oQQJ6J/yprH/u
/Z+V8YuIGCCr6cBj/mSUJ/OoLHivNlfOiQqAoqLrXwgYXtj+ZGqI202ZkHaDWuRrMBjUOOeZtoC4
iJm6yVxXu4W3glVKMH7uJHYt0DQIDMu0hxueOaiaaeYvsY6Ti26q7GYk2I2zZea9YlGuRdISxt4o
RjA4YOH1xjQVhNujQUhjUJLjc61u905yP4gjb3SbHW0qF7kPTBUyRkpCzBljSjFQZIZkIxUBnCNO
bcMZQNTIBUv8qqYm6F16EQEkRPB9TRW2r92M41KbAaigwkf7FzlrR6qgg8ZdDKQVf/58QPNVBXw1
7//aAgohcqARZHJEV4+iH76nwjzJokUUIBYsonMfdgSLqArZJRUVSfowsa+5fftToLcHz41m1BLy
xMwldYv02RRip3+Dtnut8Ig7vgvqwsGPwEvTzvMPUSRjF6EMUHMGBGDyTbzpYZI+qmb9hGiVqi0p
mzfC4lDtFKlXOgksvduq73GzpLWdEuo0nRU5lwb3Hzj5mDnY//bdf7gryb382wgbF/9GqWCPvf2u
Y4xLqrkVG4i5und/Vi3a/CgLZIn43Pv7o+OL0Rlq9uQyeNKccC0Lx2LYHoyDloLtXon4Jlq/NxF3
S1s+H8BltyoHCaUG2uymvLNMIi0Zm1Qb+2Cs9u01YuMKkwTRfz4iLeZqdmAUIIFrTslUxuGnquFz
tLDuatLQ2rK+/gKQ307V8TAtMSYPTl0SGIHYq+8/cLTPHdCXI4311xB8LwXiIF72b4mVr/eX7YmC
kPp/ri3LCQtyVSvNisnh+GYNCixoO5YEw3Y0qCNhSxzNEaqx24Tq3yJ6NxCZQVTmH8xuBMoFWWSA
6S7soUJhhLurZz2/PjnuIsJRNZbOfC5xW+Z0ELCaa+rf6kqo7/aEpWMbxBTQcG3FMQclWLCQe9QP
4RrXr/rGorrhD7rrIB4jO2rAzhBLJaUDt8rXnHczCxAFwdHgYS+8c3QAHzgS0bUlg6hZmYoO6ULD
CUe7cPnZTTAdQAM3wCYKBNxIhfTzhalq7vojYJ96jfn++YzeoStnbulfpJBtEJVXD6vnUZI8uEwU
ItgxQ1ngbAJBDeib0yZYYwLpjsjZ6/MzkGZb25yCQqz7Ion6vOJLLiDD9eTDkzuDV8KylecLMH9u
v7orwNUcgA4nJbaKIkO0pKOIxvnEpSInUqNzh1OTznx6iexi4l4G/nBsPWb9CVILeVqx32W2P7OW
qGiFXCz7JpjRW8+mOtqKCsyhgO+mH4HRdP30eUud9FU8eOluxFNoTukyBFnRw0W8U3bkV7/3ztg/
F91KcRMQAuDDnRMioB+huD/GjUEEQ9GrU0JjDa+DiAWxvdxGRxXUgTf0UgPZbMmYtaleENDPKtzw
kfrxifAWFJDfaDvA3S6ZJ+Q2f84tld9I5pIu/LerRVHmZKcU2aXt/sz1K1B3mowTBb8of21YoDC6
SUX9INgign/KHYYaWdbK+3g8p1avoW081UrvQl+J4RKykzbTXCii24YxrHKjFhulsdb84k1W/egi
kvnLOLLxZGyzTga2Wqd3/T5WrEDuiEWiAGxz9wiGo9fZpBdPIgBhzYCN1/sJexD1m+jEXG1oTk6j
Aw1pXR9H5/RikqZXGEqLTw00BwOy6CDoj1qnaIxNNzI/e5D1ADz8zLavJboWysS61MTNoDQheavh
j7sapxuPRx3AnSrov+RFwuF1cQ613cC6rilfcXT/khsaNd48K86uUK9NK8sI3omQxcDMknw2dINB
kw/G4CJhaUadGQvAhS2Yy2Z4bhFPmyWZ1cwzik1kgkTaT4g1+Dz+h8JLbo6E+piKVK5lbBPvkXVX
6TPeAx15f7CmlmOiVE56YYthxBLu84yiuzrDbGlfshzsm8oaGJfXzQKKA6hcjHPBOEQEEYkf11wF
Lo45ctsYvniSIEUjF3uSG4qN46guMFjZ5xIj4MxEsdVigNyB5ApR2mlQbcK9ywPEPvxT+ot4hW+U
ObCTaqcSwrTQJ11AUwFFVHKZLkbjFYdBKFE5VKPyXwQ5MoQK/oNI5Ssmge3S+Nn8zP6f3aqR4CEL
FPn8JYKYStwaO56yMXrg0c6ozpUY8YQcnOKKOUYieKgTfKkakdR6mUbZQBB5PeDW2wGW0fmIYHQO
4BaZgfP+37bQerLVkTYnjfmjWEpSuV5kemCUjyXPjit2nXjmTDmer8SyHobmImcft9/TBh/ZJf5y
+3i7gOwPpWiRSwJlmqG4U+oa6NMovYHKqxR1enw99dUWHVU/kTr2J2CVW6pGkbZFMDUA+XF6M6yb
NzTZW+y14Y4CLkzbzqLrIEAw8IcsQkGv6OXvfwe7mWGXs+/pczkzKkmW8gdthr9TJml5wft6K4AR
MTbrOVdxSm5LAXHG8zaDsJOPZohxWG90gJne1LZRTQd8RQ0Xam+UjRDtBosM+Bdc4qt9TP7nRfed
MFfu+HPNHGqIcFXSOLyvnF66kLUWxJQZw2LJtqoevDXjXPLvYOQwbpm5kIrGwO871LK4eJR6o4x3
rlAb1mRS6VoQTrS21bkd/15FJpLF5h4vV1DNCZx7hHz0CH/arsw4NuS5uA569B7P6TZUNPO1pgKl
/u6HtgSHghDbqOpPcVGvIVwyFFuFsgToICC8XpKlgYKaysMnR14la/VbLUE7djCX7QIaG36VgpG9
3W5ghj7hAlZBbDW2kpHei3pKUS4Aw575b/APXH0pZwJOTUQGfzTrquvpGfVdVwFyMim0Y4QntyPI
5UgyuRBfjAZmQ2qoCF19F0K86ehT7+zejWCSmMHKM/QHZzEojzawy5uSXPPYSCooifShYIzjlUIr
jf2XfxZ4Uw0XaYbBWJQ/VmDY4lTr8guY69oFLNZ+HOpdUelgEeUW5wfFnjgKYrP9dVAEKDb2vkYv
+t57UeRbf7svYdvz+Y+Fv9UQH76ab4pm6qIFanSCw+KjAh33EXljy1V8FIvJ++u3zvKmvyUAIHeE
2sJGyvErEd8ODbvDYTLQEhALh0Al2t4xjYVR6EzVKR0bGlvnmT/ZoDKGdsjdPo1vbUZbB0BPUUuu
+nJWOp079mxFgK87Qz//8EZNeg3zHk2ok3g92i38yoIO8knwiaqZxBV9eFqYhC2DiTlTizka9UfO
AcVtXZwMgErDsWlXzwlID1Pc8ES+y7/KWOWLk6cn3E3WOMer4py8J28jI4LY84vuMtmKWcba1fI3
xl98GHj7kZvRQxKDshMBEePiFQ/7wxnKdtHI+Apu3MJHDMifwvK6h6exaYF3Jb1qaWZlpN50pD9F
cLjzN9s0I9oBoKMXzh9la0OUUGlH1++B2GBlNZNWuAvPRhtFNwSnKW0221SlMIXrgwYU3J7TrYre
Sz7ETItNdenJPsbG7zPNI+uLi4m1Mkw5dgWrecmoH5gEH4nYcor2JSfRGFi2oLJ7o1up6XnBFcpj
oORjg+MVwHCCLB64jZDPDWY1pPeNKUdtmnjL82jBEI45HFs1UrgYAWeUZxJ0Ts56GNw4Hpp5XFFO
zfzCls/GLdcGqP4P3N6EswFXU9KiCpLIFfJizu9fYSd68/UKIL8DLOqON7hnn+3ehV5Ll+yGaD9L
glQtsM4qF6S41MsE3RourOKgifYuAsg8DLUTYaM49xT3JFB2HGwhYmMalW7gmq1zndHpXOdqMomo
nbHju6pc1NOR/K8tPtJFtHeER7VYO4e93l68fzbsJ8kzxCjotTGzCJVGTgY0MGSo+R/irByQ05GV
BGVvAHkPJCOQ+kg309+wqjl94pucgyHwCSk17T2iP/eaBBXoYguM2ix/M6Y3JGDHXkpGmivTi1c0
fsD1cGgns/9iGbaVP6u8xqLuHoL//AfRYb2ooGT4nOcoqQCYlL2DgAUcsNRICSzuvy/lTf1ViqA+
a9Tg+gzeTp/9YcNnHbyNbasQSUSdaEuVbqPxptQ9+irRGkfxxFf9q/x0Qx6+hcoJYrH2c1UBnbGf
wmFNFCrGiIIprrgBI8YnzTXXxWxuLlz1JUqvW5WME1k2EUqWmE4HzRmYj7rvpF7PnXbC3nGRYyWP
gxJGE5GkKtRy0sxIpoeCafqX3ApNIba9D4fWsMixPjs44cTF2mCMFj0xTYpVx1FQzXDlBOHHBwuh
8ro2Rfo6oQH5M9ytHlsnThK+cFeouMSaBDwqrKlALAmxEY/5w1sKKFt2gYXtay63bzdnZ12YKOZk
iICgc3tk+BR10FFilnZOdHr2JdkhTCxs6jfRRErcwAxwDYRZojVvhysyMH4nMQ9RA3Uz5oO3dHfx
6nhTjx9ttJTM5IrXiNm/4JaXOLcgl46s0R+SQEuGNTB3Vz1JsExb2utxUFQIK/DpTOcV8Z0xuDu+
6eKFFaAAeZwqslHuky7NiFl3JWDFyfOXKdysT09hJAfejOQsrY6jy9nN/btqeM5YwBNGSex7APlr
rDMCaniyGUAEhooRpAeep5Q0ygIbaR0hYVCcLT7LV0JEVI3RQGrE3SEPg9zguFx14e0F7MTNGIMb
npL4z/6nI/D6h/b/0FBv7kvIxQJf6C1fIMVaSYRF27ZdRou0GX23TfhegC57RuPJ6JwYHKTA7QkT
m6s/M8GoSuLaZ8wZqP6YMTyOxg58b6L6qMGa/Azk3sQhD4KkkFWciqYanaBtxhOpcMoEhl0TAJwr
XMp1ve1X4CpYuo8jQzGqEIZaA7KuARwshSyhQqDd+RJgMh6b6Y3OjhqefLSKkSIHMW0pH4pqJmnw
EK+A8NN5SLP+vdsdQnHxQ+xxqfMwN0ZnPxe4g5LKPchUv8dHixHEDsPLgGD+tEm7Q8ogs5YhWWlz
yzSQjwEH1HsTVDAx//UZj0ELg66/porNIvADV/5BONwly4wzMZrVjf9QPSlj8su93T1uZJyLIzX3
4PPBW8/aMLQZ2q1kxzpfvWUNS7Nj0z9yroEQ0hz8rX5a3djAiGxq/2/YNFkBVJHbJa8liOhSGP+H
UQU2XKUPuMvpBy0nvcoLOVOzzmjkZ7u605ZSaKxgLXRtxDalwb2/jfv+vNmJkTAhymCI8CmJTRVj
xsBORHUlUFQmRHQBmRMVxWw3mH7mE8l3fTeoWmKW1J6MJk+0NCqx6mXgFzmXbUDsCrp8rbe/ZqZY
i5TDAH4wU62DV2w4pR6Nn/QmKGkXRVmv0rxVGPSOf3AUyKlVx/Tubib7pMyMY+wZ7xTGhbfJIpbA
rX20IjFJ5YWhaqRdRCQt6Py8OyWCOhzavXqH6ZXncyT4qDKMG/Qt1rQYA89NkRx6w91auV7g25oJ
9u3ztlCJZeYM+VaXqZvwaMcBAJtrOWovnnehsZk5slleCcah5NjuHbUlXcUHJf6fUg3KnNKr4Nyz
JJta2zcoZo6+2eINvWF6zYe1Z/bVdf/Uw3aGf8vjn2/J716NOyzfQTWw5oTQI3W7LEiLBpyhCThb
0Y7ek20615BWUPfXQyWt0HNrW1eQSyGoY9Wt/a1NvDnmmmanjtT1D9WqbVzUH7s9P+X/SL5/1mL0
RxpLDlaIBdWwBQfOlGD1C2AMriXoxJu+u7Q2pr7r5u9d0uF+P+N+dp+zsC4YlKzZuKEaIIAyh1pC
dydthLMtG6a5nPxJTgulLBJKUZnSTxQP41R7EtT2kIvx9dPWijUgbMqwt1VHLiha5Jj1vfBe3zY9
mKIplx0QPzO6fJTfxZ7w0jP0vejKz6+Fvs3HIlsU8gKOqgPUkSQEdR0FymSrYYSsp4o+7YpVwdxi
mYpnB6sIpKuBaxIpjLSkquhyWQ2qgZ6YxcDVnSicm60kD46ZZ4hkbeSlJj2RMWvM5dXZ/gQa1kyq
REOSxXDbNUgyLg5ZseGH+3B40C0J7kjH+ZHB/JjtKyBZ9lJAMmQjwJRsB/tpcBEFIkl/qKfXU/Jj
bMJZJVmiXbLNAx1D05n8JXBDP5/f7FpOootNiujMoYQTdt1GRjxrACqRb4ytQr3vGlyuZfaSJuln
eF5KsBzoHDiIOQsBHtOO60mBUUZqEz/iw+jb98ol3ziqZbdDGBvp8usLwsa+p31zKg19k9mqn0EW
mrLdECo9vT4kuFlNLS4F6epNAfMZzBjRbP6duCuO22vl8n1/23d4WkhOW4eDlXsrdxkcxYcgD9oq
0mJ64ifd02MOco8+AbiQCSiUEuwITpwFvYPe1gboO7TICuRIdMDeELUZsCN5gL7nhzLIjxcF7vxe
617tcCah8H9kjhryfzaz6VuLBIMkbU3FpgxIeIwHxCYNqI6bEltMwXDBblOTRzdTTRk0duxgeOJo
OElfNb5WEk/DTd1QuLmVxa5iUML2pQAwLdud520JLjVVfDQJYQn5MhCvZaywyK+m0wsLp02WvJjf
yVDnb/MCbbwDIaD8DhfQoiTFJhfv8wvpoqWhWftofU3CsNRKUQmowye9OG5Gxp5lC1LoElBmy9xS
IfFtNIVPaUlwlGnD0SLSOh42hHMesf3VDkYgatDeq3AzozVhdfr1foqb06F04fA/aD58G42wEecY
lWDaUWmNTleK7xbU7cSXH0y+D1E5vuXq72kh9e0lpabwxwGOHjwNnw5Wyr3miZAOl5LFI9uAS0Yj
Q9AiddCWHl8ZWgpRPwYBLNCYjZp5EpXLQqRT1AGpafT8GQ6qCfG2ixtcirXvhsueYzg/tDyHLWEG
cVF0ivzcpA9CZGehcaLLhgSIUBBSDAOPczpuNWYCWDo5CJkBBlRZaHaP4Xhf5WQYzXIiqhL+J7fD
6ntUdkB8HXz3QOTa1JvjR19O9OAr5DCA3BKwlBVttGSFItjtnCSu49qhDrnmFC0fd5kbnUsbCsht
Z7ruW/HxrjmwaSos+NPnmzH1pYNte4+y3OcuYdyGIhPiQjoFaUxP4AX6unx7E9E0NSUMgQ7SuBRo
oKgv9id4UFXSeAuopO/xgpphNbcoa+81Mv6YyF9Aw/g93hMYVENwqQ93OoVhjYQlcNIcCRwG4q21
y8AWlDL0Luoc5coNiH6XpaglRf95Z+Wz+8JnIqKxWvHdHFMHEeXuwEc4NUH4FhXvs4DibqgI8XnZ
e04ykztBIdiKO3HYtZV+Gu1OKeK3jxY0ryGozTPTlNtEIVrolOHqWkcZZCPb9kd2arNuoCXhAtHd
LvRHnPhtBNJfEO13QVgnJOGOBeEfeLOuj6W/RmihJBQHHOJaVgFKRqS3Bn5yFNG+5JQxlpbM+1lk
KOrAvnRTYJBpCN2+KcjnGInL5uLJNYRgfeekLgYmR8kI9ppcKex+gffga0xZxZSYDA7+NBIOmPb9
S2ksKlHKNnmaXi648GUT0/LE0GQMxDNDtF/omIQ1ckOZInicPUKcf0nWi2WMVg+lfRyzzXevUSfT
r3gYiwoSed0wOum7tjkbPPIgyCOzGIXTTPdsgKp1KUdxSy4JmpIhTZv9sLgq8wu9kCQwcUhe2CaQ
HQJk0b3sbpyWqdy6NHSVVPBCk42wfMnM+Z2Ez3wIsCyCjW1o2nmuyhJouEu6ggP48MtFXCezzMxC
swh/bplJsUdf/a2SJ+0QiVI5ohZn8VbwN3eI2Z5w1uzMWkN91Zp2PLqFKECZPBCFGpvJyxpufFYO
nDm+gKr5Rmrut4Y3B9USogEp8zhwTzEvM9QKp4wUYOIgStkl63AKN0zyn2NigqB7H/lIi4wNXa2y
CyFYS1R7U5392NJ4GUu3YhZxhdyLB7/3QCRzWtWLroPCyKlPbdpqohhaN0rn8Hr2g8pqj98kp7Cs
E9jva++iZlkdg1Q2+1m9kzuRzCBi+trmCmtMi7nPNuRwY0lq+ThKlCFfJzUr+E06NTGxx9y1BvMA
rLNqT1Bpugvpk77K9rEbVP4drEuBDkZ3RhR94GsFV5I0kZX8YVUB2y65Y/ui/ZcJFlOroAE9+92Z
9QUCnFvNJD03mJV0HnlzdxQwqEbUFChbDnvTzgLFiS4I+rPYeBwtpt6GkxT1BDw4X88I1saDETNR
n6Bw0XZ3SJwPFaNQhtpCvc8SSW6Tv4IeqxWUd30rLUvoYyMYG0G8+go0PR7K/DWyS1TVnUFyJQTn
freAFw//Q6+Re2wWq+MW2M16v7iJqn4ec+yrvTDuMRUqHTKB/4hVw7i7FL7RlTjeGIrBWjTkfRLu
Z4HhIA0DfsnOl2BL0RfHb/EY2Bn306q21nR9hi5NwbnxJgmfNHtk40n970OpgEmjc04Qsx7bPTdi
CgkD2bksfZBj6ckhmEfV/One3Tu3yEX69zv0iEM6DYWbTUxJxMwBJIPKRxtxj9liv+7XIPYnB7qk
rNSGqNuhtOwB/wrDqOGeTmyQy/5NYwveUoN6S2WtJ834clX4yPYNg7SjTTeN6FT4Q84DAxihNeEa
7nx8BqShPjLmCwBgtdUBT2x4srM/kDxpbE5fgjYwuVBThDoo4N894TC6FyjW29zGAl0LL8BA5vhG
BvgZuXeLgE1IEmYstQwfv3mY1rq304D7no+Rcj4xCY1IIzZVyR6HMZGPMLFNeqzcRaLLdhgidoan
FiWV1BY+Ys/VL7OyzwypShFAFNCSnV3pGhe60dJyFWFrxUqErnKLEH2/M17oS0p91ywp8xLAu6/K
nCaOZgCBZ/s3pCfL0kJSxB4K+V38IG2yQoChj3h9adiT/iQ8UFRlwx9vl3QCIBFKmQeK5GKW4EY0
qQe7JQd2HrLtpShfU6+C5VHcvlvRgEdfUeSEnvnPCWq1xTgFTi5zT2S9ApDU5c9rgoldr24vG6rv
rytXZVGxlwZKzGrjuxRoDsIFQLmRHqF43lW5T+Scq7P3enc4ug2P7OLJCbpMMkqC6SVzPdp9YgGv
afDPxkc2wFOtHZ4BHY1DQ7Ozz8c3dfN4WN9vPdMUoAkaZDzJMFHC5GdkUMY+r9FNxvAXmIW6J9Fd
rVKIAFD6Ds07QAx6bsr2aYYbXmvOfDIHFe3PyNcwD/gBQKNrM7yF4rDGZD/1NILHDw1p2ptTb3F2
nISESQastl83l5pWaBW4EaIQP2p/Um8cQUyw2SeBsNuA3GVnyBBnKcGo8vgie5Nnbi8M/grI5OSN
0cmlzBrDOq6a5oeHM1e3H8djk827a/0bh0yPf5eF2nggyfT7CZxfrEUc57TrYdY3JxFMXECSIHM8
XCc2REa6yj3ORCTLFJqaUb5Mmoe/s8gxo4ycT1/Kh7J79zp410ZqPh70VHzW7FqoGFCyewvssXEK
iQScYTb/AnIMQ66XLxiNSHrfk0GJ9hUGY4rtQNq56PaAHrh0uNGYQo9ZT6WNeOOzRcWbuqTNOWhR
AcrEzk8cT71P+N6F5/kzqSwpUGv108Ah/MFpdXOafZBBsauc0AeU2VDd6Vq5w2BFuIWr3xf1E8/G
tGJIkIFKmreQtD0umqU81v6PkkpW8dedeyVn20uS00FM1ZvJbSQ0aqDiQnJ5WIMFPNXRGNTFlweJ
6u6ZAAc+0YtqdqKVYRnhfoWmHWuK7qHP5tPGqUMVxVIapg9bFxmSte+E6JOl5P62jphnmK/A1RFZ
FvFsld+GVSB/2ixXYFIxquJS9Ypc1K8jpCsbsJnrYFKlczcwkmihLKOu/ojDtin9S/rx6stS/Dfo
nft8jizhAEkzt22Njs4uTEjEHD/vHYJsYalTW0IzI8hWEzqAsh6PYFw2XgupBUJtWXrEEd8c0qFS
Py2eDl0j83IseKv3DOYNyfO8gxn0Exc4F+/yWSqNKbvNH9woU2WSBXKDEoN7Ik2XclllfTaudTBu
bAn/o85rjsl15LD59G3/qpiqxbxaqYTfshX9P4IsF8nufPADcpm0wQNp8j4pgnPb7xSLoAtQUZuE
HGeVTshg9tXOOEANIOYW6JLsTI6E83Bvwxbi8GlAU28cD+NFQFiFz0VZMKQqESKP1dsjhSG2sjbm
bz8rJXHtXytNU/nxr+0gGB15cq+SXajGEeKyKgRWINz1fmYb3zIfXRjh+IgrnLjuRbkQOswxBUbd
9ScZGi66QVH7DPWwUSQc9Koe7ItuAhNlRhZ0+Pnkvxg4ftrBJtZY2YJ4FTnDmQOklyRt63dOfN3c
1xsneut4+CoSoRJgm2KiJoTuhIj/mvo+DteZVJ+2iTkLfcVoGqAR6868FhbYEbnYVbKIKsApJU8J
dnU7IgVuMFodlWZCk7MA+/MniM8OQdc7IwlvGVfhBco+mxnOX8DIuOoC/8JgGwNTdkFZwW0B5Mnu
EwBz/Jph6N1PJUuogYxjSrWBXhxJjR8nyVzm+mOiFYwvjCVJBAWA7wlVtviuqxYiqjkU+sDslOt2
9Rfj6LNctDUNKoKyuju5d/Sfm69ltt9qSCCtxPBKDsvoRzW7GNnd5ZWCLjAo72gN6l6OCCw1ut+1
hhSJ0vN81e/lEo0cwfe1OXj4FYWgEcTiscIdXy6dLUgoWc0hDatfYF+s8LoH6Iy+lBd2ilfodims
aQJUiouZ3vx+siEUYvy813YwkxTM24tpC9oGaBgYNdoVLgRAa2Q45EtYa0A15ETMJNFWCNPMniXs
YK30lAQ/ydzjxQbHiH5zIskbV5Odm3535UItZuQp1azac5Vr6hnpzes8t9rcjuJIVTAznPF+4K+l
3xK0GFOYzrXb4Gmdburt6nZhvQeL3zimGu2okm81GXL3ap9fpR1lhGawpFYxNQEVitsm33WEuRQK
EeR4TVEpp/UGjarqx8T6nYBwIiJRf6F+1Ljf47wdJVvrxV7BmFcCd05E/toQvj8hLTL4H4abTqpt
l6G8KGhAdFaUUjI6aWG+iNWQz4CCdj605w/2FB+ulF6aZ/SqoDZONfQ9D+NaDQc8ab+IRIBWuwuk
FPn/ZHRzx20bzRMmgWtuyL4ppH34ulooGHRjDGML5JxvhXzlFsuhLMP9Z948zCHFcW7UkSr0WZee
s+BX84/YqXAShV2OZcygkjA8VFfYsEXkCDp9j6rOFNI96RWbPQlYo9fcmEaTT9IGS6kdR3JJMhPe
GcV7ge6v00dOsQM+o92fLlt6pZ7hbQEp4QkAgMPY3IFhyxWrgVjCPnH/kZcHSaUpCvagxlTF8ghS
9a04XUXsQzA0wpotQMuLMmOHfFQAFUUMQRKw/4BTUKDVyKl2xrQU7TJlYPUu8KJ8LkcgnY/SzTH1
zM/pYOcDzUrzJnIo6Qady3VjPES0yuW0xzHFBoEtP3eAVdE5v950BxIBSM5mzB4/WeYwr8XNM1/B
R2WRdGdCmnjuzuwMqw0Xd/NvwT/ydJKt2rQOIWOWMoAKLzauNR5VE04OyTK/GWufKSd2CVDyzrU1
j77FPfid3uc8gG1IWj+JUf3+dIsn0blljfZVLV68I9K0Pudo/Irk8SNVgrhandzkLbKpnZIkOibk
DLUP7bUyw4OFfRomePaphBxE8+Ve2BjSiQsItSHcO/ed/y7T05GTJ6WIPXEdOBlwfOjDcrPHgtaz
p841y7dtpFetAIUdCb9aJmAAQVnXxyyPzqYlxAZL8OQrPXfiSBnqRjCs4hhWip50McVTCXlnHuMg
5zdGUgIaf5UqDiMh5PRR+rwD5QTKiG3TJQ+XQUMIEwN0c8kUgYsktYlnNzJl2Xto0Hk9xWM0rGE5
GSk4oaxs3u56KKlALFpXHnfwmKlmLDc36mMhrA9zAKUQEU0s4gcvF47ld2BTBqZyg3dLED/2sTfc
v3alaWsoxhgh9KvnNvcDM6DNkyf96osZyjD+yUp9qij+Szo3vf7c+NOcXQDKJ8eLtAakoGy3Urj4
mcZZx5UjWmOOouHxUIHpLfVryyGEq8BLSJxEn8ltw2oV/9ZrX8jWvVDUTK4gDsXQ+52nAlfCij/2
UXholwyJOOskwnC9sXnhzoRJOUVM9z76m3hZi2oQtYKDsL1ZsPDDlNJzs8Fm+zfHrAQejBjDr4wz
7+AcB271OSMg+pRWhxlD7HEeO5wREl0tDjPQLavvbZthb2ZAOF1shfSyoLHYf9/lluutls95Izax
zvmTs5kpahPEjCMFcj0fqfUVvLHsp04Ang+5IDH51cycsFeKI4BOB/Pev09GHjVaEJa7z0qddeSV
q0qAKVVfYxBm8F7wqvHCgp2ptyYAYVPyINN8XjrlQbbRpEq5qbFKIapzBiExJ7ir9peQR0sY/OL1
eKzUYG/8yPXpsoVJyza+nL8FHF10GrqSzAO2h+vv4/CxTEWnEop1ohhZ5klLf7BKhx+4LW5yZYSX
xYeu9mzEYzEPgEHmFlePYrBBi+FvwYNGptqRM1d1qsu0Cs11tO0PbXErU8dAl+Euu3zw9kaCrNtq
bu8ggBH0BGPkx/51L7vS0T6tLissGk5L1WNksPTrhOECScowrmUzqCF9+SVUWcjyQf1azXHHCtZ3
9Ju4tc2mm6n2oGrf8BtCzUifstFIJABFPy74/6uyLoovS0L0IObFo9/ghz6A9D3X/mzcR1GaGtCb
LoRgob7INWhjzBpC5SjoXeohWr+Yx/j1meS88/fIUpBlQH5CKLzwhiO5Y3EmB8pOkcB8ADFuFa3W
RVSzlJCes5icXuCnN4DZ0gy0XzxqipDUldhJ8mfSBaqVI6OZrCPUAUPspaF/vAJEHuNTaemVxN/6
zHp1L6LWAFC0Hz2hKP1f39/g0OYGL+bo3r1k1iDCZi0CoqRegRtepKDutw3CVwjfO2Wuf1vXnDFW
2Y3QXovjBHzzazjkuUfxFHY7wc1poS022cEE9wFyeCBRatQiaGoqlBIW2U34wt7Q6dSDOLsDBZPJ
FJ3SU1EizNm25X2oDFUDltoc6tSy6NmQ61kB5RYWxOEU8+3UXMBvapOI9OvvMMclNUus2ZFDpRvz
ZhHeDoYEnCF2K+46oZ6tbSF7bPzVQmhujbiMHKneQUQSjdn4axexWKGAimi4hzLDDGO2ukO22KJP
yvkkQIZf/t+y7ciIoR3tauqy3BMAM1ghnWkr5MYJhkhUgI1OGVDeT/J8OwfSgOPUwv48mOwf08Dg
UOD6608cO1S3CnQ2ORyfvmCiQvVXuNhYw6qCmQgzTshgjp0Na0dHPRW5G4QifkvB+kxIzMPNlv5H
5ux5ndMYO2e37hBZCYUjvbDNoteUxUy6Y6UXbFzR0vWP4f79UAb47e+GKWsksDW91GWC6tYlOQQj
4/deYaDak0MImw8Lkiz2Zme5XrvZG3mN/wULC3WXtH4HLwmoPkZkoRaC5QWmCLt4GcMj55Hib8eO
RozhcIGyGQVV6NIYG5w/jddHzxpyefd8XcvC/Cr/QzpRgDyNu8OdunZDsp/i/aK6WjVHxxN1B1B5
7F2omXInOgxhtYOplW8ZVD3YX/7l2GeYFhqU+ZZY6KhilpeuBbUTaBcIImfAlLxttolN7pYcAtML
JJ+4Ky1ikQ4DWLZo2kRzIReKBeYHR10WTkzXnzhtFdU3nkeMhpVz28vXFWUz6XS2DnoACszV6/nA
8+eArXm/493kYg+7PYUVqzgbeADqVc3GSUyBiMLimyrNV4XM4Uri6UAYwQ9zuB0Z1ciSPw0ApYhq
nfO7r5eHaFtv8DLxIjQaBbvidwuajoPEilLkmu4KrRNOzFWtxLxSH+nCodNkyYRamKcWyL15ipj7
itCWmgOSyissw/fMVKq9kGbxJDko+3VHozlVEVeF4wMr/oBjuTa/8HZ+svBxouqA/hZm7WvhgiNh
rCPiOFzjTKQIoUF4IzHjd+YCM6F4eyngeNMAKOIDpQTeWYyfAvZkU1zVRTueJluDpCZMi3M4cQ2H
YCq4pl2fk/LPScNk3O+Bl2F16266KcgqyN9lJjlB9pXfVk/wZ2HS4fzvXGCHI0UzwG0gdcfiVHRC
/Q9ZA1W5pdwBCTrZ2bMNUVPgv/I816tGaOgCCVFHLuXW6B9Q0O0Njry0ImVof4tsxIbGCa//Y9FI
fODOSkcu/EaKveSQwTGz/RM6nj6YvL7/MPTMLL+SEgA1Brn1LszQ90vy1LlUKtNOBhVisUVruF4K
L5Cs6ovxSpPva+YZ/jqLDEqp+Qr6+5zs6qjg7dcH4T1kkuDZdd/+kVYt4x1gV7eI7fqIhO7zsE/I
6rW0nHLYghMHTozBOIDxZxI7Gx5yNv08h+mRfeend4Y04Z0CQdqTMihHaCvHtcrmFZvHelz+A0Na
evUgXyOr3nxt4/CnU4f3zsj0KVgU8t6J2z3vHkCc1Pt/Pim4NTl4bQcZSASqq9JNGt91vg539Lyp
hOhY4xqz64gbXVzpUxpTlXB841MyS1soK5C1KTR+Eu9jQRB2DeYzv8xL0XqlP5OFoiX89rZA0bog
TUiVxl037g4BDS5qkxPyLuFQ1IXYs9B9llo79KzvW99T2rfcljRlwBSb+mPleYeQ7cuHYo3kmYg1
deAPiViveNZEtl2ASIZ8iUuz5J12CVL+EsKBIm50CtCaLpPH1OGSUy4mKl+qXb2677sE75e9uokD
CUoWZknQWJW8fHE/r0z18MmF9ZxggatHN06Ywp5mcvd+y+w+tfRiIM1nbkq2J5NxaAQpveJsmtVk
RuWF0DGmt7q84dFTZIHFUZm5HnbhVZ44jmGHoqKwFVuqkBE+9xFmGqV5S/7oWulVXA4cocPbTlaB
sx8MKLnX5WC1lxZ9+svHrwcEd2K297DUZOYVNL8VB3NTHZ6Tw7HFEJ/af/CnyYXdoapwd3Ag9v+R
7KuluevfcQTTM2YiGawp+0m/DNYQ2jriYO/5s90GFuwK+etANmL2l9ZUbkmtYx6sLvFoC0eHk8S0
6hL/V0ctlicSYeyh0xOxPSj3EC9h9kClfYA9ukxukNKYCwwXm8UrPYxUc1F8NIAe384ewPOAPIIR
NOEXW1G8wfnprrt/QVm7cP8bNztd+6ZXFneQVZVKbKb9mxZ16vaMH77qGbybO6/Cwo6W6cAfso2l
C8Nuy2Yq1TxKKNmXV5BchAlTpPtfaHSSUUZtimc42enud9rJEAdoE+36+NacTvpmxp3Pim2BhQUr
h3b4vXqOmAaudB/pC9dlwWE0mn6DLyuxvGfy4nFsvZ2SzBW99R8y/fsxrwf/750TjGM+fHcofmr4
1GnZPNB3AaAonUFkBafBhsIlDYbZxHS8Po3V8vUQ1neav2lWfOfiqLaAqq4/Q5ZtygBJUZXwqmK6
afIEW1nhsIYRiLFPJcZBOWDNUR+d+ZP8GWZkqsvEP6gffcE3+vw5hLoxBc/kykauK+lK4xd6fo64
n/5r5SwkpgWuRcMkNzkA3kxtXcPeLf/JxEtT6quVDm90rPYTW+wXReZXrIlDg5yEGwagR9djW7Iw
xjrZgFyqag5HKQHj8Fowml8f/IU8ebJIQiycRokFuuw/3wmx7Zzpnix0ElnEYmoR5vCu0ZcrnoiY
YCjvW29MUloSxhROsrCrwkqEp09h56oMpcvnicKZfIZhxmTIya+QJTtetVBbOeOM++XrBJH1Hfq1
9fFn0P0NrPwEVReNOVyx5IQ7kgDWh7rP7XmjwLM64zJ6eR/bKbdKPXQ0zSFywVaa2rK/xw+68lXA
3SwC0tMtZDRMgine4/fyUIKa2E3En+muj6Kb8ceQnw1Qdd8HLlAUArzpfu2tR/3WbEXxjFbmc0xV
vREGoxquuS2p7C9cmVWg4088stqyhWvpBxBV4wzThrsLQ3m27Z9hKUDpujs7xbf7O2RlTWSXD09G
tDou5gHBU7K3l/MJudzxE4ppAr5+MOOGYp6Z59GjMymUOuhl86mngnuqHz01P4GNDzO3QZfPkQLD
4Cjf5TSFcUs1DhHwM8USDr6KBAzgcaRtL89PCOjvoyVm/3E4DOa9Zy4oHHnHv5TYDIVMYjdEc6nv
7wsgSEJH0yH70lgwBoAIjGZwLZxnPapseB3m06a36xfjBwOPeDeQJGeuAXjhm5zMYZ5b0pKCM9NO
VWQV4SQ0UAvK3TE5l+S0Faqa3AI9VK7hLEH1XWL4i8yB7EiX7Q2BOcPgxJ7wkiqbVCMcPA2v2KzX
CQ6LZAlm91gFmJptdAL4IPuRUeFsCB8eb0prAACabY119S1At8znqPruQzHx8Mv8qsDzXYHOJ26o
wA6Lvzfv+8p8ti9ZoF9cxnw2FJcTUsmBXm3mClImIsHJ2ZQEAiTvdrjuLDQPKFApIKbCEF+tNEg0
GwkuP3sp/bFXqe7w6eIfg+3i5eGX4aYN856IrzRWuGt2WjDJC0z+geDgX/gyfv1kGqb1W/nC3gJ+
Ta0p2UuTHYkRZXejYxvC1gYRa00REtTnHsTvv6i1h7vrVA390TLP9BY1PilnK+svjOTj4ystRlOK
wYfadfyT3vmrNbdhf5AdfDgTu0sa1mLYG9iU7l/PuBqSV7bJ3FLRjWsCwCEXJcaick/WOPe3gOow
qtmfcWUSbODM2QBdY1r/9J+/bYU3ARtuVu3ZKz+X7nD5409kXJJd7udQREiWmyl8tXQ9sgm06TjC
kVML+e39UC28K/bxGTyQnBVVlRqIx0ibMo3k5nndmcQQkhrdT6+t2uAo4cfRauMw5+RAXrBFHKBX
7bzR2T7cPPlB3U+fposxQjbtuOaLbxoqO9IKKbdd84aML4d/Y6mrhNzmRiG5Bc9hMnuyc+YJq4T6
n5oSCMHcru7WNm8gJ6W6N0RrlTWTGMUHOau7C2OaGZIzouJX/1bjo4DTxlj7AlfZiKztNK1PbLJ7
48Z0wTemLUMPO2aCLNg2LYW0gzWx8PQ4cfHSnx0mA4HQmu6MEXqF+xo1gy54YP59+tmFgcuDoKZS
CuUYY5TxMA3YYIBckgFAgHyKYPvyfMSsa4acsrOniCu/V1R3aRIAydBfpCM/eaYk7TcvLSrlbPuD
IOc3SkSdYv2raWcyNjfP4NOwEAjXVg2hDijUiGTbMRT2BhlQolIem+8+nPFaNv6HGKYuJYaJynTC
66UGEKByy+5oNMxWUhW2GKgfBgRkPSQWlNJxGGAXSvwUOOdRtqvbtJ3LKnttBwSoDcjaziyAFx7a
gHdiFvP2Bd7M2/IJ9PJEUO5U1ZQoes5Hvb8+kc7wIS2KJfNlG/HhiFWxHW13j6CFDhN/M5z15bua
Sa9XPy2edeQd1Jv6nh+wYB4EUy+L2exjHp3d/oE1kfdHUvzRMzmowLAt1OgXxoDSHyj4yA8x/UAJ
AEI+L7YFQUjZGamhIH4gJWoLGGJc6MuIWIvGG0WafOg0UVuqhCqyUJmyiB1EOQOhWtHcYxPH/hxV
SjDki03jMrZ95qZjyqNn4JcvOeUytb0Nlhsy97+Ktwa8snKeZtgFfUwrPLuDTPE+JgbMQBg2wR4d
rdVD9cUc+Sf3Z6T3lAIJ2SMsKynUc6rFDJzodfB60+ccnXJ7VkyI7fFPuCWewqglLqQ8UC9MEdYD
GtYCXvNyaRY/CsA8c09ec0R1K24KFINrPb20zj4BTM7KJ6YXdP0aklVRP7RVW0bvX6D9xjLkopaZ
LxdLVK9KnznV0LUoCRzh+cb0qg1zoQ7IKDNC6TQTxTqUassImhZBQCCBtd/5GTCyf3rNMUH1p559
wq4U/sEGbl04qe8wWBsCFvJGqASHI7SFQsGjdsybSW+0V24r7/Ew/NkwJjPkenvsQuVCAmn7DVWe
n0T6XOlR5x63pvSPlcnrliXeDFXdd6O1e8hfR3zpu1QY2K/ReKWDGfEILmVRKjIcGwWzXxEaRfce
MDEu15A4S5NPUiYcdSz7EY7+aTnZ82tiS7+w9NLbuGjgsza3zJDea/caPOAEQ5ozh2ubeaYQFhxl
libP2zV5y5CdGZ9d2ZtPY+q/ukwcG0Xv11UYZywnfLD4Kp56UVaNSZbLESs0mITO0AZ3N06RBYZB
upKhFTePB+G2R0xn3F6zxhKmhnde1OXdobDZw8FbO+zHiFQ+6eoCC6+HTuQsxIt3ZMipvbGEJgkG
bro9hGwmL28kwYyCz8jimSpJyCfJLFsG28T7TiXKA2eaHU0CFBPaOaaQ0zV3F+qRZuwCCIvIGubV
GpCyV3W/u/usKXDic2wGQnrT/ryuTcm4osOWvDdarpWPAimwC/BS87HHhaf2xhbNQ8zVaFhaYw0+
1tcCpyuj2wFR0h8/p/vnHBWfJS9gCsjayV4hqS7bto40chBaTuNd4YQkCgcxrMIS9K/9EtHJ4oa3
kvL/t2TXWIf4vyk8VDt70W4l1wwq53Fkmc57ZDLb6mXxiCSK9o9SzoceAaQI9VVjtfAM9ig083z0
sc37JZXdPhaB5X603uOybv2YguQb0B8ZtlHNLTXeAScs95taE79Z7BGqlHda4sOHlUCHiO5UGkX6
V9Qx5rWKc5hqH9c0bbVrX8rXlIVDmzEwGBIqWAksUYmYbhILgecrCsJnuoUWj+TDcRDYH0Xso6Nl
xY1hfFBjcpDgPr6ZzJ5MCjev37aoYdKeazRW6U+/ZRjCt4pSsOsQRGqaXSQSao9VsJdd/cq9R+aA
8tvza3mGCyhJ9/ZYph9EuXxMofPTCntqAMRKFNICkiv40PhA6g1nYVcNwKIZHSpYMtjzGkwHX66w
cfUihdhXXMCOLM0P8DnrEZzzOHW56ymLLSFewC3tk2+8YWnLyoWLO57GyH396ZJ2yJG4/T2+/aJp
tdYVQ3kwTB+Ukhx6oDBhcaBBNPJqajLs2SDszt9BQnbVNADgTClYW723W9f6z3F8ZPgiQeOFSaFZ
SPrWm4E0I8oJca1H1624sFa218/uvk+TdtW/fZXtAUrI2HZAnR4IR6P96QCEhjoDhxC8Pxu3P6Sk
et8kFbJrdfownt9ZAyNK7F++XDlnJPPJAl3etOatVKzI2JJTeLp7zQsXMCoddX/U9WrRMWN2IOT8
HOvAauMrreMxr7/IixvSQF3hqSX4w5bqmYCjPJcJWONonZZ3Y635GGUUnbiyVvtiOXvYns//K7o6
7hKinFVcPhR9HkVZpsb/HBz96b9nm47wwtUDC11ZN9bmdF/2njoCEDLkxVtChCPmfH/a76PzqZJ0
zorYsokANvR97W4S6Z38YdvYDxQvRclEBMTSmOBXa8g5OnADTdoUgxWDr8IXQlJ8yfQHLb0pswZq
7MjlrDNZsareMqlKfRh+x1lYQH8K/YgfSWcnTu9B/FmHQNEdMhcExjkbxGuuSzyPLOJoTyXRYe6o
dqiT8wJtL5SESphKyyFBRIOJV31+i9z2XszcKMtSrmwgo75YB1yOkO/osGhUKjLFp8gBqHHtdBau
ZgoIk/yBpED2dGwwN63bgV1H9jHvp9Nec+Fk33eFVoKJdPBLy+lT0NEtJbiK7hFd054pMBMN9kBv
H6WgUj3iRoWKkQsKBLU27FP5yRYHMpqBDrQd7QLLukr+b+JHKTxEQxGkZwPe+sTh0WLEAKgaIxkI
MNJSjT89p0APH/ogXH7md+NrL4LreB/HUPGCNwL8ehZ2GibErVm0NLP6tALakj58suGm78+Jm4+o
C/LxjWuWWLnVZnKrtjLBhxnje+nrTxMXeU/FjUBUHdf6I8tWpf3E6z2NibUm7qM00QKzsHgDx5Ei
550EWf/ob+cHCymjZVdRXU5JEoSPXz0QhwdM3XQnFc3wDswU8vjpmH6rwDCKxPhzhVVlgYJ9HA4t
Nno6dYrLBVqw4eye0PaCNmgKv2f712hvNv+JSWwd8B1vk2f98TWFnDC3XvBi4pU3X1I/jRB/dU1n
Q8BRshv78rJnS2O1e1WAcAkcJae5oqxxK9w87fFlvM5fzgkXYr9MTqbpPdDoBhxxzA4p+bRMSBAB
lW5TLeUby6nIZjhFV+/7+pai+iv6mYUjX3g4LXfiWehc6uDHilIeGtpoyW2xzgoNr3IatuJIRbWI
I6OtdeQ1+vNpEmZDy5FsOcumZS1bwN7JI4rwGn5uIZT5CWtbaJmBBBUTb7+UmbEemKmF9xTdrlge
9WaVmX7bWelB4yUt0JVMb3I2PB5RdJzeAce9VFi6tnZACWawUFLYFEjBorp0XB1M9sPuCxPDyo6B
CdGYSWlhFeuBrt6T/NrfIyiivaqlzlJSM5frB3BgRpLhK0RisjurhNms0CQfdocD7AeBfhT8ElV3
k7cQgSFm9ZtRRNiXOzoiXpK0Bq5kT31S9vAbuaTxO3keeeYWo92TI/+9AgbsvVVN2dqNBv+p4utH
WF0racBjbmVHGUI11J1yoxfRw1ibNezBNd7o9vmvSBFIx1toJWUAwnfFicbo+xbaxBBAdKjZpa+d
iohET0bCPsId6EoV+lFTrbsVL/J4lClZ/cOpvwRU6MpFWNv5lybiayl+UZ4dN3ZWmYcT3qKI3kJm
s5P64k8qAFVAtD++FMSc1M8EJ1ckcNFF5Tp6uynelAN+nerqrqEJLhLJW3gzUfNhWKfVkZBp3r22
+BD96jQWB9jlmP08qRHlA9SFJMxJ13hdew1QhLKuDr7KgDMW5dNWmaWW6F2I4aBcD5wb7a8f+Dgc
xKjQM0Q5GKVUA4tHemxYR4F2V3Zy58tcTC9jcCFCo8POoLxOprev3IOK/Hf4IwTUCo8YH1JOFIbj
gJcFBKzOCjvGKOEC1ckJGEJfM4pyHZ7SUDErSS+LvVJZHy1IJzYM6hvNkVQtmOrCWs+xP9l/xY5Y
hjFyxaOrm18CEoe8Fc78K4T3Y97/vtpVZeeMMXIz7pnS6E4IB0gOXV5q5ttey4pn93GdYGR5YzpQ
JkUzBjakP8Q1JCyeIWzHXvP0YZeImz/Mh/mfitVfhn+e0oa4X/TX4BDtltnGjJSa07GI9iIIr2iT
Jo3orBhe4GiRC8kuR2U2Q0WCvaxZI0dOjB97F+jaKElYJiYaFlJmgH/pvI19l8+UtOxOie/xYOpP
5ScaZvbU9df6WJ8wGXsWzMkxZjbbpftJKQp+294Dq1IJNtHWOj7+uFscsYUyDv1IWamaM5fCC6FH
jel7OThp0NhimoG2UQaCnt2nPeAruxkMxzblWG06eQxEU3kuZSYBihFvgF/1U8ZYHnAtJt9ihUNY
IpY0ZR9aMr/bM9MPNEBmihDJ3/zIZq4gLkNYluLK35YdWGX0neFU8LlL2xNAvKMAo18m8gfQUcEx
vq92NH9YJgqhhzZxZtzj9cRdgBKkKcCwUqkq8mYRY4Hf6H+HSDD3hhdMg+ySWX1QEavuDe0TGlv9
tZb2E44HanJnJOqvB9obUCvAPEitoe5EdtryKFTKMqob3eIvg0LvPMnFGCYoJ63gN7SiCli84UzG
aH6VEtoolPAaUZv1eCutOOsKSip9Bq/b6u+weulx2ifAccgTQyb8atTmisCrUrZBCgh4tpk4sTEB
D/dD3FrVu9ymySyfbX+bImS78GYoboee/GJg7x3JtriHI3kcwjfaMhebnHyYw0KUU/sRa1rJyAxO
capWx0ZsPkrqaeFfBqbkdQVtemsa6nu9H9uzm/qzRGg547Iu3NmpXXnJC8mnReSDYrfVeV7gMJ4s
ooI+qAVohuFGSCC8htcqBZxDVcOkfUFsA7/uG+OFwJCvbhSyPYbvoLl69u+1ZWEAjpf58ywR/73A
Imz2bKUH4JZTG+iIr66muUVXfMg8FERZRz+NXb8EjrY88GV5ttlyIm4LWA++XVpHaY/uMwT2TUCS
1yeJRnHnbp6COgJ5ZZjISKqanm3C7UuWGmwBXH5ti60tlEVUM3XgUIEgDxDiXADzmbWR0vfM4kRG
TJJsgFp9M12b+aCXWcD9gCcY/4CjTgqfTmB7V9fwbt10zHdOnKnk51G4fCYeCWyJUl/22FKOhS0a
F+GiY4ryaxt8oLsfWPvu7W2t24t/MoeGfRavkDU45AItl5IXEMGskuB0TJobGN5Sby4CeZ/CQCKF
o+VPizNifh7yA+DznJ3Se2zQk5alRVfJ/HczSlYJumov9UpeLL6wI2wbed4nw4D1YDe6gN39CGES
hVojYEHuSIihJC2hIPsWX8YqtKxWx/Mxe62babaO5OVU9dsAuTDRDG8SxSc3/qubuLXnk5VORDfo
YOo9emyexS4DynUafuzdvTadTc/12umQDcqZYCYLVBuu6hJqfAOZ9sxxS2g0TlyQ3YlZTpEh3hcp
EFv7EUVciwoClbC3aK/43In1WzvTgcmsttQKwsdS5xGgiSYnZlTLPNadJAjnEEgBOGcWKsK8O/up
TetnWSYOlgc3Ov83gHTuIUMV85MpH8UOen8JqlDIksiELOyy7NfX4PqrsFqYFgT7ssCcT/ytXtyZ
ebXBaS8Bd+nVcj+GhXcFM/dxw0qPPJCjL3fIBu7WC1fb3FANgb0xEb00n+8YLvGRibbHm5G882KE
w5BJjpLhZ15qN4mnKkBRdXA3ZJRGgCmzb6+yOqYYMYgZWdmBVBHXqqojFdgrBQcgwUL8NYp5xS75
8N3CtsgLMWYSaCwdGK1fRmDjXuxPj3nYXKdWdg9bQTRtpGfK74JkoOXbQ+5Aid6lOFU82YnR9/gB
YpCRkhteJ7lncT7QJn2/njOFIMQv4k8O3hdAABj2ponBj8wDd9JaD6uRAyUVTUZ8yc6TXJFt+G+D
b7iWfLZoQc8awxumgp78ABSn3/yRGZSQtyTcX8nDKA0zo3VQynRpCJtwCjNV8Ix0EQToNuQkjahu
SBOnNlDl4UOsuH3MTBU+Id9HUMa1a3kWVUNyGWORcEST3WGcy9p53MEnx5xeR/44R0fu3geNFYNf
24mDMqejn+zLfV+xhEte1+DJbMv7DWcghbHLUsWMGtkqTWn0WnCzUvwwgJ8Ur+OEP4a4GCOkWlYS
42VXpAqwV2kESvsJDWRsOH5pfejNUY0HCjtIj/A1vi+f81AEYmgNjEIsnE4soQ6DJN60MZSD6Arj
tGBovaSMTnA1TsTgXT1sTprwEE389zkmKC0akwYFpLkCEBJm9z+Fr4pzjY9PuPbOZy6gUxjHQi+3
Q7VUvH3ZqOTueDzTPovxajva2dtqy6sUrtqZ5TrQNnC/RRtSt6tSCLc4PQBxkS0kxIhHViZ3eT6K
LTthWFMCyEEOVpm0RxmLhuXxYjZ1awZJQBhWz6XTZ/cxoxDTge2SrqAxfE71RbeG+0Ut1/e2WoHE
fKNLytgJCwmdXB/LOa5JYvQ/7RHeof+N0hdNWPo4ZNi+FD/yRGm8dQI3CNY1ENxnI9eHJo/AfE5M
fKjGvEJBSbU+9dPhWrkjwJZe9bmqbhSXdid2y01fKi4Wsq1b0THcZWRbZ/ZwB9TpYyOjZOEHglLk
f9Nr2YLUdZ9vpYPR4nO3e4aSJNT+N0mrN8CMtaqeAPwoDdhjXETB5QJhl0TkB5499EahRXeaARwk
Mi0CPXTgDNFiMnoG3otnIC/SBTbJ6sQWWCjyQf7DFnW3sCGh0hugOtY2joPdgRpRa1c8YMYo3N+m
eBs+4rni/s3ErgwGBz4SP5UUi1k5Wc6so5JaER1rpl047FUZ3vqQ946jTPzectRFsOSGWUlJgtHM
J4Gqow4VH1Eufsz0NLCDcQ8Wf85tj2OeFmZ3te3MDoo1SW6vdZwR+6G1NFHWucqr5rjCjUmSDK+l
3sNnm/lhK9A4cf2g4moZn2kuVhKmzpkJQNA44OaXcx6f/g0pLEg0ZUgY/Xy4vWmbf8qGPxo9+LqM
eINQjqKz4fkeh4EjEpY06oDgyVd1WKVjJb1YWxr85XN0NjO6j9R7IeI5fyQxore+fzzzqhYsyWTF
phAmDpSUF8VNqt6VwXiSQjKN8+QvC/p1r21ydjGIxNh0R+Ye/+EC7pZsWxl80G1W2xYPaRj2pl5M
LkKBthppp1atAk9pvHHXhdDbVgQoLqoJsjxO12FHZiSHOuzEGJacWvO1ysMkBI9Sq4TMpAfh591J
R42F/FG8lFOULl9e3jwS4vrHlYpYFQIPSVSy/Ic15ROhDd8vYyJzMssA+pOqMSKb4PyItL4Spf+z
ECgZQ7C4Lo1Ddat5lMzjNjs20lA3THsWqGG1I44MsZMa7R2zM11sBJdKUZWVt5meCfwecfHbaSfE
ZdxhDBcl1sv9/wmND5vzmuKzrz8O3NzwXNs44pRKmvkRoggg38MzNKhv3WwatFehTYLziG08FUXL
PtRkEpcWT3gG+cYZf5CT1q7LqSnXkBpsGCubf4qAY1nc74zqvdd79CLs7z1NgIFLeoDqnOkzBQc/
DECMeX/YrwIA0WvkJWLf93cl2sjTdYDA+aTfutFwahpJTnCkdiI4aYozIrLpT1qOQNLsqQ6j088C
ruSEmFinygYKa/DO4ewJRAqkieAk/aghX5l/wONYdTHhEnEKxmVXLqQmNouE37OawQ+6W0oubd9u
kY0O4juaiKUDeUfSp4VSdBAnHEdQSF9D/heQ4cX+sBqKsFk76pQ5je+QC5PbDZ3ZQ6A3CztzvvNA
4fnwOXDAgM8Z4NP/Nl/GFQSCavNwEa7n+P+PGaAFr7ZVhBnUhuCrPIeYl9m7Jsc0+G5juqjGjtsp
LmcdpVUPnJJaGf31AIFLWhsVS+itjLhwwCDEnxIuuhMr2aisc3Iij68CqcERHQLN3x2JUvjMCdmU
0AlCLNmHYGta2iwLHyLBfhlm83JhpWe3hsq7yevbo4xoC9WbHWYGn3zuUlr0VQ2IWFB7q+Zr9a9X
I7McDzgp7Ne6ZqRqKkd+58NSaUXtcwK6HQsqXyX8nmxEW6GLjPVf6ihBtCFkj4AgJ2Tqin9/PddV
nLRNiuVceMEsuMtW/3aXs/Q8DMLR829an0GL/geIulAevB7asgyS4nZCBaf1bu47noYoD9Mspp2F
qrcqRfe5LCGFuLxYK1+/+5T5ln2ibpyi2MZCaI3h8YXoWfnasPqNnBfh+ol1r7HzJ8wsJxuvn4pQ
0Q90HkC7aMrUqRuEfgfkqAQL0LvLWNKLy9NpaC5ZNVCrvfTDQb0N0vloShEnX2G4jmFbGayhvhlU
6raqzJ9qI1C5mAMQiXh1SEdPCaoLwoI9Gf+C2lrrct+LP8Zb/2by0MC/xbfK+9ioT6wO5b+Km4bZ
wwVzLeAjSLgc6O0KV3jCEVK8lqi4ixuhYFyytGZaTkEgKY2ooIFwAuXlIlY4GyZgAp2Kwssuf1V/
n7KNrq5MP57OzJmhLkdr9J1lkCM8AHufaX39vHWKqOTncdUPEPF/cH/NTyrOEaboz8C6RCcueO2J
FixLlLh9q77R+Q1eRDXJCPb9BpEtzJuU2zJNtqNVWunh8n+o0B329BLRGDNJ+6I8XCjn83GNY5k5
8PlwHPZ09CT4LV2zvIKOsYv6/3O+8kr167ED4Td+NwfOc+npreBPNC4zQJKf0ygjAu/9W/MqOtv5
3N14pRzqraEOShnkVGxF6oBCfsIunISOK7g3THErlSHeUJWb8go07Z/CxXjrJxW6egl6iczUzLfF
FfVuavlwXGnMQ7UOo9S178ZSVz1LqFhywfAOvSBG4A8UQPQc3Daabl6dB4yAF583d8FeWG/ThScR
aMQScBhgnRokESLJLEJY7K7U61yuS8kNUF+lr+gRwxirR1iiYrfiAEKRt4kcGHJNQ6uLeTLJpYX3
xri6FURMF/erUbmHIsDAYn7gpC16L36ER6zAtKau5ROvxcWbDuhsAjWGmCD7GJ9S0LwHDDqQ0iuH
tFSJEPsCs7uIZpvQx5z/+Bq9hnOszIQAI7UKia5Bfo+LuARE7ONKlI5edsgNBxxn8CVd8G2RfKpo
7G+sTC3HbmZFjmUEP+aBfWmSTMwGOl8JtroH0ChClo5j0cCIw4k8SNSzAlTF1ozdktXymRBZ7nNs
3IBMpPFP5ahbjkvUsKCiJzX75N2MqvUE1XgVLPMYWWXMlC46C8n6B2vA6WKXMyXBFNd9HmEJEq8J
OT9wKKGeQIv/uUU8aIQuQ6XyZSPU4TI3QryTsYYFewsR/KFnaM41cb6M8XeL20DKYY0j2Qqs5ZJx
Pw0RaDLNnpslmX5xeichW/tPxhO3Q0GWo/lYgJw3itRB+Sv+kZkBvVvzdWwnCnNFzgAbphQLUaR8
gENgUgSHSKaUsn2fbAsLZGihnBvUr8nfyq+leyiqnlv8FwF0G11lq7Dh05CsxffgBGQvfNpl8zpU
i2H2NapbBp2oc9gjAZ4I6mRAJVoVsuoPkHfGPy4oy8QVywWCt0NCgyqlJ8sWwBQ67AM0nzWG2pbl
Cx+ZJzCx8jDCCjz696fvFJOsMU8ToxLs5U6z70rdxaU49ZarnP1HsnqQrUcbty1l2AqMzemDglr1
E5OuNb6gziXLx2AM/q+OlqmZIeYyBIxADhu/CmXlQ8cLpfYY56EK7gKjercY8JY1o6VMq1IlfFMR
O+xjujWUh23N3H2AoZurY/NDwlNnD7Kpuetzlx43Ka1EYO87us1OjQBydEcNKbH+IH3t56LmM9tc
f1u2FKaEdZJTjvL0akf8xIhAKKvichZKWE07wt59og0MMMFMd43MYqy/l97YoYcTl890cx6G4ZS8
ADVEvbln0oO+FoZaASbmLsOE3KpuXILL8ew2zheDxvwhhc6YQkLkrmBzL3LN72PFY/AI6S3pTq8/
iUr4k88ZjJROfSP6NnvSB9jYuvu7XzhixSwNeZHUKdxSJ6CfmyS6ive5omdk+g51MfpQjs4B6GM7
jANy+O/JapywuzlxMVSX0S1LU2ZcMhhQEEVbd4HT1HSNfhbKgRTBD69C0VtIRAq4+4eqRPdKMAF1
t2sfuMDi2Ts3U4y5e/imDheUEuGb7Zm95MoR7k/5QzF2lljRBfYLLsn8gBVgaZWY0V7tRIltYw1C
yhSeAeUgedn0xAEZa7yK6waDhMgRhebPBEwuJj5zHvbG6P38bNoy1QO6YYh6NUPRYaGxrd73yhaZ
GnETe7SmpLREzo/tTsdz/E8IOuvrZBzBWnnZzsyEwUeYSSYFu8DiIU2o5hrOgVhqN030ld7pO0MV
mlR9ycSNv22figk9HWX5GQo2lBva0Ui5uU5DYMZM/7pIGJxry5X5pkBD5SCgNLnXIl2upspYCkdK
y80XQ6Zj4G8YtmkHFA5cDQ89+XH5PJrhdZBYGzoGF6huOtz/NM5oZop8Y8rTwUtVJCIDrnMRK/Wa
Wu8NM4LQ6YTSJsLsjSQc2yf685Zb9Pg/wACmN71i6KDAN6aBX/EPbWxLsBRZcmmIr1iVzi2ozY6l
xRes1WqFl46N0bbWbl56p+TIcMU0s/qfQxnAACG040xhmVhiIBIkfmVQgxkQQR0ddF/vB2Ncu1gB
nRsOhIx0jVim8zmqSzigEU23fSsnISwjf6o15jhUCW7QFFlTnF0I3M6RuOO9dQX1H++m+YDm6VXx
y94gBtJjddU/p3C8Jv4RtOsnScPN3zTxcVR4HFbBQzIuLfLwkAFW0HOqGbXW3DhnaAIN9bbqSODZ
+T8T1FBNjOiIDHZEH4BuUJp6N64m5CUsk9tUy33B1BFwV+MHdIQ6IMJ5cDYIiSathgnc5DCJLkGG
nFEP8BvjQYIk5dbhoIZF2RDWN5AHzEqa9E8Z4W97w+d+XDACmMKc2RlPCASgOgFSIFgUhAdhdEmV
54F5LRT5W8Du0o9WpXmvvaS2Ypi86T39p6Q9C6hMMNEjj5KiZioxinMI0byO1IRWevaPXIAYNlmW
Bkn20sCYMu4rOMz7ZlEc7SxL5ADSGDjGI+zm/TjzzSDxavZWpD/gKljRF2TV8BcWW9Cg+9j81frv
8+/pUw1Si5wBPib2xigHZh4BHK2Ge82oO26LkLacLGtOO23NUdkNijB8oZNGVdK1L0o6u1y0R4Yf
kkNMKhmuSRrJbWG3sofz4OkPl2qpbtwK/R6v7ObePvI+5dIRwd0fFe52UEEhoEpkNel/w3wXBe+G
KtszFFESR5ew2zuM+5QCz+5J+6lrygz6GJ/gGGxZlq1BS4OTqRNNU42p1/x9jOFLruczl2myYbrU
A/IcutfrYWnPB6FR/VgRXZCzj8WmCZMKWmH3uQeg1eajHkvTcJdMRwfKntx3UWz0ugVhA7mM3yC4
u31SMaHYLZ3RE0y20gwJOCroj32g9t7qcaVEhlmIvz8TdJKueVGD48Qlc/zZQJj1P1G/14Z7ZNRN
q2evbjHp2JH3cZq7iwRYpoGZiKWelezcKLaOI7VVyf96CpqCqtvspLIqyPwUQw8pB19oCiqN+pSN
dWYIf50hqawrYKlmMkhECq+bio9KzfVtn5tjavs/5+jecQ9xP+e7Z2/Wk4EACRbHnvyG9OwYLaAU
cLEOhQUX0hN/2SbWbI2RvYK20w77t7HxdzLjl57Cft0MPgRk5AAtlmpqbnbWVfQYWHNF45TnORaq
EW17Q4zi7cMwKSXAjHtI9+/G9OnriHEnlYj/PtGi/elUHD6DKcblSs/Sc1hSGXDcDQ2CYowzN0BG
cthYabUHdBat4dXM6RbsZjcgZwAk/MyDsecFnv7xjZeFM2cM2TxZzQz1JnoN7bFaLRl3WZZM98e2
EryGAwJUta1TKWx2KZjt7kIbs7OCq04gBKOaxVpxjJqpbfdlXD+OwG87jsMry4do3vR3hHYA/3Ww
/GNdqC3hpKedPxxMJMaqhNDa/BNIyAidIaTQHpSQj0qsqO0Yy4dIM+Ju48C+JfWUswmUoGDdV+Qr
Aa9AhvIgdQTaEmY0thkAQYRKWWLtKsYKW4JUUnA/lFsyx27UpBpaWp5gjxwq8+6e+E8pdbfyMegi
39L/9i0XvT2UtdESTgJHYfJaLUESozKfpuO2JuCl3EmnIdX9n6ALA1Lfe6dk4Z/uMOdIqmbvCW1G
UQDdoq7zX/MdlHBOJV6m4z3BN3mEcOltfoG33viQfVFuHEw1VhjAv9DB2XaVJU3vNYX40bvwumDk
DEUbrpoXX+LopY5rOnP3oMBRdKTiTSewC7smI+zvA5FLoS6YtjPamnzgAb8hcy3cTDvOG+1yIO3H
WqRuqbJVC2Oif/mDq8t6UWmqUEW+eUfAK4XKiOZsNfyTqDVYZ4LLwM5QhkwY68zc1OeLQE5hBHkE
fMEqByG3NoGhc0/uvoRtJynTnBFaH2kkeXPZT85K8flNcZ0Pjk+210onSbp+CHWOPHLreoowGYYW
TDdPt/0NCz+6r0PPkMaLwM94lArWuxcNRgP5TMtpLo4Ldxt58H3O4ldgcLH5mqCe/VkZYQLn4y/4
fgJmZcq7q77PiL8doz5yKHG5xQ7qzc8lxGvQ//viIvb3UyA85hDC12xTeSZaQL/DdmMIaYiko+hA
8tMm1NMrDmeDkxXewZA6V+dYBC3EQUYUmJNli1RpTV8f0ZK49g/jFZ/PV7N8gws40YjjGjwFXDob
4cNvvt8hAafvI2ZqNjD3zGFkLwyw/n2X6S2gbyL3479jMenAHJTYkpo+ZZfJSh5pYOZig9jlM+nY
i+j3EizxHDGqZMdhx69hnPziBs2E6T0mpVHLQ49HQleLbRlsVD1mTzPd1dcwCwrFlfS4L1Gac2sn
mr6JZsT8lVLaH/H1gJ6pCfUwreswcxzwUvK1K4qRoio5f8b54NWmGR1V2eYtAkcTnlooT1atqSfn
o+GPfdwcw0gsqoEsG8Pt4RPZQCXngbkYC/TH5bWZAsPYRGLoStEV+il4oYvn7LKjoZEBOtu6qcvU
tcQH+iGYP48hpzBtrQlFLgN75oqPQBrdroVFqKlQmTg88qMFfiy2tj9aM5sJrjj5oGQjoSU3JioV
ZfdWArcZZ/p6gjK8zADAXobSYPSYznCaAkxH4UbhzZnlQJO78CSwK23e1L9GX7DNz80ppqFbEbfZ
OWz4CPHOgleGUmim1y6oPBnAuT+AAq98CFzWXjLxojf2N8Dv3NPDMceDgIFPDXLnzub5ja0ddpCo
XLcAQh2B+iNPPicZ7dXfGdIIqNBomkB7NOeqyBR6yGy2JLAt+AXelu+3O5DD1gxh90o7mOqj1dBU
nLtQXyBSV9wB0cWYRmqW0eK+RRV0IV/uDzmp5twt/xEcVX0l+RBvyqLxSnwtmBO1mIYDDh1ih1UM
+2hwM2aRq5zdAwdgqG0aJc6wSuuqL+eA62uO3EbpIkQVWr8X9UQ/l2KqHamOn/bRfXTPb6/TYZiA
gPQWrN/eja6NMyexk3CJbCzjLl8z73ZlBhBAt/I7kuQoAskLP57pIztO9XeutA2aT9prWUDk/SnG
SK23eCJdBD0gkhT219ieX8tiwFvyIVl3+0ashrJF2E/voaWAo5DNXx5ls2NQaGEqB/OmwgJsqGxP
q3FVSWkyOYHylwNWatJLWRkvk9MfJsvjwFBOpq4triE4t58+LgnyaYMSf0bOY3aN0G+wVBbyVTPk
NlAiywrfMdFHBGztVksfwpJzm2QrW769vzYY15ZJcskYSrcrZ1iOem7vItvocpRG3zSnLgyyB+ZR
0wvUSFzPWEYzwgIDb18IuMSuvpFeZ0H63WEv0jniSnl2hMBDVll6Qo2UVNzBc9zh9Y5s8nTgMx3K
kFBvpteZUrzZf+hGp6ZiKeEjpz6USsYjLaQsjdzGJChx1CKnnlFiefA+WeGDFef/j1dnCzllfjdy
qpb8luqfYaZSjq9StngASg5b/B2bI0gK1xRUAl1hC1/toXkRj7et0t8m7V72in0oTULT2XGGZeG0
84RL/xRhTk9q09qa7o1wuDUjcMrAxhXjYgx0OHBGJE7xFmZlzUapaDqj5bzh4luxg+GTkVJOlrA1
wN5vKgIIsdEf5tAWdlQBFvxgJTY0wn9ID4xApAHQimwUSdXMd28dqGinbNiRRs4++PR1ixBYExky
s4npw8UXROVtUd0QVdo+vXu5z1dWsuWu5tuH4WpWNxYbFTTvj0Jst6dD0iueb+JWsYTWtLcXV9lt
SZF6ctKMGhx1rKfVor/AdeACVMtfEgic44ugYBwr9vVy8JXYYKhz9f1YpUS1YtCcxgMT1pLi8xDV
icrP6WkMCVMIs74m0bZDh0iqvyJAQJNlN8lTZ6IT1+Fw06Ry9sAXCVkkwQsiacZIFVXCfMnQEGFd
2ve55i/L+BlgJFoBOz5OlSlKbOz1Vg7wAnaarmlgpOmqPrrFGZV0JxTLVMQ+91A/EivJWKLaawT+
gpE4KxxY6ly072ts4GPdP/Ea+WfDynMcxCXhPk6MI9c84qkb2KCfEXlYMlQzNwzjC1mAEV8s3El9
DTQw8AWnNwhLVwFPDIpNe22MSsMfppaHy9Ng5Jf9AJx32sCklxtHXcXf6cDyrd+stAVFQtE0nnPN
dp/B5OGOjv/DF4B1GMn3krg6g8Hrl9W3WoUoTgMq4p69MIpUQJhvLRRLnkPOhdc0bf8oob5NlU7K
ARh91O5gueKVeRQJr97htyf0ES5jMbsZtRuxBQnzDr0Ub4L73UKtMu7OuzUP9Sl9Wy32B/wbXeuV
LuuVptOdxHv1Kfl3KbS3c1j+hhEQjivovOs5QQ79eT7MnQaEW8gbRnHcPBA9DOmgbX6VLkazIKI9
g4rWYj09rdlAhd4+oTK2TMAWsx/GPywVyZ5388CgfcgiHpHEDslE4cZ+eeh0YbwCQ+6MSlVhRr4c
bB14okYpSpsJgGQMaeYs9pemhz/DSAKSXNGcGmt0OmOO5U2a8ISBSidLXay3czZSuBimYyGhiHxo
2pvDvBD9XKFu2djgpN+rqdr19CjKf/C402Dp28KAoRNSj2lEao7CIvBw2JwG8fak8jjikcmAYDzw
nDA3rLIIsf+8qNps+oV5sJhTig6iONWL7XSpmSYVNNnPuwSbpjOjPDHGWTOLCNLwGded+rdiUMtH
faZCovKhSHgjRq2DF4sTwQ8nAoUJ2ymCNiBrJo9l84WtUTKWpQu+xdejAIAEQVfpY9vYYNCGdQyn
FuynZYAOJg4Q3tcIwlfVcF6pSmkLb+V9bKz1xO3ZN0uSfKhHvH1DX+f73PbXzyJUyucWPjCaZAc1
8l9xyPxc42N8k+xvMpA/TGrD9vOC01mhlasDZeOgQ1lo6KzF6xYVquJ2jqvK8sMU/S+BW6c/NE+r
7L+o+6ojsorXrj9k/0xHFzCObIEDlsq9z21wQEEmQI+4XCKKi09eE2z64yorhQygCqXkmttLLsUC
OeoVkG4GMdJvmUHJp5aPrXIOhtWTce6g4RFwQMN8n8I9cmcFcbU6IJJZOnoErwOER8gPwoztSI+k
lEh4U6T0rBKRmpX4mMy6OzScnKuWvY2NAH3W//mA8zoJfdizXjlBrECFel/Qu60yszAqhfHISYeN
5eew0NY31PVfP8KENlBO5bboEUYEcudBT2UuCMytcR/J61VjVnDI4pCIe1Y7+wXKE9O2x5JnYS6P
Z8FEX3WSWAWJlNitNkvq3MziHF8ZJPWK27pu745wI7qWNkFzh8RmS0SOmfplDaLYgtNrPk3AFtDI
g8DJxVXHM+BfwvQLi9v0tFxS7YBh81JOCtD3LEiUIrCpvGaZTnLnsh8Q9VYmCTnKaTxNct1v/fgr
kyWzC3M7a48Znlmv9qjIbscEivL0ru1POMzo8QcWlria/8eo0DCgHATb7cKUiiTzGVa1UrjJ2IkD
KoxTSHq3e0QpdHOt1FFE1klMGPQfzJqx/i5V+CS1rfQZfIV8Mg0lkTTbDZHmka298oyXHogA/RGf
IARFwqGvjUXfP37B/cLR7qgESGMb+4beC9zSkbee0E6En0KdWw+XcTexlyxJFuPNBHqGKJBEphqD
U5P60wE5OYfPaML1pVaJI+0MJopVLR9gVBK7UJHs3RYPc/wi3dOQ8yfYDhuvEo5alWLiH0Ev21uH
zv01PBdM4YW9dHpCjUbOcRWPu3dRnKOTX1qq+NCdL+SbyOKmxIvutRGyc0MytntBYlmp49h4TrXK
nbdUnR4Tr2R0zEac7YSPpS2i9qpDC5BMpL0K9JSW+chg37xPPqtTXrm/KeFu+t2Q7luqqLiM3ZhO
ZLkU24iLBvx9PcJypAE7VxGCiJZ17Y7GglGQDdHVdqiEkvQNAH+OVD+/0gbHNqbAd3v0fYeiRbqk
mt6jaPuHStbslZVjpFzKwmQw+L30sUtJplBQg5G1QKoCXD0fXLYFcMR/fF3BS16eelks2k8Vkdul
QujOx3rKLxZX6zKAj7IzRxN6/lqpLsp+k3W2Vdc0bdKSAc+Cdb0jAXRM5zLvLr3bgqFScJGIRxc/
CujtgmQXFTaOVIPft9BrUYRqb2UrCyahKhOoy59QHNkBGVzhj6+nppEzedj590Q0xFHp8wB2Wx+M
DKQQF1Xs+hNL3jV09Ssa1cuiykZh9I/dyv+0mYx61q40c+1r4fKDQHC95abIkPYo/aGlwbTSNU8G
5slseRYSeKQxDSFiDyq3jzmtT8IdJP09GPGk6bKq8rNyy1rTXuSe6H9VqGnO8ridz64c/GIoilIa
R2FFrf+1LivkFo4xta7+R7AjQcYOKMsZgMXCf7POGeoTqqfeShf3diCM3Jd0H3qiTGHsmpSgbPbB
X+0m3UQk/582OtH1JeVluS2eJCzdHZQISeFB3Qnkk/xBZk0k1oWA9kjQJKXijtjORDhY+nxw1BtH
5r5DMEQn/aM5lG0Rfe1nZaDEkf0Ohn3wfWf3ikzrHKN5BAIxs5GM6yC7lU7O2yGBBkNfegLsFTlv
LlgCj3+3BR0Q01WqJ3uj7Ulxe3RwEhsi9kXjRQQ/ww0qv2JAG6daR4FTcn6dNcOSmTOyI2v/tHbF
IC9bMtQ3yT/hmbMn2QPahs8ub7/9H3ObLRbxpuz3PWFZTM4qj8raT/5jCUyM7Y1hxL9BZY4mykQR
vfZXAUscFWjR965/2Jxj1x8q2DR99/kV7JY+N9KNAon360/0g40MqFqd6a1sRB4akx33/b7L5c1+
FaBlvY4zLNK0qfmt+Yho/KUbz3N2vVR+fFXOTSvy9IyVyrsa0/QgL8jhM7K7KeyTelywfMkkHxcd
EqSlld9eH0SBR+vhFmd63beNSvMEcYWilxTnEs7bAleiEAxtdv6TIgvhurNaNeyPraL2/l4JzT/J
CV+jYy4w4vfCjyQoLRteKQZTvireaXOCopRdW2yapGyyEd1RetRZYHHIEpHbz9t6DAW06HVMhHCz
j+tW5erPiYVenmltggJg48FhBI9n8y6tqZU1e+38bR0f/QBn/Mb77484ucQtsAQ/BmPtn8vU/6lu
nuLx97U4TveXXO0qrP51DvgKuyOxRcq0XRIT9/ijgBzDlvMKWl6w6G5DdF1PSI68DIjdUFyc/hbP
pBrGu6vjnljq28Mmd6bqQHAaO7I0n23GJO5eoU9YoPjmjeWghQSbe1y6QcIcJw9c8NofvmsVNz6F
wmsc6EnKo5c9mXBNDhXFGLMl/VDzhiwhyW49mN+jjHJzrCzgqs6xOTy+KwXll3L9czTbHqMEZZmS
Idb95x32qAiKSiyFkscSGwGhzXRNE+yNAaQ6SHWr3Jn5kic9J/0EYnd2Q41x1mOcy3/CH0ojwysY
EmwcIXQwDXXHko6bTKab4y9phQDzvSGggYAEGIM8/a9eV74mfc/lbVm/Dm0AWwcwJrd6WJSv//f8
0QHNU5T5VzUma/yMNVBs/mkes594qm+gRq5T6FpE/OqYb1S3pbREtqHMztE0ZAXb3Sw8IiYgFZpA
aE9YmlpHa7B6c5/wlVfTIz0aDZMB2rXmqVMkjDEaWEWt7D4DPkmeyF+TdcaosSIXaDZT+PUYVnA/
k2XqBOK4MJFJbaO/oqi3HhV5IIOtL88WV6PwE6RxIBjdHnvV/wqyl5cTW/qfLdv5HhOo303j+e4t
zi77Dq33zn6avGzMI94XDEi7Vo/SrQr46lr+bGu+u+FFKvdFp579M9hMxDJD51xIRM3vPWn1lG9c
TxfcMX5JOpzYe+XXwIjyX66z5AM56TjATTHsrx32YwxFMr3g85uwoO7kl7uKXaKGxgElnDxYgFYQ
EgGyo8zDiduNZIPS+f96nLfgBWOrD752vTqn/zpiizmfQ9I5AnU9CjzRuqbs0+q0rF3n5uzjNC/g
JQorI1AnqSXIzeXTsNtYLlWudyxhI/KZKIjn6LKRhrbPZcEtf2o8U5KCony8AjBM9yvcYlbF46g3
dghvpi6qYDsFVFL9wbIlrGDzu56C1NfAa39idbvMr4CO6E8EIFf2F3z2QM+ozZJS2BbUkPhOciM3
xHhueg8xNRu3KS/AC12FsSFjMsn3o9t3pQH/jPMfZIPJ171jbTxpDv9wwhcT3TWgl8NIEBD5StUu
p0beBeSUIyuGrvU42v39tpZvB8b61QiecXZokYjmbWGLMQXJawcilr3RdIZ1IWPN4t4s680ZXmjI
MOxa6XlQKnRLLSkohL8S3Yo0km9xHQoqxQodKt6RysA4BA/BkgRrSa0gKEfipeM84bo2OY01wetb
2eMibxuiJFGDGtwgs0dn3gBPZejM97+3SHNrlAdu2/5A5pVcww/WNyw+5ajKD8RcAEMXJI/RBNVB
F1XBFYtdj8CAXPYPy4LEujbOwZVuoMSEmJRmMzR8rQ7zDBfZh8MBOeaR9uUztR48/pKGWmybJRGJ
lM3xFRtIm5RG8X8uBBrQWd8+yxSO7v/o19Fa0WLKSpy8/K6P83Ih29VWL+QVriE6ff5L3FW8Oh2g
yOpzmPC35Hc+Vg3aQFMRidEtyzxBgCDblL6SJtawD+oquyMisuHNZ7ckRQgfxTK0UbCwdXXi7oUr
nwpXW08YbM4ikt8TKx/Y8NTY5O4euqYfGnZ5ENpLgyKQ1v6U5ISWp2p0yZNg9AZbctgQ7C2iJ2IH
Q4V8YKPrsXlLtmdsXfWiagYa6FqA6ULD0t0RNejqo1ZcOXmTSYjbFogYvop0jyAL+lGHdmxVLboO
FR7Pt/8gmHhYLeBhEz1jMefEbFprygVPegArY1/EdEgJxCL2shuob2wdij2IZ55XYyUDlSg03lYa
sTBBHXO2bHaVzIhFfoayfh9u3dqV8mne640aRlgZLPhYCuXs4yLhWc2+ISDRtQRVQHP6mSG9nOT3
6WCtcay/OoXFPJNmZWCo23iHJRTTqBmxUrM5yRoFn4LzheI6takA/u5te1uI8K6e54ZcPNQBH5ye
f0iJ3y+UE6zBBxXOnZ6JP/+I0RLDtx+83I2ZO2VEhsZOdz/OPwtTnD4FkzqVkaabPDTsQxSD+A5I
yICe6nIr9WHsLn8Ytt8T/lj7jnPEhiCkJM+VGXvoGs8i7VirhxRBnOZbVtZA55CBTaCSLiiG/rM7
POtDG+aXoLHggpZuJPGpvBfEXSLOjQerTHALSbKzDnaY39gGPq4J+oO3tJvoHATee48xwQTnyHVF
aMnQKBi8LiY8HrQ4i3RH9S7z5KFZPVTjEs33xlNosiHizQyKxK2Hq3Lyr7fmDMV0hytTDPndP296
CRIeHTcwnfgcOnIPRUpwSHermQ0QUex6BMe2wpstWdboB0C9hJLeTLlKtHNdr5XxYKPym1Bu7HQd
17DHNGBMCqc46A37Uzi+sa0JhH9eqGy47zp8b5/XFnxHQ4OGEQOdK6pnlMFPu7DffKBsa2v4c6zX
tu60yfZ1p0ky0IxhHSW752Ev2QcR2RDGDSeUuDcnwHnR9XZTyGwd0dhH0IWxo0mHr8G1kE/dnEWB
oC7W0ozx+zVGJys4fWNttXgF7B0rWtrCeVkuLxIsK0xTEGZNbnsz+c2ID62iXIn1pWtuBYnEjGSd
uu1AqEaR3UKTEBQ1/P4eOda1p1T8YKO9bLcjIXORGpqB3ACptJavPF69nb2dC8fr5XiywT1hvA1b
h6d+/600y903UJwTxehO2YiLNN2wXIKimFc4Jqdqpx1QNHSj1VBE9MLLSZH511FII/vNG3G410rW
tSQy8Xqorl/JvvwRFgFK4xdSazKoo814Jg8wVbIeqamMQheWFCHKY16cHdsv9licrdA4hC9a55c5
udD1cMiON0DuMarQgEByLe6wTq6F5+uDD7okdqeSYcKnrdOfERAm6UqhNLhV2ScZP+eUMfEElVju
lDLHogLPTKpo6ijhQjW9dKDL9ixhmw4HpoJ0LgnKL1nxCamZfyl2BgU95CNojdhZKF7u7uDrZRD1
ag6Aq3xJFWM+wmXn66L0uSAWVafOL1FHXolXel5qFZPQUXhbrC9cEg01ZLQ54tbxCWkqS28obYU/
OmCUKe+ksjO0/16GqJUx9xaYM8xG7HKRAoJsPysztJmKvFWcWYfYcxVPLRqxyc/Aixzec2KO8aeK
x9EBEq9vVnNNCEadjBI3mv9haRJdCrOVQ+0Va8M/1Pgfnzkbc97nrtW6uJre1KACW0wT5uO46a7+
GucXxPPWOf/+yL2fT+q+nW0TTFKNiPru2jKvAo8in3RFl1xRzwYt5IuPPRIe/Rp/Y3DUHyGLrZ3V
Hifhu0c+RAO93Zf2nuDEQXm6PqArg4mLxMD6Vp0xl+FJ9mqDRN34f6awqrSuY5o87O9qQzsTkHDA
NpnDnAy1lTG5nvecc//RRjjza9o7omo/vHnMKxC/V1+bfJQ5Xvjrrw93okYlRFqv9jQZ5CeXJgCM
eBLHCBDvzXNI3JK11PjxGy9s+QIOtePXMscJgDANhcoP9pX3slzMIAB/BvPY62cuE3WphvYMwqoo
2uIrglKx7M8ig0h9TH5wbZstrDtZqwgy/BTJa96UH54AjjJIAQlsRGDd500fIWUm6sAz9slU/HzT
ioqgSrw47PWa4ok0fby8qgv317Jk5zR05UPXh9nE1MIvlx73j4frBVbL272e/Cp7sfE00ebvk1zW
PKggRXkz/vVWH2K6EEF2jWk1D409I7jnyoFeY78rTSlvyIQ3UheK+ZNvuDj49y9pPb7t/AdEG7o+
vk3BD6Yyg2XHHa4APJpRQUfK/ojkr0gZ70USDEwRFZeh792F9+03wD4pCkx+AlIS7mXM8C4uOopf
vwCMuGj9jD93iVretm9gZpWuJCewTFXECsOjXNScYwhNkkMOKaYKqQjsSNsoCmGS1Ov/FeFWZFIf
a7i3HXUXFGc/QLpCM1zFGuTMF3vPFKwGnIgbj/H3Mv7BXjv384eSOevs8/DKGSNzFNHcGVpJ5yPx
gwOg3lfxl4nNiRBx6qCrLz1TCd8BC3H4CIXEzIsvDgmrMj5T7HtOeHiatsI893LDnTcWtbiJ841H
ISj01D8ZSm44GXGK2MmLX1nSB0epme7CKHiRjPpU+W2lgexbPTmm2FaVT0GNhZFo8ablsytLcVGA
yxRh48Xm29azR4T4UnhyLA5Gce1h45TaaL+0H22lvSKMNt7P/jk581vfBJjBB2mAvREfOyXuXrVF
bdMdF0TlX1E3PEwEO5NOgEMNUzLO2hdIxNhHg18jZ0v/XKfZ3hMbU1R/E0jnZ8yyIlnpeoOyF8Jb
IlCbERsVooeHoXVet8oG6YhsZM9jnXO+VO72Gckg/9B39oO2d2FNZ5Nqdgdg9ffTRnOz8/7wSWG8
AB6Q+Jph8lk0xoEiwzF5L42byYM3i7DRGHps8z0S1kx1A24q2uXDgDxyoJF6MdB663iirLqs1otO
4VO/kofAbroubYXdASyNfbxFOVAiRzyH0HMWIgAJbCfQbqA9WzerAxvAfYnDfyJVyel46INn7vLw
N0SutuE14zyjoaI76uCQdagY5AXn2CdIGw2PRkdjzrhcmrftt5Hy9EOP/Ht54BBw5b8UFfmOxqVV
TTsIUkCUwoU4V6LVjUuLYRyhSaAhbPwhJhAw2T+GIHoYjA9ozEI/TW+CmWvad0TNfdOS2iuinP25
8j3qWsibBHqVWqCYaAQhrTQPwlNTuhhkFeLbtyVNLhQ7yeSOiNFIE4aX25Gk44CEHObOv4/XLoRU
3IS6R/6ZJIxagHzJGloPyxvM5xDfw1djG4ny7T67IXmayTGkM07gKzfXz3tfilJqApkExVxT0JHV
o1SQsfYyUs9Vs3b/wq1k1hoDQEgT7NEa6AX1DwUk9i5uyAg0gh9NaL1Q43SDnTaDxUZeOS90fbR/
8X91aDuM7vFzuJK++NvbUWOnfCr4qtdA2PFtKv/4pkKs9PsVvuY0GiI/lxsyAQHQipYbWcpACmwG
SJ731e7xcuvsi5SEluHt8AWk8QnpX0vpIruRKc5y745n3ML9D4mXu7PtN/NJt4gcpGay4EOCtZq7
aT9BCfXmesfFg7zqkfU8xQxggGrUjE7z6cIuhR9zvD1/7jDzgk1UAwkxifjH3yyAQiraav3FHnTY
2bdnRKXND76B1wyxyjU/VzmTOtgMY19bSVrIbvu24TafD+mpUi11UAijH9DpVIVTmBFxLvIpLHj+
igNLu8k8nwT+jPZTwPlif4gMNidhW/emntUyFRaEXEX0TDHdHbXViDQy/1k8SxtK98V6mQ1a5FZ9
As2zH+YF9GOkIip0CqH9/thBkRauMyeacenDBN9S9pJk6CIxolo1FjrhsAMIjvAjX+WNnCt9abhN
xl21LtjLus3I9MEcKnLNpD5gmNIhYe+nIKjag6xftfmg2uCu5GbCcKtullWmOJr1q6xO+I7btFfY
y+tePqRX+zOMl1RqIGkoNUgk4CuD7bPg5KmmyA392C4m9jmbSu5sddKwzfLFAQjmFnXVF59rzOby
lvUPnsLkF8ddYVFdxYWHByIe53qSHWfkYPKGVCWx78hfLzRtBdI6/JlEYcJSZeCAv/aXA0uXk8Fh
WTdql1Yt8Uay/BOh7r7Ej7HBNOELnpS4GqAlUTEI37iAnsWZxhZ4obPG9ZuCCneQ8WHXpZfJLs2J
wahe23HiLiQ5rrqXE3ixV7gsd5aoLDz0V//A/cWb0FVqILg8XLBIK8YQJgzAyYjx6DXzGs3wLvMP
JXXQ2NLMhQ33xZ98kMy2bfAGmUWMssMoaxs6YMl5pDb2GkRET1unTG0DDATZLHEUXa09qUoumQcz
WVvo+AGtTRmXjLa9ugwDHBKs7/XOfPCrVUAVAhbvJsIhwLMo+mEE783JzbTJDHHrRqjRVa2ezwlF
qvzWcMfe//9j/6p2iBfaIeW0+9CY7/SqTuUMZNqycWcVb44FnuZoYR9eB+izbNmHv4ZOGwtP3uy0
o+RjmUOgq0qJJSuVsMj4iirlgnW2LbpUr9hVjUyrAwohqrV4ULetVyWQNvKNyziaLbZXfBMn6D1M
J0hrlOc+ZUEjjn7Jmu5YOQ2PbNoY78IZgh8WVnR/UsnVOySxeVo5PU+tovWVfgNxFPT5wesH+Xyt
t1oGBdQ9smYYuK3qsD7R2li12/nQf2qszhuGRgJ52bolVkc/q1VzFYby1LD6MHclYRR8ZCRYUn1W
9HrUieYdiMb4Mb2BgfkkHBl7Y/4owNuokd2WeidJ9fwXM4I8KqnWo6dHUwFeEO6UhaKhrCnSz5YK
GdyCGGgCOr8s9YKpjTABQpXKFoeapER3QhsKuoSlGkmC1ze+z3RQMf+Ml/jeO4lmMioqOk5y062o
FMZ4z3XE3rpW8rO3ptkIVhBs4uv/Od1pe3TI2ScOn6v5Qfz1voc8K4TR7iGnyTJ1cHiS9SF+xJpM
drLzDzxrYEptjbFsjtjuzg2cO4NsWeSfi3vvnonOoWUtob8T+OcTdY3pkbh+ajsEvebydPY2SYEx
Mqun2Yz5gzGwEDbnPl0EKlAdfHfvAV1UZ1wjOceA5jm0XDbJ5WldO1m1+azi/4u5hXZrs4KYI0Kj
tHRc+YfcpZgxMqeFWxwTBFbVxK0nI3snx7yLXsIDAUjMkOPnP295anBTXcdrBYRHd7hgz3s/8PUT
lMEdXQkZodotY7gJLVL1Al3sCYNXf72MPxo0PbR9ngiy0IkkeuljyHeecOdRektCWUgxSplj7mwZ
lqsPWeV08ZNF81W5Q2MsQK+qRsVjpp8Pb7y8EAAAp8It/w3Rlb+ySbpuuO1f29MT7KOABZpRu1Sb
ukenkWRvEJ+CDXs9QDApbB4ygxe1ygURYYmcmgi/4mopz76TI9TBcgBZj/WL5zF/H+jS06KJueA0
6CsS1LzFaPURLxkcjW8JR4fyGIpSXJ5GDaG0aSnnlZ2FaAZQbYwZIMWPLtum6/S/GSwxhMNOPMKb
/K7yWTpqqxn0WF4zJuhVS50MfQbVIJWoO1ficLQ/xu1WRkze+rJyAIYGOccsPKLOno/ai4+ldl6n
Fy7Y1f6ixrXcPK4UAYCmDW5yLhMDZIwaRNh0z47yca8K/vN5iDz4AhlYb8FbFuzARxujdRKyfFlt
2vWPHV5Ymo17I8XYwNOXl25vMj0lzjUo3rhxWPwFmy9iWFdFWdQeqoF388SjIEkZfbgDWW1aaZOJ
tTw51+y952e8C54sN8QqXWiMI8wbkOih7VmKGUXVVdOi3B0tEJYgmwZ4hM36rqz/aq2YvnY3X0lO
Dhumi4cYvQMYGuKYh1HHbl2grsgYAuc4JIO06hIlrcKM1yhTLaA/3+6K1zaeK4ZreV9RJdarIhK9
fKqOHWnA86OoSfJPyIsqhW+HT1M0AE/Vf2kR1hwk3gMNhHEqAQJLIt31PqgGPEQPm+4wcQL39MNz
rKPmGiHoISb6jDdxQ7oIkz75slRxhMczMBWykR4sVipcsqsG/YvmcMbcSouxA0/62t46hwsMb4ue
YmWZibjyWfrYATcZNNBOKl7iwNTgJASk+z8WHaKapx46ICIFm98idvgpKRYAdx0HmbHW8Nvf6NYA
KonJZbUjW89neZR2qU2W4OUxCAvFbzxrZSV/zP9ziNEf3uwuJXXLWBHo3QThs4FAuL7SJ8C+LtX8
/pBV/663aM6L56FwnaSvpxpkxnZVex3ENoa9dlwVSmxlT5U/crLGY0lp/PzZ9sul33GcH4Ghk3YX
Id0TkDU3fWggX7/d3sQ61meX40EKB1bFOhft239Ggg+fBi0Plz2AuM0kowHoUL1YqDYuV090z/k9
d5yQfGOockR3MOnILGvwZtbaeuZEaqDarAKZfGAsWxRTxQpmpzvaC/Zv6wMiOGwnphrSFo95DIWr
eDj4x6t295qQ2L6/4boDuMsu4VqSeFouEeTPtNa8bdSqBWNRZGtVVf/yP7Z8M9UuHAlbXHNUTBGa
uQuVbIOlxLndQctaAwn2s7wNe+NsYouFKuhvqOF2DdiCOePyJwj9v5Yqcrs35oStk35bIhO62ybf
gYxewNoFPD4zEnq6RFs2hvAAsBHt7vLsaD2uGNyd7c2Ob/RIX3lUwpNKTKVf3+2OY7Nji9P4yCkA
hqmh+t6aVhmJz1nMnjVpss1GEA3zZADen9BxLHH1BqB+8ugHllO3OhaPzG4DSBdZx6aql6Z6R3Cz
MBIwRMgoVJWKZUzJIyYEyqwMty+QR/bAx/7/bwKuCQC5J9h6mH1KV7hU890pSpUhGoVS+/9JzY1d
KzHNC966REQ/RG0r+04tmiXc9KB1DZUU7xU5N98VtcHPPN83BxS7zCDSzmTyTN5IlP0Biyqigs58
nT4Pg5+7wsReG2F1rFpU4WAqqoraqWhknQwubxVLmHEh/dU4smbXwA0cs+eJL0ri14fTYWEpOn0o
M0sDZZ+dzSYKPvpcNKFaYXcytg34V3uF+sm9dcFJtCrY9Tdy5/2OxxEsRSzf+sHABAFwoQwASwD0
yYwNmAkwu6GvI5F9vAB4f0TMjRlKeAdzrdo+dKY0iQyBKxEDa+yk7nBHluDkV/CK4RCDimbkYPSp
VgAT4VSWFfHy21ld9dHNqqPrGhfqE3TV4agOvR1ikT+RxJdZ4mJGmF5HavoXgJxD7BqFxoGxFJGn
bA4xih9/GRORf44AB+9RfBsdBspNL9vXeOUp948fALwFn5sSZYaMtmrpraKPhYqCuT3njHBILodu
JCm5UrnuRvXQbCw5VulhysaAxdC6GeC1Z2ycyGg+ioZnpsWTSRtk7VYqdg/BEfiJ3n+SGFGEjfTq
HcSrCOecH6waLLnzUjOXGgKBSYOS5Y+CklQctSAQEOh8xFTv7yLkxywpPJhS/maqRzVxoOhne7gV
AXHFXwt2bxuP0D4VALtKRjpHLBtkhbACsSDXtS/Kp8eqE7Z0VLWZcaiKCdVGAuz8MKHrmi8JxxuJ
djkaOSKyzvZzraoXnsUWdGxOTdY6LlcbpgCitbQuC6j3+XvBgjd33/ruO0gdy06eHQl7u8esXzvj
2ZHBX97nA+6/gVrGeA5DrZRrZJTbd9X990q0sF0oe+Cp2RLmTomV14shekd5Pg1P4GahwXPj6Npo
8W9SuTgQT3wKYIvObCaMcbPJGz7QOrhlgJX9A2ploSWg9UaNKuwwRCHj9ZyvEq3hKu6G+NB5K0oU
bnmps6C3z9MtYTivNPUhiKtTplduN3Z4MqfR22f2v32r9Ph627XSKbm50IhB7XHx3jtSjJIFzdzf
PuAu0drkmxUNQX9SGPGhODJ8Q3fVsad4zNc6dPOsrYQglBFmCFfQbEQ5pSOif5ev2TpU9lSE0l7z
SbQwr657zw02Sp1znk0VbOE34ZlJ4maJoePzKJimKCSsyfImr/+ZA0vsOq7NsLjSPZiDlqE/Ia/i
N//fYOtum0J6gEgXujMqIxjTigy+kEi82H9nblKyDW0Ueqff6zsAbeNF+D364eiBnLgaDT8VI84f
tKlyUeddHA72vu5SBKQKdssN6n9k2V3CD7dpo2Qyf7XIBo/yfvAt3DFBSWDpU5uL7Wpc4Zv+BNjA
0LePzOjJb8QlUpRuj4NNULujVKsXwznW43JzX74m8HCvtyJFYOqXmlMe+gpOUcw9ORzw9F8suy/Y
JbRZk8Dm451gQoGU6iK5Pj4RN6YtUzIbiSPHytmjBC4KHHmG/QuqlDhc+gQxMOoDg2CRbz5zBtNN
rgDCs8Ubzy0oPXP9+jsAB2R9Pn3ehDK+HK9kREhYKeINonAGupnYSO+ENltd1pK56llTgpWknBpP
inQWZRpu5jGNHAmrMiwrhOrukJsjSmzHBP0h27hQB79Uoyg7AtxDWy2fnQI7s/isGrdzxeeWaONm
LIVon9FJgBL2qU/OpTdPjPr9DvfQWkcsN69aBmhhlUgo1pmkePBF9g9WrDBSoCZuDygZwK4coCbY
FrMveLjKkETH+3E4Pc6TRI7ty7r00+83Bt+/2CmAMb93D/cysJ5Y1aZvN+cG2dYCY0gfPWPRyROw
ueE1skUroWRigWRZdOC044jIwstT1sjxLGQ5LBWvpdJw1YISVPsh/7WHQ7AnZKBhBVgOkqlIBUpC
PiCNWGPGEKHa1ievThDnP/YHMqdoHLX3Jnnn5BLI+j+QMfEwNTxG5pM75WLz4Yv55CCKOU6tBzx7
vRY8kzSckCFpN4wxKXRVOEoGN49pi3NJYJm1+6upMtaFxWBRjGh49kFLlidV2CTodfoa7w24HQeA
OMQ7VYK1+I+qJFJjWODCDqfL4pzR3iilfAsre4dwzSayjHvH/r68aB29pMpgqF3Tjxxcxp8oUEpU
TMKwvyI2dofPq0B0MOrLRD6W+F76NxUol134Hl8DJyZGATrmbwZL/VK7bxDLfu/I3ZdORspttxDZ
I9MWFJQMWFT5wPHM0vEehkUN3qB3A3Mv/Iiw5Z0UzvgDSHrkqBnR9IgYtF9STZ8A7LeT+afuPCG9
0JxGTIo36Nfx8h2ZS3xKg2f5NBE8gy5TsktlUHbwNXONh5n2aWulfvT0p917zmiEcVgc6n13d9XS
dwOM11AmR0m/Rf2RuWXTdizgAKT7Lc9f+WnuRjnkePQinTGT7ZXYNgC1+Wy+SCxhEZh4VFHG8/or
egcbf0IWSx/qXs9ulHemMfbHdVdZPm6tWuvfCWKMxRDQyDi/3/YnYfsqIgvntE3e2q21PYF/Nt+t
2FLDXii3SVdaPeaXpY/KnTTTv2s5hCQRMdjrmth6Awxs5LQahYCRPfJqaxXgfsjZ9WNvXKouuIP1
jmpKjf4eMrBMh//gvQqk9FEgEU/cX0lQfSDdF/c3/Z7icu2Kg6QPOboBdtTSC4jxH6UAT56kheGX
gm3yqYIrnZGbDcBNzXAe0O4NRmIf+U5vzgrdy2qNjhGEs6Cz86Ki5r/Uw+aJ+r77R5ocQebIrmYp
/7SFLk55dBd4rEGF/oSM7nakiSzv1V2B1azYpthHgnhg/Y5STWisa606Y8IK8LElLIKj/xJtp069
NVYj8OgAn0Y+bxwbvlp/9usP4YNhLYWcQ7oQUBcZ1amtR0k1TpRun6ycJPrUEsJEF0egBveVj82+
03pJ/2k3PQWpL8JAquu2n0+JdkJ2IfsTBayx1BUscGi+UyDB32wz7DW0D+Yv4AsbqKxMQX4siUYi
Ti6ln1OiSGOJS8LZH0HHvT13bkSWqAFUEu/sUzDNaEEl6rxprean9wB3vFz8z0VSLjTyLJhrlOoP
cExPhtbP/xL37Cc8tgLfKtsWDeJLaOivz1i8jArew2EnFFuxjBYecNjhkihF+AZCNvPHTF2H78ql
r7Wl7oeuW0ihOML7/nt+W7avDHyVB08hJdGCVTTYgTCcE7HjligjwZINIzfnph7B+f2g4bfefddV
e0Zc7icayypH2gRi8i00q0lq8Bigazr2A3LGQOnT3QI3hDFNBM4aZy5mdi2UESDrUJJ4vSd2uc9/
RN0/wrJeNlANQbJkGpdool5k1mAlByK548+FkxoMWKr7rOgeAcXO7/n2I0TKEJ+icXtU5ahndVZd
hwVNZM14etapA2MN0zEq2h//SN5Vho0jGua9RZ/nomUePnMoXX04TucYnmMLliQHfQX12aIbZWsq
65W6a0DLdfyPy0Y4DMAGo7hPlvbCrH3mH/VI3YEiti9QF07TBUTWINe2RB8dJ+7Mhqmc+3GerzdZ
uP/27belYw5rSZAAamg74xXS8JZpHJ8N1SlTCp/lZSf8xXi87GbAFunsLfWQtDDipA2L1seD/zsu
6CwhTPx21V05u8YbW3f2F7M1oD0eLygyc4wZgM+sQ1yEAWWKG+18KrGES+AQ0ktms87tgwh0kZKj
Z5rHUs2iYY7RXV2jB19bn3n0jYUDt6iUh1F16GxYRssErdUkIhyyslb/mp3iSs43IGx8romtGscE
rAJMHMUMJ5poyHqLWYaB4GSklygRtdzF3rqaBWLdzY8vzUbMBGbHPDK44xCFuzan9S3KE0XJWRoW
+buch0QdT8XZ6yjoQfL4SdYLi94aROe3PJjBe/rAqfhr9p9A8aAF4idZbSpI7vbDyDmiLrRnenGP
x2r+XgnfBaqHM+NYvGg+jyVwuVam/GwXIFm+xgUD09KMTkNbAC4Y0T9QOUIeZH6BV61V4zHe990f
VQy3soQRCPnM4A3RBux3WKolObcJojWyAng02OZELyummHKcR9pnkuP51SCwN4cNa7iyZGN67iPJ
PKjNEFcEASdyH4q1uzyKoNK6plPicvwNA2HFakVrdS5CXZkOg9AuUrrL6A+jsnJHoq5UYIIVnhbv
56zoCnSdlTXZl59dTx8B1Js32O0oklvowVWfnuKBCTtZak5diEM7gvG7yF+wqmfli27cUxbJ02f7
KfX394svT2AktHYrX5eaR0v7uLUKF2iJUzEFDd7a0zzLkYexSeILlTEXyDpZZy29dZl6QkF0zWWg
BJMic/XH6uMaYMNL4ItPK/0MlprfZGGXvaiVYtnoLJYGLm11hHw8EeHbWmnJNt/KHEaw1VZ2Nghu
PBjYTEM7EFoNi5eK3ctGYcAzIKhqzg8R1lu4LIUHpMg5xU2uq1cTj583DJv6ALwbIwMRZ8gyR6Mc
JSjyZWonuVpgANh2XXafOWKdBitRDuv3RPe5iz8TihjD4ZvBQD3Q8UaVmzywn4+NKFB/KWUEmqFn
1DWtSEMZi2uT91D3ZB8Yw4/jAbDDIuNXKfZf9J8AdgX9zn4eVpow6YjhfBtruOJNiuYKze4gmQeD
CnBhDWv3HbW3i0/NSXCtqLt9PWuM2OADo+nuA3hzw3LNFEZU+9g/vXLy1/ztDO+meIC/tujy7bBK
eNCUrxRvVbQlGMXUqcMlLPDo01+tR9u0PhBOgpYfMECtPo3RaRiphSKyPd0DTb0CynMeMk4yU45M
7jKDf0CDx3SQkc1vAgxHESk3bt4sN9R11ASsiSkyYx91VUKhoporVOX1Gcl31QwmoVh+lorb2VBr
bo8hzMjewBkuXx1zSH/KgAV0POs4NkscodoGIJWsTgI3KZLP0BtLCGn676UyTznCu75C1CJhX5Cs
MWr1zRZZ71Q/tT4nTBKTHqnxauqoDamvKKwPQNEjFZ9F+JmL9iJDfwDYGUmnHJPsXdw/PXfN9NWW
m5h6h8WYDrxQ6dv+p77ie5cVuGCiwQeKONfyM/oBdw9IeBNrKyZWUEmJtMjx9jiuvF5tyPYBNylY
wp5L+ytjzHpYVe344p4GBb1KXMpqXcUAuv2xQbup28h/iMhrlwIEXsGWWCsqbQ/f0XC2uDg/luhU
CukffiwUeBjrBUjes36ZZGFBR/88qGfawbUb/PgViv6EWdhD4dbKMCytwfygtMNCU/Fo9BT56HW9
fU2t3JDucuZrFSJyCTFBLeP3IP0KbMfnAzkKiadEiYLDtBfgVRBPYqr0Su/RlS+v+CpJchmbKEQX
fVWpTaEfLYKhMemlZ4bafLN3msYKaArOV+M3894PM7prM8pdwghKqHQlJo9kM+Le68vkd+S36PkY
nv42e/qRR3iAseapF6HgboVtuuVbH4nwKXNMCP31NTUiTpTiXGCG8+lMLRjmlOo3X0F7QStNkPtf
P6KhwSVcwqA7PdEXScxijq4fZ7sSMpioCGeMJq2BadpJP/HfjNXpziLyueBlXX1zIU4dILmvgiUP
7rZF0ejuYtgD4jAsTdV64CwEh/p2bq8+ipfEG9WQ0qTLcDaW01oQC3DTtxWlOsp4TZHzg70mPPJk
mS55gsd8CC5KwogttOKAaUpFFXv0rDq5KJ0bV2vmWQPJObbQay0chrkD56PIplupOib8USGQ98dj
CnHPZfY7TXWJEblGyVDoXj+lNSoPICmevdwcxiQUiL4/eMy6fcKXwtoCKPAPAfHKDO1aVElpgYH9
B93qNcj8kEEvY9pJU8MDsWFJ3uTjYkBApg99OKImwSswTVzEkRHBaTMJXMk5cU1HAX0RqtX2CDWP
NTmRR/OeX0qcqWTBx8vofvBP6wg2iVFjUSiTCEXrdrNcvCY5iIm/kQJZR1Reuryp6UA4LlzQnpwB
TqhCmc6qphrL9pF0H5549g6a8KdxenvHNDWVdr42onbSMpXVxpNMSPm6gLwMD/TYok+QX4JOP4hv
x74gd8aId3FBIf2elBsp8rFtT9bw9Ts2rXv3YdMKtjn15/zQLiYSk4f1l/P9tVgrj6peglxQEMc4
psEs685FOWSbwnYu+UWGy59ChPD98ssGuJe5OCstRw1yUzIH5bD/JLW0x04w/utiCLdTuc35Ld11
baDFcyJn1gAOljm3swI5lG+VvYpKIfVODc/6Hy22eWAqkMB2vFhA88HOFg5ExVeXE+C90gxIscU9
In3ykV1JZra9jRkHrS0xRJc+pxLwLbJYL91obRCmgShIspUfN2aTNNfxujb5AblviSTYGclePLm2
QwCZvaSFnxzg6UTnz0rpL2CYYyB1eBkuNjUDWAtU9fUaW8HA9BwfoNSbfz8Ok3oOO8ET0xSP0j7L
KqWM7qJOWZSmWYGSCzuPxJ6h4KvnA0as6ehhJMeyxzvdFKMU/kiBVaC243IjDhK0177+pbZxs5VN
zZHvgykZsoEwBZYZLslAVAOr/d3RTaisCSilVuneIRAJcb88qcGlBpTwZNKKnsZc1BkPiiQZxL9T
YyvHNJpK4wNz+iKo1QUcJtSK/MWYE3a+veJB7bsyrm+HVPgO72tVoWWnQKcG2sXbGF7zn1ofqhfT
IulFF/VzpRLLoMX4eqshYoC8JfauWaiGw7dHB5U9qTBI7avyxods5vqbRjkAvHiND8K5XlM8uzRf
0QS2lrSARlTAGVt5CLYASWDFn+gSDe5QP6QsT6rDNIs90wKCHU4aXaOhwHYqyj23AEtSLpb/avl6
/pBXwyZ0Wn6e3NAlFbNrHdwplDRGECCRj4NkEaymDJpjOA6Z4x0YKuh8VFGfqlFN7k4CtdrXKgCE
NTte8ehZ3fSOc8phr4XpBMEmg/wNFN5uy6cjWgs6BKKGEc56tpguo7Zbcz9RkGVRKnVpWKLyhJh0
IPcAXzeGtvwdRQabuANk2vp3DQNSDctfog9wzt8cankdFfjT6HbMg9Ir6+sB1yOeiMzrQOPsj9bV
dr7ORQSnkCRDINuXjBnOSNiOJcuEVr1vMAEuTkN08BgCDwCHcuMRtFFnbxSdlwPhXDdIXiA6TbrP
YgChl23dIcfeQPjZddrorA3D1kZAvg7GIVuTDS5Rp0lOjWFmmFQSfOtp10rjScKGQQbXn+ekU51g
rWUrIEg0g/ezUxKcD5PgHiMtmSQpYfribMFkCrrZYFctzJT/GVJ1ZpZTWMkrtF/tBNj6Rssz2Qpg
shYbJU+Z+fOr2G4gNuAg+z/nzbvhAWel7FVVSiIYfpw9yB6yDSdw47rc5lIaGMfX/OCeP/9r8WF7
PVbZiNtGR8xIGbBm3d5xQ6mI3qGbspkyAvC2p9YdEL/YnOHYx6jibf2vZO5RIB9hlrCzeIUNMoO0
/1M6mhIu9XR36htyovcHkGTtghkpNeS0Jx0rRrfgiZqMZxPStnSMmb5CSF0tCYtr79YJ5nzdZh2P
+jRbEm7dtwKQaeIKNELhLKNDXLQclDfPiHOcM9vPHsDKSBinkyNDVJgeCF2wTlVmC9f2yvp+InJJ
1kyKsXkrlP1PSLToy5SxKzeiS7vEjvnT3hIBOA2dUCd0QFql5uXoYCtzMLGUZRWlq0PjsEQaicSi
9Gi2vNCNP3qCWSRQi1TQahs0RjxVUVUsKHp67/h/l7r5Cs7RZ/BWgm0l0rzmswdreCbNSlmPkrXB
swt5hds46g4eqz4LuaO6c3AvfUPuI8osYS2oLBPfEDCeFB5LH7k/rowXq4O9oEqJJbTb0aya67HM
tU3iBM+ybXXYguJtH6wu+dinD9KKBUJynitX9rNBLXcChheUZkutfgkLwDZ67Mv7TEleB0xvxIKD
UQzwXuJdv99X+XzSa0mV7Q5SlZJ6k+C/jv4E1Fk+CX24nvT2qigYCPTr9IHcAsD42Klwu/lDvCaP
vTCDXwwRSfxGP0mEkfuhbd7j8luzLGaxjnKyzeBI4H5wGHv+iZVmpQaXEaO9D/7QgbUkYqtNMaXM
sVHTo8pm7Xn9OOECRktLKTXwcKm7XxD0JIB+Vt1rIANv/alDkcmZxyE36tECVuk77N0X3iCV61Gn
itdLtgrdH3oH8AlY9B02au4qhZ/dlcQnET03eGZ7eoN0fRSPWmbywEWqWI/YHaLGEDG+DFd9gdmz
yJ/xZaEQLZ4wA6NM/F1K7+Z4d4epIxkoI7nq408NXI1n2fDgID+CoUIfvFl1ahQ8ebHGUr/n7xKZ
LtCdD1ozPezQUynjwYCyzyPKtx+0nfY6IVY9b2enCxk6cyjuEjwRvK4/qsMljYH4A0mFoUlTs7v+
MTLrNovoXGI2Jr9Aeeo6N6JtQvVwfwC7PDr7w/sC1XR5cus7mNA+BSl9z3iiaqOq0K8JI89Ypm9z
zJj4TTrSG135E5NizECKKBgEIGp0b2IPImTtyX+smczd59i5lQFx7w2yyhKEI9wic8GEYJN81PC2
Mv7eQov7rTFjnhK9RkTCc8/epVhJplGUSjO3FJ7tn+5C+Fs1E50tBUVANnPfPgqR7CbS7fW2oiXi
OFFQly1PHiO+OOLDbcSj6awNuPz+jchssYK8Zg28Xcft140xo14Wo8kSsNw16wwRXfQ4YXooe3KX
i1JqbgVkz/tXT/sA3CRSCFC6AmUNL2NTsr1Xx1agRhn7lPN8KUny3tim+TiisPSjKQNLbAo0Udpu
plB+nZJj7p5vOBxTnWGmZ2+SmTvf0BP5EaI6NueLFG/35iXPLUrRdFLQps7WDy+eOfL4xKkFuZ1Q
z4i3unGL3o2AwF7XdAN6MK6h2v05lA/ylLFG0nmicAfOKpZDt8CM9TCPHzAzshrk/BFwX13jNzg6
i4x1y/P0vDUe59NTmFeduY1c+fsYgTig3Zh7tpmnJGiUeEZXiWAgJC88tFQW1WOt0PfnyrJ5/D9j
2jxIqBFzowAa5ak/bGmEL8GtVvz5ukGBFF2poxVsdlh9h6R6f0ah5H/oFZyH0wCkx4SllAsvX3WK
YH2YB+7dMIByh00a6PrnkBVSDAicAzy8liaIINMkgxFQ+bH9wWOteb9LCgkDd7mAFXgpr6+M/E38
IKB7or7lDJo7ocmsK1bpcTNWDUZduwiS9qBOVXBkR0ahOHyGNkXtIb6d2sLfVZ4lwTNQJOkBUghP
PYC14KOfMqQ6X82471fBov/1PE+eXwVwSJVi8nAI29ofjMkul+r7QS1y+CKi4DeoX10raFYc3IMm
0O/pY7rqwS/lTOP0RqiQ2sEEei6pNQ7jJ2giloJZuEaWT57HdR+2sDf/s4C1Jpm/J+uvBbi2rZg8
AZK3m0atCqlVoszTqXZDEZ12Tg/aublD1xVh0ByV7OQpzGI1zxRuarOdejfCoNSVhj6Wgxz3ArKn
6wIE8cBbkm1d2KiDJQXD+LGw6UUnaaXhLSTbEz3UzAraPOfBR9BaThUAWKRIIkdp6NSEJ+QHUzpa
aZR9F7FvNbaW+Fuj5zoS2pn8cxwVbus0G3yhMNgU0xowvxXMM2oktQILMm8RkwGI5DcKRubh/NYk
aQVHq9x3SmzP7ZvZ/qT5ffHuBKRAn2BvyyWUOX9HaxcBN/9ktS3J5yp2bbi4th4J5zYQR97pEdey
Kksz+qchQa/hyYAfKMZpGw9debTh9gZyHv6WvVqKM7hclaA5C4vbyQTMYlwGS57femCxijIoHmHM
2eHDsiGGORNAWI25rGxFR2aCUk7HcVvw9tpiT/DKtK6GmqFv1GQdlKYMxb0QXCYTTc3xWIjnJ2q/
VfWthJZCeYCrxdQKKpvafxqgjss+gv9sCFt9QfeAZWMzgboRI7+LLFBFHUumhcchSxStAv6++e2p
k8c/OG08kkAVOTlFWtkprjg9wOAQ6mCcTXTj3AaJfvNSdOJhRYUIcgLTEZCaJBOVyUFUBD9zTbyf
blvtcEq70sOznshgBV0hlyJE6W3utfTqS+WNL9X8RfpCbk/GDF0Y4PZ6gjijBtoiJlm6tyiqyLRc
5WSsy/eb0yoRITeqMUPEoxStN3HjfKa8g81dwFTFsgmUvjN7ASw4582xQsdejUh6OZgkifhfkkaA
8/0yXOuuWB8euH+1SewI4js3VCF+Hl2aAE12Wruc8CHZqJqadC6PXuMQ+GKdf3FJjpJxTZb8mndS
EQ3MEVYiH7p12LMwrdPCjyqXxx9c3BIFvJ1rUeVuCm94XtlWiX5gJMxNd4rEwpPjYJpatXxCozyL
1+79CdRhnEAF4PcL92HE/vMNenjKvZY06ptWgtOvKQMb6zsUQ08W/6F4oRMcTVR6tAAqoXOorbIs
ixD2looMXFdg/RwE8S103iNm5oY9CqFHqVvGuI9S8TO3bEI5tybdZNrocCk3PDNnaWZvfrzkpEdB
7YLGZTdUaZIQo48JrEXH10BawGjdo0WfVYqhtPm5WKB8VM5VQw9Zu/32SymksXiZKdVE/w3xh/2j
1kej9xbAHkwjmSqAGyUjKxreElMNSvB9989UCpYh/b4cC/w6G8TKGL4/TfvKb0Yme0an2Lq5EMbN
7KiSQvPArmKKOmZKRAY/K4eJjQvCLNPHShNThTfml6Awa4c07i1C52hmJ5ilmM0H8bW1U5BL2LKR
KHt2gxnTUHd81iOWduijzvQt2rNmWVrUyvcKHXoov7VM2nU1PH5pvOct+opas+vMASRnm5xSAK5e
8wxChM+k+Rp5EQ4I4aq1NvjUISDwYKb9Z8ZcDzGxePIjpSEM9R76F1FM2K/v4dwPJgmfD3NQcQ1v
0zFj2FQERgxVjoK8eqA3deT0pWgQApNOqhvTb4c734kJVbd/PPGGQr/k86zDB3duufYPRMkb0XJ/
3NleLuE3v0qJyTpqmPONvrZxJ/oNF9T7+hX1gMHpJkEGz/+8mZuUD+vPzUE+A6YYPbODalxAQTjC
GyWRHdPzIrm+xNoKhtH0xF8dEO5gTOmQSXVTbjjPMxlQZO+bXlwg0dwwRXGMtQDcjxkN0SI0QfFX
niQ5e9Y6qgw+WJy7kQmpJaYrU59U2M41YwfmTIXCPZ05AXGggXnoSencSg9PE9rdzJYB5eGwO1Kf
VyoYeglTidFk6cbC0juMMfVxY2LslGpTiuTAPplfIYcaQRLqq3ccdsiEqvDROuf+jYMt1s4Eka2e
Wjq4nSkdyDXj87q7HhcJKKT/6pAQbLdBoHO2c+7/+nHz6MA1f9DlkrOS6NiU3GgKbfJEwFF9bRX+
UBmTicug6qtZ9Cv2OGrRmZmMhPcW51KTW0P8w3JlvQKr0pqVEcC0YexRurWfT81LCIkW6hYA9AyN
g8R+pUA9TwpeCQXxH8I2eGZrUu18CwnrsjONsC2pT5/XqJDuIMy3aYOOZ+YRTT0xbhdp51aRWNZS
QVp1HO/C6TKa8ja3GMOWyF7uRKTUZDDenz/GN4JbMsDDN1seNqrwkVLCme41ZbYur40M08mP/jxX
eGoODozxDwVibXOY/NFY5TVPgol9aUth/xYZmrh68EWiE5rHlGZW+hAwdPQ5X7/IRGqH29dcVVA6
YFosG8j5zrC0tcr9xkSS9vYgYownHk5CQM2sE00wlXEiHRNMoog5/a1sxPGuX89LM1PeLCWJnztj
uEeb28mL/GyNn208vVs/T2mFS/TGdmQ44sZHKIPZmecULeF11R6be4V9qYzDIIi4CN7BGcHNV0eO
xl6vqS+rKDWiLTjkmncRoNYs8yK/OIMdhNHR/yIv3uh85pjAz0HyaFP4ao+gheBbvy7PeLtp0ywh
Fl8fMPmg5SFXFHTNgHApY13t8eyP3RhGssTAj6iQRIz140HNxR+5ozQXK3t6zpORsGLb/P+4KaLg
AYfbJYDNPeYE+NNAmDFvFxYPKRY4fPSiOx7W1tbOklpK9tyEC2Gl12cfMQ8St+cDcG/o2ii5zAIk
9af705e9R4a8b9Ne/fj8wXcimQDG8fqhvOJw/SJbk+bCjc3p55LkDsdsapoWIOLdQt02tevZhRQj
2SBWtDpVOi0KVWS4TEUiXApVdTrnL/ImHMkl/RKFpFITtQNzRghN6fOqNU2Lq0GxrwfjlniMAgBw
1NwiBiL9FbYueKrthcfzIlCgVbD6mMLgRHSYYhcID5aPJyIjHsLeARXzaQvOREvVOJOjeRT0aDHb
J7mXMVBmIzAZ2i8V6sBYf340QhzbInIPd8R5Sklqftp/rdg0ysFWqRWtqV6TLU0xYajL7V6fChx9
v+3pOww4VepYidCJn4IO47B0qHV+YWVyYcFO5lHkvMH+NnHFl9L74KtfYXRD5kfFoh9OrjvQnIdt
Uh59fBr90Ba1Qd/9pRzEyrDAP9NsJkb2mT3GIJtOoQ9ADY9fAB7iR8UpZE7tcEY5+vKNPQWMjRw4
mfchN3gMcL7PTbKshxrqy98tCortvqgbEVvYQ98qXL2LyQvtezxltUiFWtLzU/AFWCIWchM+zJec
sHtGcUlbVR0STcXOP3lQC7QYtI2/ZrogZ1dbf1exDvU6TQtnCjC8CRGL1fGMUdgecVmFuRDd3DJx
Ym9wLiJM6c9vXKtEnDo/x8lCp7vbFvRMPLkjFChJQA05L+qq6at+H4Z439nHM8V64WOBCHofOzWe
3HK6Ws4/jv4LTpaZWuzRMiv5Z600q8kka+ctjFm2FT9qH47A2a/OJBVkbLie6MgCV1YHN7Y+hzI+
FThRzsdx1zVLeZt1fm7RBIw/DYFBUmS0s4lCenm5WKgn8j37Dn85HMW7tfpR6gHMSDPprojJAMSE
bRPB2vom521kvymZhWlZDZFrCdoFUaMNvtN/vzMpe5Q1mLedWOCKpDcAqy6f+Q7zkpBWA2XdTVWW
1JLlvApGcpPmUm8uDCbaR0bAJkMQxox36KsQRFbT7nC4s+Z0TEq3EQ4fAbe7/gfBFncDu/wUzXSy
5G7xrWEqFu5846CoBXEKqeovTajZZ4fd2PctolG5jklzYhWJFBhCtTzF9TxBmup056iOlqcM5YSH
wLObX7SZht0RxjEzgM2kVELSbDkt+DSWP5UAB3LxhbJrJ+d3cJtPt1k7C/WeE4L8TKPoJxJFZ1dm
fcxrujF7DZTqlTdB5iT/YvydtF97jH/pu1911C2PuoCjHPoHvrrS/CUyOt6G0kVNrhcy7ZcMbIFQ
aI1UVa8J2AQYIurfccrnrW1E1zm3xNJ0AhtQH83hKrWBnVa8z792hm1DgBmq4RuV/3fhqYpke7gW
4K1zdNLurF2JIgFn1N1TlMsqbZcKEynGsbQW00pIdPz7Jbdzh2a/DVmFpjCbO6L4FbgPHFRGUKSZ
R28LZcJH3k2lwQynTtbEU6/HNNyERbAAjMPWZOxAog8eLJqw5PQxQWvtDJFXD2yxE2rOXni1QB7D
anoWfy//UUwgNhKDDY01+soLt+LIolmBgYxA6D9KWOnZZX9VouksTy5qpYEM5D7mVRx7v0PAYrHV
Dr840WIco/etx4QwE5wVvIL2GbzOD9cqSUD1vArMHVoOyi/xh3TCjTMFXrtZ1IXrRtsP0J9YeHU1
p9cD+nClPQQahDq2GH6TV43d+jfW5VQ6fh1dpUNYTjmkM2wS9syaQTcFEJCkhLefOk6StkvqJW2H
pFToQS7nIoeA2KTnydYz9+sSH71nH4Do2VUwDUdhxG7hU476CyEhugza0nkR30/5LAF08mLV5vqn
ROelqvyZMi7EqqivsANxXPaQDgnrS3yXqRdqowV1rzAjZiQO3/S6pH39yBgP/3QHBHVRGGQGHCW7
sBfm6SRUTbUwyG1vYNzeIZ+VDyp/5xjietoJprpvhB0XLTSHn9CF9qUqYEyEe+LQ/xbDe7fiGpxH
PYTWDjXy2110wP1FYFRyGCYb01YGyZ+IXVG9UatPPd+auaJcw7VoRaOltUbbU0aT4iwzbH4zs9uc
qf+clbNIARtDqu4Wj1DFFiiXWMIejsWKFgGl+qdI/ps7d1jjv3PjQ49hfSIBg4KCS8RcUavzk9Pm
Cg9RBPHXn+pk9B/sXnhfSMu8LdRlb47VruMWRuebtfkvi0YTdMCOKHbndfHqdYYTerw+Ys5CEZX3
6KNvu9g9ga7+4nHzg8Vm1P7jDdUxhKm0p/eIZhLpXJGOd8EM7bW6z55DlPJscrhIsnzCDkfeSuYI
R2vTySw3Cj0/5OSO2Oxl7X/UKhw+s16wIpDCDt/xlqAsz+x+JMLrz2u3Ajqfoz25fnlm8D5L0JV2
Sxmd93byDiCUZ+a5bQIUtcwupMRFPGUbZUo8dB0eOeVRlkfqPyHgNHDSTGpN/ssLk1p0JYWCAhHS
cbe/p1tQgeKRz1JnLpJZxbBPt5TEIGyUHzhWzUcbObwvUXHK73XUvV/m5AwD+oL3RwWbLLUtiEwu
/TbaLx11RlNwypacTZhV+g1swj5m2oIyV0lwbb/WeVkTUIoGThAQY0tUT2caieTsAMpIRz4tqZBl
MPe0uGRIWxaI7Egz8Ca9xTnx+vsWCJVt8zNNYR8TBiktpWYnibu9PQwr9kodqdlt1ppudg4mvHUx
dZ6Oj8AHKNiaVDVCMqOiugV7iU5dbE4ifL/IJ+Bt30znLWgnVgtmFbRPrQkNyrUl4mGPGHCD33RX
xyGyDJcwljhK1+oFtqok6LYuoOlyNCtHHZNqD/N/eh32yh6A/J9BWmbpwyeHNmrv70U1vZlgP0+G
+LTIbuAFkB0TFO+2FP1tLwjSjcUdcPmVgJPnr51HCgHs9mUqWu/QiqMHiFhVLaxT0e6SavqxNbtm
YN/0hb4TEbkrQPHd4TPFMuKcH6AkvSXb6nWOwLhBsPDe2ZFcbtfiqkSbwUQwFSyHGj0RVXNfVkpE
WAzAmN9fgKy3M/PYarRHIJ7xYHD6MPKgOAssILwJAVyM+lKOJXh4jpeH/AAUB7o0r/o9/FmJSvmS
fCq4L9AeD24Kh1Y+8AJav/k0x9gb7OpXi4HeAPmGNTwdRLmUURm53K+kQ+lUH5ZyzcEp57MlhS0X
VEjFR3mgkJ+8hMxPOV+5smSL1n8bar8E8GiCcpmeErP3xeFreTDDXUiGSacjSt5FGJHT/b2A2qAH
I9wJHwZQw8viiTcN+WzZdRBiTIYW+GvLSxKXV5ka0SHZKFGZBW7gzwCYiNqZSQHRFz95BNHBr+KO
gmLT5tlpLhab30YUJ6ag34CXIhF+gyEVQixk44X9PKHi5PgXL0CpdNjnDbRroSChcV/F5vOEn1Gf
EbCcVeWPTy/fQxdwrTS0xLbNqLcKSsmGHUMtykft3pnJ9quHeFdu21hjI2j/QAuMwskbwzjlxSJg
iDp+WkRjIkqsp/Bjaz7cOY78DS7mCsLxeQ6U3ZUb7EYsDVQ0pt/cgnX4qFSnx3iw+CuOaNjUfYNC
Zep6GygXq29TjyRWpbtn0QLkWP10CbDwFRGCPv033EaeyOWzsHwFoMZZfMRB6mvIeOVa+D8NvBOx
BBxG46JiFLoX38QbrcJjbVcqeK1jdx28Cfd25frYWYyNzSaGqMYR7adQwtUdXGjVe9Sye0vRGUHP
HWKSwFspp+AxcEuwjbOl1XJYQqjyzA5G5tyYox7e1yjjMGgskGQqxF+hKCaahF4ctQAQP6imWZTR
xir8OgtD7nr6h5InieTdcVplm+ZV9QvSrC0ebZuIrHYJjG9k++JHh3NNtesqICMSNnw7qhWQHcm2
CVKAtaf1bxJfqeuz10ZqoT6VfxaNKDtkmX9gwFENyf0sKORaOArTfsq1XaWkOafB6B/HM4+SMs0K
51RVE8HPyb5k+InbXDKOj0QEmNNuzGAwGj9+ziin+g9XGG/cJ6pfj41+K581wn9Cl9lN1yMQ2nta
IhJ+She/6PE6hLcpV0VIjmMvv+jr1sZA54drwzvkPcrlc90uPlxOIQCp79/ny9gvcplESW2rCCmN
ASKYoT080iMaxntVzicGVbIijw/6bn1mKHQioRPMcy9DgQx2zm3eyr2b8XUZQvGMiJH3cMk20XMz
pXwxkfP+Zyr7RHvq9UkzMEJi4T5srUG7so9RtX9srC6+18x94MAF9mTCJHeM+VPGBFXFR7F8/2M+
QNa6WfTRiBPDEDAxW3k/Sl1IlqcFr9o0bo0Z+84V6yEDPWS7hw2Mf1K7h6dDln38bS4cDiUjhvpf
AoAGcgt2Vor0cbNLA11Z5DCMmAlp0BnyU6yaN5G+JpkYc4VqQW1EyFSxkC+fDIvzHpaRtUtT0Zmu
V4xtRUImQ0bhFfwMBj82+dNBn9Fsu8qqRmzY1vm7KJtLc8pHzzPHsUrA3S3KSEes5xU+ZHZdLH7R
hJljHGqVsvEpHk+mAdDsOnN+iE8jhpWDxVPgyMUUb33P1XEV7mlBv0dkp1LSp1hpsrCWV1+eYnbt
AdKYF3YAG9Ef/tifCy4tqaPjj9p3D/WWHB6vozDa43sZ53zXBrHBMSpzE1Na0UiDSm5xu/q3ZZOC
spnl4vYzMryTk6nhknc5DFkCrHac06IBVioEWBtF7+Wwkt0BQ4ubIDHZBwcnjEr51+kDNvdhJYmq
WbDUKwUJpRiZ1kJxghAfcPB5PTbBOzOTHKsuXmf9Wxpzaj/j6gpVerx1OyLF6YaiV2L3na5ZbTqK
bh6/2rpuZtaBw9i/xzAkTvZn72z5Ti8sTeGfvUTbayuIAObCRzv76k0XZbY3cyFBgVYwfFuNBSeW
xe22IUhmpe9kXWKkv0dCr62IIvLOSlqSPfe1rTBAfYAYs5cFAlw0Ag1ozSQWs3gJHj8oUg9MIljs
8AxS/bdriesLz8IIlWsVQMd9rOWH8GRsj684s2RdtFq3ijBc1VLCbXZbS68bxbp0XdBS/7aLacM6
wBN+ellqI1L7L/9TT8fmtsy64NLjoo3jEw4hpR1HIT1C6592QqWLm5OMGFUfPlu9IfpMDyPtV4pW
gcBrYYKDHrhELhGjFDotq/Yd22GWIlSxYBkquuaQ6UOXBcF1EKXopOxBGwvUqG5JaqX6u9W06tTU
W4HSlImsWGtVwNvtkzdfsrptd64YwJPWXGKJYazebCuRW0aiXce6ocyjyaKUhngKq7+L4ICLydmh
tnvo+DQBDpbT2rEH3y8OgZ5VpRCg3PsbgmqI0LvqCQDE7jvQeCP7xAC4BqZ1bJbjmbB6ZbU7KYnU
mkAD9fhbrfeYFH7L6v2jVgMBROshjkERS3EWNTx1vViOqQUaanRRzl2IzS1y1h1FViLw7Mf1PmSa
zL5yiZ5tL0h44bx0JTIXF9otJ4MyTU8sjHmR90OGKmXO3teuGZtWG/ni4YSjnbSSJVtzntoyNbca
PPAj/nDC+fVUg02zjsAxJHf9ql1FaE0YybivwgeTllSLODqSoTTax+zYBM4Nwh+KTgvcZv970U97
8A0NcbyTEuxBl87r4aYfLpYlFx/prpf5+v3TGc7r2yRWw5bMpKfUoO38kDBD2kwokI7KYGHPmJID
PAJoyL+GfDhU2Pwi7vpfMy26nSGCEdnry0KLYYQNbCGyyKZo1GwExZUvgeeGOOImo3tS1ZFifoNA
iqO1WLV6YiZYTJnTCxSgm3IVc5GD1DeHKabx2h5+hMsX4VKuylCPuOu/KAm4lF7CFQRG17jPA1kR
2jW/uXziReH6yiAqie0TNuTt/jPuvHWnbFkjGKnFvTj4OveXpC3HAgxvhcQUx/OuQZO1+CBuy908
UtcTCwbh3pNtBI3IB+l8RgWpEJ38pxmjTyHxE20/8TkBXHFmIX4wChnZ92tiBU0IBuQhwQ2an2oA
B4avxf/vJmFVVGTDDP/esNf1EeosAvG30TQ0WcW/ZWUKuY9PCVjnQVfAoxOwJF7ZJWqIdQg2Uk0m
wVsuqd0FMGhWOQS7GTdirF80rcBALfzry6y+hVYPWB4ph4JUhQgK/NZW20fwG/3OKu7err2sY5ne
He9xGyOA7Rnpj5prO9PhZtr11J083bdWEho3oFmE23l7Py5IXk1EVh7YpMmmzn0tlblEb31UEWI7
6QvdS57PnXbs/EXXfcnfMXUPfbJQz4A8azoc3LZuGqLSfvufAors/O2/n1blZQ+MzTqhJLqKMi23
kaa0hbmJXQ6gEyZGDwqGNG175/ZUWms3nMjsbrKwlpAH0FDSGlZjGD/7rgh2fyRoPYEk69nw1mfw
EW4L+E2oL/u5WMcUFpCbRXVW2h6FvHY795hXUR1KpzZt7qqMeO5Si3LcHaDg6RuVQ3h0SERE7HI+
YN6FR1kV9z368mV9V5ZXUBtAjSVGWGOmfmKhvb8cFq0GN1N7UgbqyTrKZ36lCyIqVH3In0umDIrK
OnuCXBDXpE0YMVd31UmnTtqigoKUniHy+IOV6nkdnr8Ybv8uLD6w2hO57bGpmW/2Ee+Xi3XpVj7j
9M1qBmigEWR/1MMYUBefC3vHzT1d2AEwK4qamK+YqBomdk9HhsXtWk12+9ovuCXfNlcks3caT+Cw
xrHQSKMjwHGzgIFZxIeKpnJB9fue8/ei+HyZNAY93KKgs4H8tGjdCBL92ThUygBTOqPPqw8R9RFj
qMGZJSMh07KJeaHZs2ESttmWU/6jdH7D0hqsbz5aNaKiWPyLNSRzq59jOuZAv7Jcb7C53VqUmPZ5
wu5pM0Q1ufX6dfpbSt6ywwoLF+eI2x8ic7mTT4oASiPmpyOEnj/j44njKJHjuAG+WNO6c6aenEt/
sPmCSbzkw/C9ea9lP6dI8aISyIxn+OKXXKa+GfutV0SURIIfJa1KZ+XZaIgr0N7pV/owKbvtH00j
8i/p2hrJwkJw+h7oACDZdKZGRo0L2Mv4U1mvZq00q4goTzmpJ7nUT8uvmpL48rLYCkNOMkYyokaK
eJNKRpeOhyMre9fYpbRtQl0wZF51p20SEQxr5r4q1X5D0foQvLIgBx3EK58dzVTPqawEz2BwCngL
JuVt9FWtvqLcuHZjxdQt5ZOpbkw9VP/qH3zSDg80hTXMUN2F1GI7NV70uuO9nYOsBJCAv73Fhn3I
FDGNcwVGXZnK8HsUoSXSZgU9aD/mhS1BpLdA4Et32lp6ty9G87tzomLiWJladObj2occDcQNqd3X
PZcrwSJk0VHmaICHMLbqld7qJJhMVvxQvK7+RNcWAIU3Hyk1hcVlo8kLCBLw9pvmFDRCQCu/cb2C
g+JRc/s1IWruLKABoLifFVlI1vdkfAdIe68KKKETihA7PpBQoJjs7c8X9sA8vbVwP+CyPSF3Cvm+
O1URx5II3xRgRrKbfPPnBenfGyMRB2wBEt4Ln2NzmnjJ38uK9SmoQmkYULmPna71D9W/vQ7cM0Fm
WVGr0syZqUZCYT/xZnL4SxLDb7l6cI5a6qC2PJvRc4VK4K6jRW1jkg6rFu+mgma9tJXhAvlyWOQc
jTJPmJFsRoQcZCkPDxC1vJwuedBlGMZRhKyNjrkaOelfwY5VhuikqmWDCtJs/d0Lho3qK4uOJJGD
/lHYl3PnTj0ExNrgxZ/3xnQiJYuvn+2iZKEY3WgJ7VlF9Lj3LNGh9hcC4H3T1o+hItQgMgLS/UNO
wAwMU0I+OmNW0vcsooJO/Rdc+V9fRIC6YGWuz9rORLOONKuPOF+79pili0fvMtjETiET+vAmEt7s
e/mtg2Mx/fUMJh4JxHnAY9Q0jX0P0vthHvn6+aTdCtzgCf61huABrW+mdVhghjyO9pPBihb+vpEb
ttDgiriW8ZHXXmSst/GHv2mqeW5/edXSnLQoTjaV1C0eF3C59ompJXWnUBzeTl0Sn7FsgYPwOWKT
yjqCift+5Yfp9LKtlVGx4u7msBi+/dvFoRro2Me33JFHKj3Ov4CUhxTFEyoWxMjGg8ucn8U/757i
lBtxfO7A0L5rzCvZ6wEWS8m8J34DMqwm0C1wHuseFVxSwJwVscBiaHdXRnzRKPz54S77B1LDser1
goqMYyfaRHsOoj/5mYdPtX0rFW0cpW7eFSRSxtZm+JTJ/k6GzXRT0sX6c6o0gGklXz/n2LPZAk8H
otaor2uEV+Cu35Sg4mHoQQrXTAZpZJUPu3dldPIPeDI0pxndbSm/DrlWhgpvkVjWHmsnGMEPa5RT
BlL/KeCGtR2uhQQ5dWSIVaSDtsLcHvQTpI2I3v2mbdghEXFPvVa3v+jvsX/ynsd8fjYlypCcSys3
+Xq8Kre45pp4H90tnn9s2fTWWbRaabqKYx5B0ZNHaPt2it76Pyc5cSsdEr7caM+twA7NjjIh6Qml
tu4zanroKknhYwDKfWuFXlwQh4zqrADWSWqsNVtS3I2/4tdbWwO1cpbYH+Bx5/x4snW1yd3F5K/b
T0QquYndy5dttkGAC+tSbXFNeqc/zq+r8Wlc2AgIngEeaVjDDhNch+tNUtK4K5OBUznK+XZYIfL5
j/xYeP+rzKyoRCD6XvjfPXqVHQnSyLxV5uIjnS29QYeFd/oWsTuXCEjyNHuLHEQ5x4n1DFv99M9d
sU8kh0y8tTRiHowkOnGTUIhj2JgCvzr4I6KTIQe3uHVipjQZOrPQwSzYZ4+MJYid/DNrlg3KXH4O
IwNyi9hIDIdv42Iz7va6Fk3vxEkGCT8NGUn7CKvoEYpwlLUugL6nLVNmRrkw3HwfFEFgETdPv8cM
aPNZhTC/VJ9ZY+uRk3oskC/fKHFVSgP/kCrlLvtNfp9bqdoL+58kVpLgCutRaZHCKAQQ+4f6A/Cj
BxpEmNSJE02imORQ9Mi1MaxqUsC7+0XVtlR200coy7RXtY4/dIZsMQrmy6i3bB3ZlGA27C2VzI4o
jthrb3hOVUUGxK9axfdyUzJTH3KDWQQo7xHEZgLXtBELA+NjLzx0KVm+9VFsZ994quGtpEXlazMt
z9CPjg1mH79uGSw8qc8wjq2cMSHqeLDBU74dsMLKNsQnXLk4nSsm95jbUATanJXvhUZkPE38QOxD
VZ+n1Y7qMpylSNMcznihFgDlH0DRvel39A5O+sXuUBeaGrUm2ryLWnrhuJJkgUKfUZzRj3Ibau+U
ye0J3zzS7YqtpYy5WbzwbhHMGteyiu0HZKf9GEXDF0h6BeMY17Vt0K3GTn7uncImbkCB9uQy9mOy
GLmV4YXUPdbGQAp/FdQIGXHnvQTCrrlzRQLSMcctwRcPasRBQxspKByMqMTUf9bx7rvhJRO6CbNG
6aDfVMIw4ONuQHPN+7PvnwylK2+LVR0q9gQJ0JL8GC0HEgC4x9dQgWyJx5C3M+sbmmY0k6XtRaen
MB+jUADSOhkXc6A1IntlPZr9mpp2Pmez1jN+46b0nMly4SP+rSXYCWVRHQ/ewDLT1Ja0U17OiPSj
iOgNLpuNEZ8kOXjUAhal8MLjVxhIyyRCQkCBQjj3Tpj6v8s2TXvkeoNEnkNVpVR2fHSPzgjCWQvx
ZYJyti6Xwjz6gQXhO33bPJEd4kuWXuFxA5YppIK+qrOKGXxVDsXq2AR1EpC7j4t1XGv4ReqYyEa1
4KoUc1AMipdHxXoA0qn23JmqHu5d3dGGahgVJXBawI1i2uFax4OaGj8oVQ/+I1Gfk+SdRd3R90Gf
BJeZQ4Rf1QxPWbmulxlilLuwr67fNNt1dXQB6TKFNL+cKWL3MLtgx+cHAvhzMx/PnxYH4wZI5bHD
uINKf8oN6ePYyNW48n3qzAW2CebJyZUHqYgG1usE3BZKPZYT6Stu2HoGZKh7tbs2BXjR9c1q9slU
ZnQz83ZAZSDvixzWmlYXO0ECSfEHT+uRg+lxI0zde/10BBZW300R/nboVyPH2wKBJ/MOD8bBz3cO
66HNl/wDQX0qBsvckZ4Ozh+CcUOULaBb+L3L9a5HPxU8LZYgoWxyjgt6HXpCH/W/OTHvFx+tOk6z
GIrsD2gVt9NUDbgwLm7rLGxqoSLYQEoRpAvp2CFOfDvXEsgbPnv6qtkXX1wo1IMjMjXbFjHXp8ZB
KYJFAljrom2HOx7fsNivv2Q/GMenWxfKVfDiID83q4G9DjAdEypGuSYD/66Si8tJydSH2Uu+Hed0
yjnpPt1MzG5T93ZM3iH11/pusXz5SBAzezwodvJiYzzXBPnkXMx7+yqDarqVrFyXtMrvzZy9OWOw
BEFJp3aR2CZcAAHlPs7s/ZDIoi5A59rcu5Aq8YX9p2KKtaUQWkQex9Y4K5/r7Ug62MRjhH9YKF0/
L8LnNcy+6YXllWts4f4EWImQuBJT2hVWFuwUz+L/co+zqRiasDA9BNsmI5yLULWauAVy+T5vpjSh
498KCb58HVt6x89q53tK0kTBwKaIHuFKNXlJC6pHhpwb/pYqWCfWb2HVaqIOSoVzfz3sWtstxFNk
HgPYW263pL4T9pfLGyRCvPCyuZ5xAqQn9SiTBC1qe/y0HIch0lXg9icqS/ekSGe4PH7yz1k3YcNh
XprfeEHxsNVHF07S997HC6PJpm5e/KbE7j0mZSidTfMkHBkXc44ECwjB+gsjI1Z44xURnT7pyBDY
79rzjgnqPihpz4lXOli32gygSQro4ZpTEi5dkjOfft0FQxdUTO6eysN/eli43WyfhBpUYryvbjCi
yfVfR+tqPgHYLnOPO4uScuEiWObbdEEkfKAS0opPofIUvSkYQn9lZ1FwbyqpwQTVcAHhyn87EOLF
iubCK9DKzMpP2OrSMrLhwx5dtmkn2BHxKitoXnZKM+EKAd4NYbdvZVugUzgj55vF/TTfpjMHRf6L
mAHa2lmrkp1vKhA7ytyHcFbk24K46cXLvLTMJwWnqAGGYtkcJHVNzBD4XCqQhbC/hUXP5W5PM10y
1WGlyrkbZ/qWFzZrp2dFn3JOi4eJYFOOw7fXWnkqmvEvUa4P5FXpTjPEsik0op1IzNj1sNGa0Sie
vgyfg+u05uR7QKQ0tGQUtWmt2vRKdOcUdn2qZxiTi8QGg4xI3wWLonESCU3kySlhbz56LGF02n3x
hmqvxjqN1Oo3Ixsp68vzdpc32LI/8BfXOPonshVyKLRmhoo28nPt2RVrbNWUztRHv6JkJktP0FEG
+yQK99IjTSxjp+iyWfTChzoosbDmOun26cQcvXcbB2l98TgxwVDMkFZ0F5y2R/bNIM8mujXY4KFM
dup+Mv13ljAv+XSfgCKJAtnGpO7TXyNcdsPO2PK5fww59OG1xZaW0FiT3QPP5ZGFT2BrpY+2VfaB
BRA9BeeKXVppeBsFnkMByOLTNNvH7BZpHl//d1F+9DEAsbDcBLcdXTrw7tSF6bSkKLkpc5up0EKD
FvZSaasyF9xzDfDrANaoVAV0l/ASNivBO3NkE1/GwF4xIcXyzeL33NHeGNBjMmtfb94TAsSTT2wh
zZTbGxf6oosyVMAocQrRsnfEoqaBEKtO5M14GR2N38ZAD3VD4cwA7MzKpNYt5TGf3jh3m0Yprz37
vcCdlqCB+O4hmzG5eRk96Olc/Jqkun+I0p4X20lDNBLkrC/3uX6fI/AUg6UBDTEiygyvGluFBas4
HZpRWNp8Tf/wenG3xE7DF6D1xlbIKPiM61VzhBMrxqyNpCEErwwK57Sz+ThPnvBIUsjqnFiPnMlG
/cVfdenTfc+4O4WsVyjJP3Y8PXjVbZs9pE7ksf0bzuuFWQYdbKVRogAEzx1bD2/M+7t2cMuwgse3
8IymeUIrGrIaWteJuPVcqsQ6feANGRqSYZyp1hCBKiUZX2kDk48TbdTVYzJBJHPTEpvtw9VrzbmG
pEKE6nO0csH2InAWVQMoWuC58Vny5uIAgGrmpEGCs8TSyb5U6eoyNthhUHuGVn8+LW9KEUaoyFlS
XEKIzZOUf1T06mqyUlN9iT1/7bIroUaZX1bTBn1F+PabX8t4SJXtDuWo6CGGjQzUXCSQ9yBlOM9U
j1qNYNPmhPyrYvYAzA+cryytawO3I9zQVobU5ZNNsgwKtO3g8L/qcmUFkSSNU022WhUXg9QF7fW0
fnIoKVseJRXh7CO9JsyjuBShbZA6Z1UwMJr5c3r7KmnWzL7/MUDMkbhxWd7Kuy7uiapy6o0b+oLQ
DPvjEC7RDhxG7rp9M7yyFniG2MMbC8XVXu0buQ7/CSQSFE7w6Ieuy7G8WqyicCjRAUrJBqy5ZOwg
rJHDZnuf868iZlRK1iTpkPSkXLeAuWCD+qorlYS5mFg486j0U6bJqdoNVCCNxupFDzkQDt9GkdY7
FgXnzyhcl/vfZpcRIB5bIHOMyPSH9svRNl6IFBqB+zHKpdbambqDTiuUHzwTbKE5IOYYAyqVPNXb
1ZWxw0fNyIqPHcAR77ORCsM/CRnpRKyu1W48KAnQ99U9OJaB8+EO0ROdiryr80XEtkaV4n+tn83J
ABBukEhpoc8ciakgSeylHgFB4hEIzgHxoZGwP9iOhUHA+8fm4vRtoGGKKatBBcJdOl2fVyZaSpsp
SBZ9Nb0a2OMiNnMUrkIWY+HoiG8HW43Z0CFUBhrexWCX0fFZmUGYrmXe27ZCWRSD1vM144I+WqFN
+gbNV94MzjF6LTgGXXvfb2aeVPLHP+t+tmCXpeLOZp0QJjdyx17q7RsYNTB4nYdlfUFi1O4Jb9YE
apQXscNzMnZ1B7GA6wII2/3NMl2KhygEhs+zqlelxJXPShXFvjtbEc8xPIQPear/SwSKlcj68ZRp
XuWqB7Dc/KCeF8sMGT7ezXGcaMH3yNJRBpYVHTrqbtOupDRIK1GMe29N5vfsgJF8yUyhNPJN99E0
0DrwzcZ6rcVZjWxKF/Fit8RmXLHAsLYoi2jeZ6qg4i+IzKbUybHRJsW5aM0kdAt/onl59bbO5FCC
hrTztwp4cf3n58upQV7IAnL6u+oRroJObyI7OQ76QuLGCY9eyyVzKsZduzKKSTPqUytcK1SOM2Xd
/gxvXp+FNrO8MFZn1wmLYLe4cVarqt4wB4BZ76F65nIE59qzkOcLlwKRZJBbCevKQ7JyHpr7hb0x
de5vTtW/gKA5iTOS/ZTq6UOgjQ/sXYxg2VrDNlTsFJ9kRuWe21G8x/TM8/KQh03G1tzR6YUZem7A
ve/4rWeePmCwTjtzEQzKjAqLy5fbXSHofWM+4Jl+r5ejImSO3BIJ7JyU93JgjVXpNuOttKh7Ba7a
mMgY3HDEjGPaUa8Pvc4Fpl707W+qLmgS4f6B8so4R8DWyQHgQcCffz5py/e5wX8FfXtSR44vdu7i
am770z2dkgGQQJnBalcbA5aMyt2suhh0uWR10A5EhjaNuoBQ5HUnKlqcEKs07aXVKJZEhK+RmqH3
97R6lQ18sJJoV1VoUBiWGDbs8Meyp+YeYaFWGHuasW9uCg1lrjYSpAk5zNJUV8C6RYKR2tMRzWnR
Voc4o1kE1eiEwSr9zmDY2WplBfl/kMWWuBXmu/X4U/wJwrW+5f3XhKZoe5lJ8Phsefsh0Zj/G6Re
bxuilusfth3orfNQlSkNB6LQsEVFhwGOh5WjkGbaYM10TkQFsmU4LnFSw8xKya9Gsgh7WesVjnSE
eOHNfOBG525F4oz5BCBCZAyXo8gSpJiaqUVDK8V99wYHq9LPPVSkTOyMSrARxSdvdoXh08Mi9pnU
INpdtTfwoXSniTwMP7Csu4Ms1LMq+2/dwJ7iKCipXtvVorrql1FUfWw5B6NwyAmJ0vg5o8d3HsRj
fcUkDk2hBAz1xekZNcPV7NY5XhRBTotKsGnlCf95NfP+WMOpf0lyFDIL0+fquxiOZehXL8XSEnHb
0vxLLNZXq/l5Uu4Xq+TxhRhxHkJ+hbuamzB6t6A82Cp2fLrNMHkmfbdhwxRBudEdor3K0sR2Pi+M
FukPmc1MUcESNrd7oG/OgTL8zly9QTPm2FAumljdAwKPIIX1BA8hHkptz8AWI8qOft40mVJM4YXe
Im77XUx18nFFz25QkXyYO3nBgosM7ydCcbuEVUe0wLOF6YDeApMfeBhPHquHtaMz+7j3J6/0GzR0
Hx7c5cDR7I4gFXnkZWJlmMDIYgJ2cpOhyuUO/siAEjRitjwYk/oA4NP15Eq/BDjcYcRz+ltaDXEF
Nth4OIg/AQVYzZZ+RN0fUR0gVdH9CD97gQgHH/m2hMQbtiG5CW+WgaHWmatbkt3qjKq/Yip9f0Fl
A2qipCKwV9O6SWrpPwFg+q+H/pguDmovsr1kc8BV0IwbPWXK9NVT/J6+RPy9jaMmCNAacTH5fuxd
iaURhjTArphmOqZjVcCAJY1kEEI9P/m8Dc5hgKcz+zzKfh3EHhWyvopJ4dWY9Yy29+OtEOHppGpr
TJE54IAxKusYzIbrJjMMehBFmttYKP8mttNkJEYdOHuZPre1FrBZe/iXBdK7B0IJarqRNGKif75C
1QSr86ONWgwQlhn5u4uW/Kic/aVBRAIfGMPsgBW8iuBNQqwykVut4/yGUuqfjHywqZdqF03K2rYl
Fh78c9cl3qNo0FqqTrpdtv5mNTh69Kdix9dU8IkwTLKtnaBn6X2l88SdhUvyFYkPfd2UDkWQuxCE
j6OyuBNQf6k1A7a7W0DCARylDCqJC7dWflhQfR0KowhI31wiYnTrPmdmDwEgw2H5o9k6ko9rxNl3
/b+7+G97kUlcZM+ZtPYQnVkvgEMT1iabcdff+jdZqtA5CrZLEkFbH4q1y2P99lJAVj+1D0+WefeG
8wItEzqg2uC3UaFqgXpmnzn46Rakr07s8lboi/+by0FXKbzFdDiAD9YV8cf126PK5D5hy2zQWQru
AiVK9mKH2u39fQweU3fWtHA88EqGCJB78NfGuV3VoIfLdoH7CJmZSswQYrgGljuaktg4MJcNB41v
q49yLvfrJZIInRU8PuOqtVV6B3eUQOTpUOZYaJz+Tv8baQbXt4ihMsNriTTTjY2mYsNlCHEwQEgB
kU3Nm6hb6KcTKbTILFCuT3IjZzbnWMohUe/6nkLbJ3c9SE/Z9APh1t82uUTOp7fu+zlbDZgjQa9v
fIzcRmgY4H1S2ivofC/1sy+DuQtDz704zX+v3h9/gENTtQD6zQWkj1IVAGycDyXuFuar88CUvHWC
6BScvVsiyhC9MnKQMAgDLa/tj85mqjHRKKAhDC1cbrlP11OfOFvStNY1QZZcqspJJScBifVUggNl
wX3aFk/tUO4OiXtunN7dsltXXvMsUepk7gzzQIOm4eJdpXN8VazEorY8iV20iMobyVZJ+CKAt7eq
L0mEycLEL0Zi4dwuFyWE30Q6zHZXvERIkJGb/f0Rv9xncxE6t0P7jij3P+7DYmrj1OtPnu+W2c3w
sih8uQpU4/RRv3FsDCOq2LIMHHgmkvroFAtVCluMa2n//ORVYw2tGW/UPD+JRZLQhfOHt2ez16bj
HcZb2YG8fMotlwSJ7dEbh5Oc6vlAmjLaLkJh1u5epqEG0s9NNSvxbA10qQ1nMIM8OIjIcbblF9es
8J9XAMaqABk7iEmguwdHyrR4mvBohSLkHHjQfNzXQ4p4FrOpfFPNB3JS6T4+7Ydrp0oAYdUFLbFD
+2JEOBCBEAEe7yI1rSpSXnkAriSZlzJoLFvVE/uYFs7cFbaCBAFKAS8qnzDzfb+Gpf33ZOxhT9Tj
alL1vPRqwrd1eeUi/c6JyV1PxJ3bVfXAxk1gZakz60jXOOzEdhUzPBTXa+DEMw/fDDROY/6BrP6U
HN0Ef4TIwjb+4HvqGMI5ACdvPZhdZA7GxjCJQi67TE15pb14S9CSf1loynSjztFQrxbbupiPrkK+
FnYdV4tOc+BaNk8kfTs9ccXPOdJ93YyNvTbqCFkK7Cl20xoKyHkA1eRQt1137UxZtig9uH36FSZy
uu5+AL24XPC8BRJRJrdS6MfvGicB+3SHVmBktxj8DAQW3MUnLka++P4iBVJFGlz7OyjSSX7Khyq0
guNws9ODlhNpVxFGRiMu4aduhcrZFR8nd1ICMOKR5OW6yky4z7nyJt+f1IvKofgVLPsyT/CsKwM/
Z+aJMHU1cBDKM0IkGzF+WI4K8Kkr5drAEeK7Xidw/dcvkHAJu4WPnGEGC+PTOr7sLZ415dQkBQ7r
qRY3Q43YulZyXre++iFdQChqh6aV6ki1dBsfG2WP4nkiI8COZ24VhPEu150NvjipUG5Risghxxm6
vwoICCqqu4PIlN+9tXSQWJ+kB7gcIkrIZNckdxswM9IqIS4GC+OKT3AuipV0oxdoyRWx0lOfEISP
JNjHTtENEWCmjd4xHLg1WXXJRBzSxRd8dhTtgwQk7rL4ndVbGL7oXqeieGPzAtTgSw3N7UL69pug
ME/5vsn3jFUZlZlj0OHxwLvskQoJd5mtjFAji0QDSv1Xul94t+tJY9lp8OMc351F9OpzBbYzIX6a
5i9KMVqQYd1RP16khmidz/xcmA+HBKBX29HgW8CYEQDQU530cj/mB0K8RmUBs2Gcijvv/g0lwKqM
JtcrefGZDpPdzOTS0tJ2VQJjuGrOB41qDUSEtCWgl9dgqegfvX8rsScFA/C2iZpSlqpAAV5B1C7+
nLns+FSeKDyylBiF5Sxu4le5ROTrc9m/uDFR8o9Iwetav2ocPH7Lihia4tMwstVG8+wZIz7ZqfjL
OU9jzxjyeUcFjsSoKhjR2p3Y8h+g/xpExGI+y2m3jTApBwj/4VLmtmimGOnj1QYTNJbapbbKfjyW
Ii40+I95oJ+Kzv+4skNPQ3d4WR9+4C6WPu782zjI9T1UlgX2DRZacscWNiq5GsZWDgb3JIFeUX46
Skx2cPEW/H0ztbvyItP7lDwlyhoWs/b8iHaCWUAFPsM53oOlO4j4JsVCN0yRCZhw8KB7Z59Ka/Ve
JmUUjVaNU1uwoUgWel6JbLPcW6Lma9LUGE2BgftOdShVYUaVjKy60Cy5dYalucajhgBWVmPFfMTC
N/6VsAwegu1br+LGP4v9hR7HYdbcFLMMNI1cL06uUnSoGiXRlUNO9SjHw6ySHE4oo3cFyuihJ5Fh
Z0PPHx0hIFzNuKnd/3AZz3a44w1MbEbOq6sGOlLeRV7wHzAzSdpekY32jKkWRH3xCkYrUAY6pXqN
16/gXXMq00fzU1DNvc27vxJGBaciT/X2rDThWsy7bTMMzblg5RxntjuMM4lWKDi9v8s5A42Jc1Ua
Jcz7m+wFVylttPlCaSgoMVSxtV8Cf0PM8TpcjcYxRDuX407jYtwERj5urh1MU2zLc03YazbItujh
ugzjeu/rPKj3Im4r55bzvXz/F2rpGte+s77YrY7QgfM0v+uqPPM+JKdzx/Xdt4PGyR6fuTftEfCY
xrPc0L3EDTJD5tksg3b1t3cgYk3fu4XaAf6A4smfH+YT2cfrxTtohQKkYEAmLP7OWhfFVmi5Ictc
XjVjaOYbi7MgasLde0qBNEzLTfWLUuvdIPfYs2dVx90HI+nznvY2L1NKxTremngu31coJbgU4Udb
tglPai/DJulqiAtXvXT/4zLvcmaBaQxMaURORYVmk5FWz1OiDRzyCbluWFcxE9ejvJooCnTcD7Nf
aipwcfyIPtJvVpNPsucO+I6IC/Adsjzwo4/UO3eKB7l5yoVyEXkMFyilLCA8D9GuyjKVLRqMbJ7D
gapZBsZOLW8hKlpgpKqKvoqcEPc+KOYbPHh8ILdDgkdGLLd6EdwLT4cyPcL1gpNFXMhDqf+ldaAo
plK5+I+eEQZjh38MkW4UiDKON2FdAXQDcFRpdAlWSSH06rvdMFSUItpUN4Z7aIqG9cnzIeWWqejl
Ea+abaYzqJcg2Gg6H9KDxfnKWYP69oaAefIkw50hchEQKZtXKxIi9e8f0G+w+c+4dhLoWZis0qFM
0a+0OIc1HqMUshN++gl2MLmrut9hg1IG0lnQ6IBPB3LX4rywzas2EjDWjbBL+QKtdl8D05hRS+Zy
hQbSgt+d+AB4mArdIB3O+XBvAzszK1X96wthW8QsYFaae8gridkZ6EHRkMJbsI7oxEqzagwyWDlD
4Sb+dT1hmQBNdmH4VxZDOJPLE6HXcw8LKkDES3/T/VmuYKe5jCYVUY/eycvkmDg+5dQBa9Njodq7
Fm4lb7lUrI3DKNQXtJZSw9YREKPnZSX2klbOSTQ56NGkxE7nJzMBSDqw+qFYXs2AjVTz3ExtHU4n
Ei3MIoaeOe9Hm1riZqrsL56B6mjL3z3eXj0DX0qA8Y2jZTxuKrR1oxmKO43f7qQ3gsahyhkpoCXq
ht/o4bceQNkLl9NNnPYHJFOMdAn+Kq1Qk2IHWTw6uY10rbJMiUQjqKyfjt8Ca0rFaYYw44EP44fB
4wrmr5tMFZDd0dqQKNdabmd2yLZj5y+e/zAy6jk0pg7IIxQbqBhfXjT7cp8tahjvyTtMR5C1LS+J
zX9w6h13ZaL5IgF3tFoEulXQMmye/4Ew/HkO4Q2Ul8qdSHr98hMUNIajgXdc0u1DcYPPmwsF5leJ
oaBcTp2TUNZAjzP4REp1WoXKZjC3mlIOeEmCG/MxuR/1zFeW3cKc8tEceAKeFrFNtTaS1xnWVhel
vDLTrhaEolqxhv84dHxHGzMqjQRRZCPNw3iwupgbmHKqVHGWxyVjis8S0+Yn5/4GtV3FZj09E1z/
dXpFyZ3lDkGCcCCOBP7hykw4BSsY+k4DIRKjzHgGuQok/iSuuLleUPcrd/4K/tLI6Dotyvz4nR6O
jYTjRtBFakFPqkOkhLcyca+57M3MNuHDrcUZsdOTR2HWSZ8dlEkeGyDxILJcrmr7yORyPO8m/cC+
wyDujlYihSbCQuEzrmd+rPIiVUOGSnXTG19+YHD2+fpOXTuv8y/+cyKF2oJs4/UUP9BsONm5pmZS
xCk5fJ5+j1E/KGdb/3uoQM8Tq8B+tBpfkPsLnF6Y7XwlN5CkK7S0Nae/FQQPaDu+vZjXRDSrgwIz
w0z+CYAXWyQu3tguU6EniCJ8AieCjKYUelRIc++qyB2ETH9o9y6QBuSnfjv/Svct8iJX+KATzrIn
DTCLhAKMJ5PCxiTMyWiquB0i28f9ZKNdy6LhhGe245LSfUyN6P/cQzRkGAp76bXIdHWvYmFqf2sP
pvGABAcOo5+w9eQqVA1DnaQ3k73KglHxnf+jmzoUwGlfY+H1hMgwzNelJoFo269IOGpcvUAZeFw7
HSharFkm1Iyc7j9RGirp6cVbpiCyCrPKw2GxQ+n/hjbW0Q7lOTANwTk5MUmzBTZKAmo97UwcqnQ5
R/dESca670C3s/tXdrwecxq1ouVuXTG4Noq2vMHCNtClgRf/Srkv2G6Fy7T5fOdryv2cdx3lEx2p
f5mnKyNKdpAGNgZNLBFOye8qhpys6xrB4Pw+qE5ty/GW5psS+DC4BGMU7bJTLWTL6c+oO6eWufzi
KV1KXxTb6ycXxdOfKI07aZ96crvfHmobe3wYdIoirg0dBFtVxBYbLdf9QSktPZ161SteuXaW3rGR
T9N3xkBaQGfkzNlJZUWedaCAP9zrjW6bzFuqcBQa2ei9tcOg5xAatqN/30fWD17tDOTe6vhDOfsr
3+2AqsMOVsy8rDJ/6JDqDnPqFYPvRfjr4Bqq/5fjMR1kQg1LOEpSp+3/1HtMZ9CLBI1KzPHkDPZe
aVViWZA+ZHtyqIvo2atrviFT3w6sjJ+0ToepkHeJUZeJLOt/KS+h3KYcWQaZUyjdocm4SvtSJfkX
WzuMz+jcW/MwUQ/MwdrOfo4bkMcGqSqbIiigqDK3rwQclKAi3dWTa9H1gh0CCNHsRFGAlj0Tzpkg
8z7g7g/s5xhEULDKqhC5aAZmIUdI5NdaxMRTGvpcn5eKCnhs60nVQ0bgL8tDC/oY5+2z2192YjK4
LhF1F4d76gJ8Ljaxd3/il54q2EHMvgFskMxaI1Mm2tmwyqKXVgBQacLOJOHQH0tlXKQ237s5WWSa
5NDp2UVW6NzI0F1352MgRbKs3+kn+f4cCwWfVhs1YhoJstXdn/XPY9saLChYxpkCdh6nv2V8hIQj
igb8dHdYMpDc/p3aADo4Fux3pz0kOkuPzuez5zhfz651fvzR5qiPtGJmDb+DmL5WpDzBjA1qoyMx
jO6PdKCzfyeoa6Q15GtyQVB7Lo6ohMkEqfz/ruT/xap3y1U1RrRmF5xH7zihMapn92qFz8VUQn4V
IKCjVEySx4nIcfRum8GyQyL/64UO9/VOjR7WWHKW+Rygh8mqRcPaV0CXit+oWgGPdMfRqOfjpmbt
ZWrM6nJkbj2RRet/n8t9axckGlNn6D+HvUxwXxTvn2pv958fUKaUFFRr0QQzruo0wrczRGEC37GI
KrbnKAzx4OckHE9GxQXBaq91WGFCLvE3K1SZQZ84IQP4kCjJ3Wu6+9M0Ej95l/aguzCCTDWEK+qU
Xx0LdiXCEL+f7tGTndomdiuvcU3LfT2Yw+laFTF6sooWPDtQlIqH5Lo9P5L0rJhEs0g0HEpDYwjt
h6W1IsbCta7XFV6RCPzcUc6YizkTG6oNw2dvtT0E1dwGcT0C8Qstc+1SQjA+zIG4nyDnDIDhMDBI
BiIrn1W8VV0BWOoJ7Qy3eBg1FlAgQKFDC5CFKnIZdGd6acKWzvD/980mls/9UYmb+6SW3DggzuEm
tuSrKtj15RBvZeFHUgnZwvfUVANUtLivikHwfNOEqGhv05JKtH7HqOjqUUNdmc+YGK+5YG4Q2j5R
qZkshK190kZs2LMGurlE6i5+y24mBosoX1JdfIsDpZDkJY7kEMJ1NTcy40XmXkUkaQxS4De/KK5J
iprbKzsqEpR+loASnfjoiS9QHAUMkbElgWjRKk89JC3v1PL8MuG+fHJH0zFYCn3joKVYNDylyjU4
jhA3qitNU0BOHe4ve/DehPVhgFBkGIEKVyt7wYvFDF1Wb9kFkHoJrhidDdNjE3e2fvHeFZ53NEVt
0hfeZcdlwjU9Z0K0nXXrck3aM2bgupmbFJtuIWpgVDkFaBxuH59n7p6l1KWBlIis5qvTCMrgXZuk
cn3Trp0IYKTZ0ksmRHjoITWbhlcLfmrPaEZ4K9tfJhg9TBJ1w1wFtgZESKh3rosO2JfvSpmapV5D
XoVMJRQGvOr3CzjpVfTbBS7oWwdiGNd9WpoXccnx903kbeFyRnSuK+3KNiZLMkDHkm9njBRuI448
bvfz6XqEMKjMP/3SpBHfQxb3NMSasl+donKlwdVp61kmv1V3OiWuo0fADohyAS3JTJ8OuM6EKQuP
TREH4fBYSBW/VMcKESeXE9PTGZMt0QZDtW4bRXpGsHit9TuSu6SiTQVjGvJYeN1g4jwT5j5FrzNr
SgEjwEt84NBRWtDYam2VujjoUGFilEhm8TKRFiHICxbcpNF9p82ZuPYfJbpJnq0w0zKzYNQVxCqz
/tHX7K05Vo32aFVcjvphwB0PJm6Ixido74p3Opr3h3uCZL3RyJgSHjkhE1Ca8l7VMzrk603jixDp
A8pIx2+gCz9BvjQ994fgQv6Nm7eWFJzGjecMzWJQaClMxSFFIcu3imoDddqP5c2GvCyZxf6yLFMa
yJI3qddVk3Ico/B+q+fiRLbKFmOs4qRoe0Ost5WkMiBIh2aLoojWFjpIa6HYVK3dG5ZfijubF8fX
CceD/madSGMYLhv5Jxn6DVFu2Ryddhis85KJVGRibovapVCTa4TxlYjfc9SNAvCXnkwNpKuVXU92
B3U1ty9DZns3EsQfykO9bq0qC/ORQ35lXLaEb6NoGtZ5fndXy0QR+6MIwWfloeIVfZNvfbDShjQS
u3LhkUUAAfjDe3IZEGKLJ6jLRUEjprsncyRbQzlbo7jjbx859TjOHoo01auorsT80ffdIZ5Xuh9s
C6bv8CLUJyZa/JNR+SwLmph51BYdJSzbvlk74TcHZiiJroapl4GddP1GegIgVGE9JkhNBltK4R9g
Zv5y2UWukxgCSBUjuIJGJc5EZNprAWz11o4gqqA+g8cjmmy2/XmIEu/Yd4gTg+kvdRUngOd6O04b
3oM3FM3cevgmVmV1Rafp5TFSl5l0AHvOyZBFz0bEsj9Go5I3pANWS8RJNFSkR/YUXptro59hGBuY
o+VXaf34OGZNfz8w2rftN9JnstImXgLR9eMLfqWrEkl2mCU5Stn73okRnbTMVC8uMyjOpOb85Qj+
4FueRXoE6roB6RT7eDOKmQsAWF+upKVoJf1FnGmRXwPhyVV1wyy0L/JVyBQRe0v55s2FMPrXeEA0
a0I2vEfy4XXkKbfSL58+SObfgTyhOEx+APLxJ0CgYBiInLPtgn7MliOpUB9DRZzop6nB2wNQfy2E
KeyKyir87JvjBs5w9TNr7FDuxajFrK3o/tI1L+cnkpzi4+CYf041oiQZ/9z7JfjgAa+Io9HFd/lh
LUoharpggn/h+KaV/r1zIrTNSeN1UVBQqcEHd+5HZa06GnEJ05ze1HnjakeWIWClPQzSjWbdR1Mk
7EhU017eXQoHRhhYMGA+VVCsnyWKD5bcZdZb9CehzKD10zXd6Tp3Rvert/JUT8Ki0v99n7zjGQD/
sbJwnmaPfK0LTQwZVfnOXEGWB7LmQ3Dw8kMacxSKgT0n2oe/hgPZ3iFECSCCUPXHHn6tIsSCZUhr
1tSB/dUFUADk6EZ4SIxnr80qHRutMBrTnu4mBQoNUWnaKtNT9RvsfLaYq1ju7sNwKOfwmeyNj3sK
VOTMPC92m8ljm8XyBHQrrfbGU7sflHjDyUs445KAwG38Zbp+3I5s9j7OM+8ZkInxYHfB6F3qOLH7
cso48d+epT9lwUDGSeNCqn1Ot56K2kJQxpHExBUfGwBfSKr5+HxGhQfF3C2jUv2oliq+rELXglEf
uiJ06YtYpNibUQDgKiLi09gjV4bYgTZNtIql307a5+dci12M7dhKXNuKp/QSalykkuCMlOaOu7eh
QIbC2WbZRpPE2/TYhHH/9Th7yIOkhbWx/GMQ9Hp246Nl40pNxtgFA6dNFFbyU5f4Q+gJkvEKANj9
2PZamb8WSnl5MwHEeXf9G1/jhysJttQc+whOM3sOw5/E9eYxvijIROLa3rvA8Eq+lNXBnajtvXRM
uzc4n2YTZT2YqdFuBTnmd56po8b/0BTrq5N+QjZNqHYW0nuCLzQfFjnBXipEb1pPFR+MY/2YgC2j
SqBqEiIegT9Dcl1Q72FySfXXGNuaBRd4wDOkFoOMywV27j8jnMI+NvTy+Gvtvr3fkqPa/FVq3rGx
qRLJ4xWUQYSYHq7lRCiOdUj6sfK+zJSy8Yh4P2C41/+e06Shpu1MXzo7z4eJqHJ0wmndz85QIdsL
gj6HzCVU0k709NS+pxBR3eFLp2hfzSVAYR480H1656ZhDG2VPQep1vqAlgUxAhzLArzugOgstwFE
g7TQe9IFVwGNz+s+/7bWm2F2iptv74fxyDNRA9TuhHj19lrr4RhJJceB9l9BsONMJqcOBd6+JZ51
rww0zl6kAEqEZCfhCDvYK5DHZ74Gi9WIoKaTPxo5D4mgL4pLKKF+kk5X613J04XvA/BJQ3YBnr8X
ctMHZsugzA3yhgxV8ARbaNpRqTV0cZLYLDFbYjaYuvDRDEX+W98WpXONAHEEc9IeMoflOatjNHGi
nMfXZu+fKjfyja4/L2XankJ6O3BC/8zO6g7KTMi5fnlWGB8By2nObJnjZt4a1jPpJZwc3gwp1x/T
aDcRxRxJbajYQnF37gXcQPNm4SmlvomcuT+yBnlqO1AD1EE8Ii22tdhHguCfz4oUC2QAkiXDCxSE
a87vfxeITZMrhZlfdPcNWmCmx3zbOZrxP+X/Sg/6sJ8fjayZhLqYDEy8ddX3t8k2D7NusXM9/eRI
XVtJVkK3T0/5lxDFzXJvj62Qmbxdsctm+6/qNEowkPn2eam/K2o35JW/Mp8yJ53cOGYyE9fTKWR9
myd6Q4WrlMlthsCKZTYSo0ymv4urFqUfXDIklt3Wy6BIrXHocKUeSo8zpEHW+myL93NkPNsyF2Gm
2j1UKKYV3TBtE/j6SR77ivbJCxZCnN9WpwYABKFPsbFMtm2wREL+ZMLX9ew/NpH09V9rr9/un3Ae
g93ROVNTmImRtFrlD3+hhmDleC2sB17rv8FBFWHa8LITVA7jDqT2QQ4npdFqbM4sbXGb/FYUKD2x
RoBuYGY80yImehy6VhYDXuTcO3wV/jaFqOhRU6aC+weUV2dbRT0vo9dAIA/nMjGHC2kxww+4qipR
CafCOGCBT1XNmnMl2kH225Yi4mAyqDwB3TBFzGaFOWSihulQl1xORWLIoqQVK/cil1kuJt7h5vB0
wxXKwCe7QkEOljefpS5IofihdvUyvx6TnjV/mUPx0YyhrZyg5UHhBMUUYQI/XmeOQ5Pg6zKlybrl
Mjhd8Xu2U/fXgfupVRmYY2bb98R2dxnwRjTKMwptBtS5Egnzyv1h+wDboY2yGNsgcYFHg98lZhFM
YPJW+lncWFOGC3yN1Vy4/+ljpAetwBgjQZV5KEW9LxU7LfUP2o9P9DHxENzH9FNlubDVDbiA90hX
Mv8ZkIPOb7bevPf76a3yB/qT7QEEGkeLU/zbjaWVXeEhBsxJsuotstbt6ipvoqTANEm8UuywSjDb
AIxKGRcNTGSi6GH0XXBcIJnPusBcuVMW3De22O/ku68gPg3C5Nnyx4J5GDO2wq9Kcx00eeqh44t+
pVpUBk8qSnINVj4WESFbEuUf9o6xY5QSTGqORDphpaEaK5t+OthdWqUUakrgBFTmXbWBrkU0tF/4
kxYex3Sz2xL5/wJvu1Qnf8n7yDqHUHa/U0vF3VKuoGyFyYkFqADDQPCLHOHJJXimztYkzrUrnwSY
fIHJzMMVbhXWU+AbjHdutcktqitEDvVRZoSo0DDsJkBbjkhrS/Zim4zq1ctyiy9rsoizgVCQAydd
31N7lCGjULE+k7NV2SI3qRcGZ9STS/83YcV+OReDyINbZYuHx22mCPhHeVXQTGOANmLDZz7spBk6
5E6lAodtORYDZJvDgAGsXGAq+6H1qDFT7nc6h/MkA2g+P0ViUF9lbI0e3VtbsgUnorwizgOJ5Mcr
SzYtdJpedrllVyaJ9BZJ/3VSDp2drznP0fQzkjNgXjpouzXrfvA28AeGr1vJ/lzqqUt40n1oZbjV
NAGSPxSuRYKQvHHB4wtetdon07bjsRHjTfsDcV8mVbmQvq3V7+bM2mocZoiqeGRT/cLuNP4rCJpM
UQ189q1NpQnPPgFUESZI36HZBLSK62rm/247yJx9CTHeur88WVajSgwS36kHodwburNHczhEWYtS
BsUp95ZN/VRWFVgVTtcsAd/rx3QjKP5WuOFYjykXzJlXpXkm76scx78Y4QaqkUyGavlp92Za1/vH
FuQYsTNFjtuNLpaewzM1gQ3snWTdQbUb+HRCQolfR4JfBjhYZhm2pFwUML+fg95oj/xSZx0w19jM
fK/siHY8iWN9rsSNH2fj14fQaHr1ukTpXuDSzKF4B1LXNDaxy8AkLYHJqo6n9/fSbtoVjkbzwKU5
A9BqlSrQB+Em0vD7LYqcVGKRV183t58SmVLJA0Pygy5Qcy8PSAmnPeXBtlUT0RIOdc0MGgN4e+L9
H/Hc2owN1wpMbx7X1qMt2oPcC7uvdD7CAjViqHcC0HPPDnjZNjOPcHwLBbtXbUHxlmG5a4FI0yQ4
heebgL2lVs823IxwgRdZynX3MRBO/o5sRW3GnxwCNg8mHy96T+QsfySUpxooCeyNqgV1k03WlC3X
/fa5bd+CCr/xq+44Q9rlwtKGLcmxlmGaRbcy0pw2dd/j7uhMSFYIKdXW/dpOFCI0MfW35QVwzkqj
8DOdxRHKATnR/STL3wzulR8uBrC212I+h/iWOcUQKnSY9nm53K0OSpIsq3nbNcq8MNXVYj7JaPw+
Xf/sjwQaCcfpC3JU4Fw43JYyCZ1+2qsEBCiVHaR9mRwFar6cX1nyMhIshRmIqAxVQDyTzUj3iFIi
gd2QCOMqT8rTPp+b6RgO3f2PhtFiuaOKQauudAtkwWkjAU0wlx/s2CBwR3w87x7KEHBkfkMBLQvG
99b33k0eZjCnpIWOnRki/mB8L9bShCa+xc/oGi1ZNL3eCaf5O2uysZABJyEw3tap4FQrUBa8PHws
J0YkDaV/UfPrpQfYB2DHwzreJBmVe8kWQgjmdZ55xpqhfNb/RXGWLOOVeOTCfC7iJn50UU5lUFjR
lucKekP6kdYMYU//fpy7M6ltF1jHWkFiN5vRc2ujckWFl21Ib1PQMHisxH6hJn921U/tPbUwf8Kw
5X91G9zRg4mBKAtKym7MBqtDeBO7KuDnrWqo5fwSKBebqUBdcra6f3iDlRJSaA3MaXJqICUkfsbM
WdtOtjVMFjAkWHZX2tGeZDpSmOMN4OfKseXHZKWDynH10nbAqD24cXFGd9zFrl/RuVfoyebaqHEq
uJDuddkMb0aWX32uPd3pq4SUXzjRW9KxqtGB2hPRBBwNuFS1w6NevEcvYQ0goiB8DA3jilIk/2ZO
T0U+AqGxk4Esk72JV4w7w4BpzUlvqg6enWk0kG+lV81rjG9pIdFch2er3ThXiAXu9WcZUbdOwib7
8eCaTnsnEJjIDjOF+2eIVJm6Naiq2G0EanSPhkED60qAkvaY8ZV4J7AD2F7CPnDgOoI+pZIEzYwo
fher8X1a73okXNhgPEieWvEb3hP/aK0kVFaJMG1YdpphympKh/QLlF7WUIMnTP+i5k7rwhgF69AP
aZBZoQTaumgIV0IFT1tMhqDOOrfsbuYA9HDFrqbo4l81vrrOHRHENe5MZchigZLmEhdNRslopzH3
z1vrJYKw/sprx7F2yxiZRr1sZQiXy5c4md4QwTYpzyNsH3dao2LbuM43T3Hwc8lErlcGUT1bLybR
9BG71fW8KU7Civa+ogU8UmpKxoaE05YmatGfZAxaSKjo6cJW1saBgAu/I/MZseQcpeZuIIz8bdHr
uTJ+zjEtZc1Q92SuPVRMTI3LgAlTzwwbr2K3gESZxQ6qbS1pNxRuI+xhxuMI3ajQRoYPjP8AmetV
VBrjGt26lvubR+wUAQuYlXgfbNaWWE5GSueNUQQ+MZOB/RnBmPOaLrtpneEmwBOHtIS33rjKyFG8
lIpRFTlhrH2Sw5SRpocwxSwa3Rw9bnJIU/bxarZsy0bXZpu/GuRKvSw/seUsl4NZD3VX56udAI6P
eP8Qoq2mx1qdfgMgO8azsCR21GiEG1JgcrmGN6Wk5tmDMHi7JlxYF6JcuML+87wNAbaXKa58rHNF
uy+PxNss/jGWlA+1FpPrhbtgNG4XBEJLEPbFv8jqLNi3T/bQJGAbRnJiCwlZbPYS1Qj/TXmypZd+
hp3G/4I1UaYyjl1sJiWCkNpCYk7biB5MDqYHJXOjiORZ9I4Kq9mph/o40Ix71BbTZSqJWjRUIPno
rqTCeoEl2GGNy4eAWjCnTULGDXsJ66tUs0Mbpw8/SAV5L/YgKRdZqHJwtiYEnObIFbo2fmei4yBu
70NLOThvh/NfWEi5+dSVV3D+GjJrLIZo7/0WDWu/jecGMYeOwJoskJHb/9AD7cwcAksucbKCI+on
Pw0DKI6KsRaVFO8LPM2JHCSBC38lUgzJ6xJvj3yvD18r2orDB6Vn7p3YH+BnPpT0gG3H0ScaTZzk
yTWNZbJq0lmMSJAMZmGQDiTOuPvAjBYFyxN/DqbdrppwVoc1PKl7q2OW0975Dhv5mE54emBH9jiZ
rG7S1wutkVFIFGYkXU8m6T8OC8vsGwJlBy5N+oQfZ9NDMlrFnQQHtc4xFXcwOpz2YWmVU9XHcW7s
r8T+IBDfDLnJyXHiODSO6i5nedIGsajgpoVuAjRa8Hs1TK6ZsrSool5C7QH0lNLgN9f+eOQ2WvK7
+4wplthJKyf+FsDkk0NVz2Yp4QrB4YdaliYHFl0Nk8UXxON14RgF26lgebQuWXE93VWnMlLQRRQQ
vggm0JrvyVfERGbeRXMzQ9dku1vhKTKoojZnmT/E0QTPq0qr0drQXYJYGy4hWrtWJBiKPX3ira4c
eCzFrQnLUb1S3m8ExviQUrfC77YFr3qGcUgTf9vUy4l8z+P/pVjQdEVVpmHub1+t6k04CsWZlHjh
euayPlt8EJny7XRM29Xt11pMqv+pqlV7sMrvRrVcM1cInbOA9+ca9/QRbQXQYg9inEqTo1bLufQD
HNczvaxZBB8igmqJTW4vODLlNUhglDhJs0jV87R8s4SDP4KSzxqQ46ydRrrJYmPbjRM+F0jcyixZ
c83TZIFjhF+10vhcI+akWWIOUlNFhvnuyPwHwAjcI6Fb3HNvasIQKtbjLL7ovcGcHZQ/lmEYiyMH
6R9VLKFMYmww3p8G73mIXH++bMjgoCdeE7f30A49PNFo8V8ndCRb9skFh2B7wYa3HTz2QnNKbhJj
6OPZJtiImZ07Wa099PfFgFfZXWI5i4dFoPdNT9xR6HUEwS90ajtwkyLLtynqzGkQua5xcPpgrsM/
QlfavruNzaZA7mOuMfl0xLimFGHf+lFVhkUnhbqyw+/AC4TH0wSZB9eW/89lwarIyeQvsAbnbR55
5oK/u4MM+FO80Upsc5mK4Z27sbrTOGRcgY39Jhf1KL4NirY7ABAKe2Q7F5Nw3kzLBWno9GM89tQj
wUhvcut/L+fZCpBU0VB0RvMNn07ptlFFJP94LRvuTiSRBTXxhtvitCyM70Dnd21PHgCqCqNa5F9q
zbDNkXMFjwWOeaOUJH+eHxNHljdyoBwqBYDNoHxFgZYe+e7NJYeO+3F9ikKWkuScLtQV5R9Pz9aR
5ntjtKQIcq6ntGMG+YiXv22my65hVVgvj1tmDI4IjEtWs54VGFFIDRmCkzdw3hAZ0hLM//ZCsRcf
AOX34Jp5dmHMRH8k/4zJB7nlUuIckcXZSs8I3Jwtwu4SpDmRyt4J4C8MAVWEhLCFfLLDNEzAhN0L
1MPiIFvSw1nvG49k6Sm9L22r52cn8PiPqDM77x1gqKZ6J5UqNMDlkiTufz6cWaBOdY+7A9yuKQmm
gjNCWtL93dQntzxNkPR6O663RKUirg8o+Oo/5wdb33MY/SsvccsJtRfOB9mHj4Uy+ens4R/5X/s0
5WI043aA2E7BZ/+8i5dLvyhjeB0CZwaaUE7Vax78hApVjPBST50ot4FV3SgH/w2E6OCzqLZTpCWj
SRjYYlOxy5boEepbNlIAIoG/Jx+PIPpIadG7gZN/3JzPeMpt8hjmxCVyxBBIbbEVDKaZCRdeKldb
ZuIJA7HSEn70HDG8f6ld6NKcXkXKGs69J0FtGT7I6Obk7IJ/UCwGBcG+Skbbz3eieOezJKDgwL66
pHIKksEcpluyfAOMO26hYXhYPxOM+901XkaAWycg2H4cepgFEn9o23KR7UsV72HeQ7+FgdaGxY2y
Aavoj4+BC+tLEnhPK5yEtqan4fXWctZZ4qaGUqte5vxepT2+HMYUKCz7dt9qcxyyvzuYHAoXau0F
PbPkEHaK2zdbD1lelVuXhokRRIbzgKSF17OkcScFDSV1dcUHhguHfjIK9nBfOsPYJlEEK225+WdW
edmm/f5HEGx6OcdB/EIRErhjRSmmH4XU9o5gF8ztetn7k/MduYYd5tmXwPIvWrBYKvAdVHrUIKOU
JsDbwz7ws0leQoVMtu2xf0HVxbkFZPDrCvq35pqQipi75FvD05vUQUeeydkMT30TlA5F34kJ8v6F
QpZU8tal5BK3qwRkWgJzS7JT8LEczO3xyZ0dYwleVbP0Z86Oywb58tuLz53Bah12vZv3Rq7HI0nL
8n8vD9F8EQsNfR0rRPgKevFKVcz4HgxmoLvWwFTNCe53owdtgNWz7vlRehAKH4QVjJEo9ixa7HcJ
oji8gQKJ2DeoRlmbi17sdmm2wSaQ300/y/Kh3wLRLxNzocu5IFfgW+qIjbQHm+lsiQUb5xJjvAPG
BOP6H6tL4jVw64Yl9sD/NuGg1WVpOM40cnU6ZkoFZr+orZ+z8ASowB2H6Da2saZ8QdN5CspTxFIm
06w7J4oi5/J3Wo25Umf5RBsPvjQ/AkIJHQLO1JXQizqAdF+/3vHqselR1m3ZRK/fkeuoQve8zoN+
g7h6yloEsgB5rjtVuw6n+OLGM0xkQ7pfEsoE7gassNSY++mZP6PJLLxPISrCoK8pfdAM7ySlh7+W
ERO9F8yb8mXSgVbtPzJO0f73Wj1Jnqv0J/prk9qx1PsM3HqhA6ufcPQAhwRY6YkmT22KZfPQtIaY
zWv12R9vfLS0qV5Dic8aSPiXhaWJPHsvKh8E35uCh9g2u67P90XE4gFsRyH8l6febqQNt2v+eNzp
zKz5DZkeGlZdPWzpv/to7mFfY5wYeM5Y2YuA4OmMwBtV7XBflqzr4mDL2nT+ogbXApa9MyCYYL5I
U3SwA5U38EwjaQddJZAySexqUYiZjv2s7hRmomXiellui0T2Nli83+1D0JqkYWuhgOW0mp9eslmn
metIuMUXGZ/nMle4hYh0cwdi4+LCM2n6hTRLvrhIZWquOatbIzU4+MwPb71Zy/lJwEwFq5EJOs8p
u6V3fOX+v42keyPOcA/I4etkbFhsqbsF4dXufbyCw12GYOjcSFMy2cZ1TIp0SusLDLVOItmFSgwy
7gK2Ya3Ua39azkz3Lzr5LwJXWNG/HFHbPj1arkfbd+81Adrh4HBFpu+CCPJlVvPioPrA85Pt+ySL
B7BgSmNBxhw/DPSdUfJKHNDTv88NxednN9dwxCb/BQrDoCrn84+AbbBUgJO55uQdWFl7SOBORyhw
lcuaIcf8W7UQTUJPKfbpOpMc89pY0k+pmHQsQ1XlK7I6kin1tSxvPHQSIhUkQVdcqifYAZwU2Gfg
2S9Hr8k2OEbcFgaeaekqA//pi7cYPYTwoJc4GnrxXy1OQjyQvRvDQ7y1IQVbRVloPMNhjyXBCLhm
546o2BmouhZk5s36UYaPcLwa+InZf7xC8ZdX1soyKNwud3AqLzBUo0szMc9X9bTioGUXfW90CYx5
4gMTKc2RUASpJ7W8ixE3Hs5KITB455e4hP5g9ZfSUmeZgYich/0C2zYveSgSvctBPfTGZHJ2zCqi
mJZ3UzvkO1cHWv6EX848J4V9VRShCdFNNX5KPAeSHgn9YnjwB1aTgWvFcrfObjI7Ly3qt5uw6ARI
drgKgBtPc9yAEg2LC4UA94wckVVRxSVG1lHvKSb5wa0P2+JfedBCGO5Y3kgpO0/BcmB8pGPEyDx6
demaMO5LBMIhBrBhH1J2C0D/gBhWX7L+yZODu3ORhTcRFejIULFvwOv7PNyS5GX5xT69shzi7SX1
sHvBE53AlXQZpSBRGmYdRrELEgAfQpIGBJjIXvVBUbSAXSzDEky97mAJ1xWXtA8RTN3Umjm4a8ko
tArAmIl0XaGiBgzBVBQa0WFQSoKYWgG/2B2NnE7i3vU+SXM8Crm5NCVGyQZ+3qgtFTS/rxV/06Ua
O4ecN4reSpINYBAbl1LtxzKfE3WMymNPQrX1riGh82k0dU4QcctWj3Gkuf5eRMKaJjZxXlSny006
B0SR8yq1Q4AOHJJXiuPG8Np+XaOPGLvgGXcGonGc8mLqXtuzHJsopoPzVKYPDtWsYX9T91LCz2A2
JbZtFJw4xW89I+tktb9b8cr7X2Rs/lQdgIUTjpBg3bCbHHXgfu/VCn7mtVTkMTYZwmH8W4Sc5SUG
nhuUBxrybiMbPu4XvV3B6vne/Y5maJ6t88rSoJVnfbuy98UtlPtalmUAWzFqNAoQxtfQdMbarp7V
RAkUV/sYYgvcyEz4iGLpwSgosp/aJXnv8rrQncsTyu+coG6X9lph8Z/FEXQB/FNZ+oeY2CxGdZLr
NAfuGkw0OpnMytieKtsz9a0mxiV0BU9YDmpVjDTwuC+u7IJuatawAbvpGzKODeNWV1+K44zY3jzl
93muat3LyD8i2YDc1Z6Siny8LBJETfTJC/4uE9F9sMcTJqdEy5pem/KhjG6NoiE0qVLWFef83rWB
m8gPF7HkEmj0eMaqdhYi++G/YZFRSTxm5IcXFjw8NQRx8oklNycSw/47SH58ir6rkffyZxJ5LAaS
dGLV43CfCtKvmeYpQSJULFCjFUQeyodRXyFlCNNHigam/dZ4QWwGlolHL7h/DK3kSkKcl28iUBoS
DQthmzFtJV202iWXcnqUUGoOzFWnJEvGbzn3Dq4AQ2t8mbpLO0eMa+5x1879W9jR/E2oZC3t+c9V
qeT22o24IPlrx9Es/R0WYbpw1d9eGR69mz25MnzJ1nOZQxFtCdf1hkefRPQqtpr8UIKLXD+ffNuZ
KpvsVK/WmBX96r1k0gbuu843EGyKnyqu3ubzAlJb1JCyZ6boQ9mirhH4ddykkFJpLmNcNPncyIVk
hgNC8FR/KZ8LWURK7mnq8TTPO5uVly/+bw54B9iucCsM+Ls9MjiRV36fywk+5gXzxcuVfLcV2n1S
vXaS4LEyMfw6iDQzpfCwJxyrR/HYhiHXHN1ANnfvkm7bAph87kNkMtnWWpjfrjHpD0xHmNjk9DVu
uqlCLeVBnhRtq1puAAsgAmTy/R/szlgsjcgLxfzxAjNswmouod0tay1SEEMWaImZ0gp77nTi+yCg
GNoHATC5QIA92FBv3LUMadChP9dECTi48FaWwinfZBKDzhh9I3TFsHcpd55ks4YMUAIdlKidb5UB
EK2tCzb/RpDWWvRMkgDiXvhG4bc86ty9fQAP2oDUaQJJRdE7e9fR4iqGDhwMf2DyW5U943ScZ4hO
soGbYU9PPGQaScvB2HNVuO3OYiF4Xngz1H5hIRP047vGVHjjLehOsNgTpfF2EIDzKb+on81rpWe+
O9TMfzxaBOiTDMfsOXLIyOqEO5ZaEkjnDQjVqAnNMF5g9gdLTAgfQXxpsRdA52oTrf0UpXrkysrB
JOkq5blDY/qS3cSUC9JhfX2xMFwXS2SiNqsfpGdMR34LAa9d9tKxLhnS9aRLmgUP9oCcMa8qz7jW
CLYUSTPip7lWTGwjw+61JAxss+Hk1b4C5HRMRXR6S4BD0PboDegY/1QSGJt0pUNnLr56xVmAV2Jp
1IjKlLLTwGLigXeD2u4cI1r8zHIfNxEe8mvKawAt05ZG9iPWGZNGO6n0B+boTV+0jKGQgQdZn/UU
cNRtpfR4ERoU4X6KB//mTvqw+muh0s1v7CtJBNYYVOtOGDrZ1xUkdv2GpvBvbNsini+3QTHocNVA
4iSUaNEZuxI9AkW12eslCvXmvNAWRgNBwzF5+ZzDoT/jE3FxFdrXYECvaGwLThY2YO5/1IO/ykJ9
8nNZRgfzabLx92cxMMFj2pq8tj0gh3hj1yJjzn3iQnQDDBrS0CthlVZEqz07GkBeldyLTdskn6h2
Ncr/3glw+vUNCyw5eay8TGZTZaiTs0BWeVRN9eyDdRHU86CxUZpl0J2G4ADVxb9i2dyiJiDS0EKU
v9XlJ4axDjcuw7mJdvgP9uXh0nTXVfMjfWLQYkXUt7aNCtU8aCCoA2tM9IdtCbt3VStNptNKDLY8
0r7UYlhBC0hK63Q/m0JdtwH0jlSFzxiC9BxTP/eAmoF/P838H7u5WRfjUGFiUXiEIo2Yjx2pVJhn
Z4Xr0vyjw8e945XXfXZZmU4nmiT17Ky4x8drstXbD8Q3yQWcRtgmrbaMMLuiGmKlAdXLtQ+pS3Cl
WtafjvjoVBqVG9ocaDHmQpsc4rx5nsS/5hItps2Yk9Xw6MsTkdArGVlhoiSB724T2I7qCBHRohn0
lKqmdTLZGlLHsyzJdfCtWYe+3a9guT887hSOyWPaYfDHyAruMP+5fLBWNqQVFU+LPxdWf7UyjH6z
L31N8TNfqnAQdanlPbiWZeDY8T8X0qq9N2Gvw7GOXBSt0xO3VIEqYixLu3hxCtELjRJbUYC7qJhJ
ITj1Aezhr3Ok+oKk9Swabq/hWlskGfkDPK3pr6soalRa6zN+C0oDA6fdH8d8Tgw5ICQ7MQuoGOwl
B9SNH9LdM+f8CDB6HNDynvtUChvGydHiG5zmAwewX5AOHEYbhoKCyeGioSnhqeF9dHD5TDQMWpet
IKpHY3H1kimKU+ptjV5sFTp4h76qXLBXwTm9dzL4BUBHs5CBoyuHjlG5xGWJFdRb9FZw5UjTAF+y
jEyQOcWtlS4/gt2knTtjPU386gWfk8RHbvJrQDp3LYlXhezkW1Di5OMiI9+jNQmYIh08br6uAUW/
F6kcZuWMa03GyQo+oUPWkIE3p7+Tb66hN/BWGEBLswcbA+QT+ZZxm6G3Jzx40JBLtzF691yJMaxc
vrZ2nLwd+q7IIvOtXBavbLuhENlNPkEnSM9MnbbYu95ZM6yJHSWpq5tux1OZftf0kXH4bwnvOo9R
juEeZ+qRW5lHKdm2kuzXxvkSrj6kBiWrzrZAaRTWX9NbxjHZwrHIR2ppM6o+X4EjN/7/THd0c+pF
kt6s2sQCqTNU6BPH8abXG5MWECOlxm7Px8MiOGhxgP58mHSnG2piGv/c6KQAX/nwfsolT/1cDo01
YqcjWPdUgGAJa4eXWVpXDckRJVfvWZr5cprRGGAghLLIGsds9+2n1aOiYB8MJXmL0x9cv3cZ/47j
+HNQ4UvgDflQyUbVZRVgq8p3Kg4Nf+1CBkWXTw1aCe6MzQmdd3TDpenMiOAzjxqqP8v8ga1PpITH
kZK9iJHVBJO/GSYap76BWLofTZU3bvbcOJzvuwF54AY4XNb8ARmevcnoIIyZCDE1XyHlSkAJRi5p
hEnuADhyG+rgmKGIxpL0+Ydz2nf3nTselLBjgcyhoA8ZOANDyc/788GxBjWY/7XnlOFFQpbj69JN
kkVnc/fJPUFWFdRIWXZ2OEYxXosrIVtFSduI9GcAfurDgrrGRBf6lxEAt94AwG4Q49pxVL0DppXU
0zOyOdkr+tzZtnDKAS1wE2fkBu1aCfnaGSwBw05AcO/u8OY5oNgGrMNRm1NDCOR5K4amANmsJN+Q
p3k/ZADF5FD95NP6LQu3VLyqZPVgU7f+YnI0w7edVReg5q+cVnD2KKvL0OYb/F1EzQtFs5leABEe
LmeEZ+9d4YODdRiA0qkIHCoLN3Gnl9MMNp5X0U0ewOGjFZEBkV25QOJII6uMEFHVqwueMnWeYczK
pm2U5EiAtpA27Q05vY6U0P54ch4VKij1LoyrHbvHdHpJN0ftW3rEagBNeNEF52aBCyVkyiNCjYOd
C57CpgB56VjqkcMvUdgp5yEwb8vDVjmWYBnBOZlSuPwSK//JIV/XyajWrQqIlYf+kpvviWZYR2q7
vORgQc9xUCuf5xp9g0wCG8j3IHXbrQq8qLx3R0mwmQZLMcXr/tESBdhRSG0+wU+rlSRzC3GabxSP
YDgipi1M3yfd7zyZQW8Wl7Yv+TtnHHEQQdlCvN/OgQnb+z4ARDxOjqygSlcscfLDZfQ/zjs9vfzs
bXLB/CQRVDB0WoBLhOrepctKq32FlJKB/4LBjs2lC2QOHxgwlFpcey4ek81k6+7E3XccRJ0HDobo
c030+7hLKYzPF4kNRu3MCHWD0Kgx96V0yGoIqsfwFTeHdNEumOpAV50jdGZGNrfJ5Y5w1Q44CaQ7
LfovUmkK5nlUZ9RWffYsVKAapeixweG1puIXTD3+6u1278iP/0V3VQCMZlPrcIEDgVZ+KBzv1pks
58hSWFjjo+GDlQKuaSssyNtG7PlCtxzZirNerAWUCTPQAiDwnethoWlBd68DBVM5SzGzYx2WGtYH
d3/FfdSYyUXutdEyglDY/k9WO5GUkPXXA16OOQuCOowOe4iMx7q8HngRNVWFvrhS2zngurDZDBD8
0YEhiS3iAPpwOkCAE+ws0tPQRaIxcnfBeShJZ6C+wzbXD97+SwUyHdW56WrZ4W6qI1PW0DeDFo3j
LgtFA4ECBPIpED74lBZOu+HdiO1bxeEspie2V6XGA/WEM8Hv0ARyqQUrwICiHErDUMqVvzfZjyDQ
cFwp6KUz7Q0vxzTcY7WBGu8f+WQTQXALe8l17302k6Ewq4DKOLz0Qv8g1nQ0nxOi/2ymGkOdyzqd
GYqEHPFs5YsxnLlYhMSJgum1nOHRVQsQRLA/46RAkWfMpPUvHeV6+K6bE4tAZligvGUYQYPtgwIt
gSk7BS744UpNR0+ydGqqxu2ZhWK6KcpPhtzL4lbn0sXHuQz89gyPX58MUcsEJxkSe9t8WskRoQ/R
jn3se2aUSbtZeY8GN+thoMBFNKBptCHAdV8swWZ7Rle/9qf1HqwKwO0gXLKba4hsVRmKTlsiokkw
Z+6O7KeLkPiVSGcesCEvyopxWPXejuTEHjYagA6Abf3WET9KmTcV0CH5DRAldY8pAGMHXcLcN62+
YiLE6fnjIeAA2VGTQMxzErGILZs1/UScj/pSq+I5nfA+zq+ToaE/AImWb9xm67u2sN33X8qRchcl
2Gj3KXIyE1JRuP9gQR5+SdyjSXqVkHhKFMhcr7EbahpA4yTuq+YKrbICsBPggeq4lyzmCrkiFyag
Y4wfnG3oWHDNDI2U1a3A88eAmLRv1ElBCRUdXNCe9RzhycOeZIbyHyzl/sLsRf7yySWvYU1KtSZA
nunsFI4sYkSFzAgcOHpKKPIMptnEz+/aOUEIjrp9q/V80epM3KjWCMMR/h7mtvFTQl8fyhYSRyGG
9scP+sORbYcKE4Iqg34HUJ5n/vepIXm37/5re3Y0d4kkGwbyQqpmlFNQ5bxlaXmqPuvyHeTaWmtD
lGqerhrjdnQ12o80lUyImYBPphRCekh8OJpq51m79IUfNBfdnIi4OuEjRj4pt4jyzopMEmZwpuFP
khggDyuG/3tAVVZ9NTOEnFljY/7BhzNwYF+0JMfT+VJphRpAGc+dt59d6xHwb6cMqOTZEU9iZIaQ
cQ/54rfsaP6GLL23aIvkY0XwlD/gb2lroKI/o9xV+vyre0jNq/8O7yGxW5yueVKnl76Jv42QV3a9
gRYHJH/twFIaAj5LcO7pmBHMGhHbluFB6BZ7BoV/pDWxAwfhf7YknzeDbZJ2lKdxGRAd8r4/cPmb
UbrSAUtWDuQZfKQjxHRPdYF/fMKSS38zYSC/DSITu6WzQ/NM9E/f82qogjtA/VMdG2v/h5lnN2IA
3O6ANgBcl+msemBortNTB9sxw6qJxe9Oy+xKd7ZkPBnpwwtxPPJwBb3riZWn6vmRbKCf7SPOK3KP
p8kR1vVN14MK3gdzzqyadq0zAmBuhi7lFpix15ia6XPAu4RPh70CJoNtrOBnLpRZZm2Vi9Sl8IgU
U8XOUtriXqSp5vnWtNhp0dUNxOuNBvAmSn6Vnip+ufH9IqEl+betxRrgQeKQpZaDiRC2uqfoVupd
TvnA7pnA8MgS9daimwLuCu41iBsRYTWO9x+zskdhw1tCo/PdEXpk9SzIKwHtfm4eTcP/0uEb3+R+
JqPkXJI517EmIdjDvbYpt+2kjx9sPjK9eCxrISujXygsD57AISI8ilfuZoRB5x4fkVppBM1K2JTX
00KTrXYgLuoj4hbJ0qbmtGOH1RBRkOhBcWeoCkl3rlV1Qw7t7qamheaWFFPp3fKzGzxFPaf/y+mw
i6hRS72Lo84RqlUPAVD+e5ugeJ5RNjLc9J7LOS6zZV1E7+u1hu03RHEM2ZgQuQCNJC5sUSMCw0nF
9h2YM/AnZCUni5YQQemaoNa318zg+xSjz088hu+aTvXhyEFcHdT6Q4DrJ5yuQLQL4u6vUVJXpweC
x7YMOyvlip6fJzESZZRBOVtOhVeLh7ncjtDv6ciUmsXqwQQKaUotwIjLqjDjmAVj58Fz9FJRWyZb
t74tgiLj9A+UzeSUQTmRkCb3DfuDWzjGWMgfqV/RaV27er2RWEm9h7EpliQI8TsGnzB1eecK6tS8
WmwHN3m1HMVN1uq7NG+s4B6PvA+2IZmhPCfP2s+tyvIOGIOV9fc2Mmy0ABVynyXrF0um/mY9bKVM
900xFjHDGlCCyBkDESBG7LWjT3wBt3wRenUCA9DlJHTNu1SOx03xQ0t2oO9SBves5GqtEJoajU4p
GeTK1Pqdz111mN6Ol219Hl+gd+gE1tkZn0RlTiX9sfsuu5QXSIY2E5jiWdyoFtJH3LxnUrzgRQeZ
KCyTs8Qm0ygrCn7b8Xg5+eLvoACvRnhwyR8ticASUwS3I/Vh7JCuDh0fEojNOfB/YJ4Tuvow4STe
ADdyL2C6IUFBVV9EAo98Sk3dzWQfG/6Gguj7xeRWlBmZnO6seVQwxJrQJjGmoFKUaNF+8QrJmLVz
QV4oUiu1QFmigM8z4bbUtHpwBGJqnjTKPd0+tn7S6Wc0rWdb7mR+iZzgQvwY0w1vrPOwGdXuWEwf
nsVeVXnpMBjXmrsdfLTMYmDQYz+kPjIb7i4ENBe51Dr4aKkNtqlR3y0jtbGjvtMADIxNLmxmFfa7
Jpethhn6nimZ4S+kQWw+7Akoo5JApOeTyKVHSh1bR2iNWkctIMByTn/rA534ryeMFi0I7ZELbFls
vyLDPe7FHL8gli9RgkllU4z9x+Hj4+jbyQX3WGNQi8MICkW7Z7X7gh58q7Rl5YysIHAWMEY9iN16
w7/3F/+bhBoOjIWqs3TTFcIGwefXUhhz8FVJuiky0KzMLTcXC9wWgTdXwQZc5W9zkUGTznkVBbZU
9H/WfjARIG3OwDw/muuz0v8SG4wvSfVwBY7ldFE0otK/iCPka8MNaOzfGT94hOzRfwxgwhimjghE
ZepP0RQthdYNsl2xdy+IP0afhksfAdEOBBu0UP2PJcGXfDNJiXcRXnpVVd+FYok3QvSGMiRp9OYl
DvWxm1Iv2QqqlTbK37U1MoDRuNtRMEzb/fGHqM0QYK4IS6NM1GxKwKPcIP/C0hUcDNfWWXSwCfEt
zCyY221wDi9siW90beLVGiP5u9iK2AuELibcCNV8rRq+i/x6L+R//Bs42GUSuDL61AbddoBII0XW
6hKUG2h/whp+PnjA3ppJ3d2gGaV86GDrCZB6ZFSdYxAgYXUOJmJmE2psbU24FTaXs1+LZe5O2gZN
t08fRRKdDvIs9tB/0cKSkKLeADD4fDSQGMnjV9FBsxqUakslzpaAwTubuEoETk2pLnWLMvJweMz6
+PLXzpG6c/8I6Z+EDTp8tSQmGaaLPLLGQKlnCHMAxEZAgw8plDqgRWkDoK8v8qzMOwBN9yYFDUor
8fI29j22VFa72jR4q3rumf/+WyPTV83wqSGKXxKG28O8sJY6txXTBgMuSAmqcWF1o5re2of4A/9d
WXNX/9XiNCbRjcAQZ02iQCS+aICJo+gOqMHaV6HO69Y6JKvGAE72wUQtQkf9JyZdqYf4vwKR/nnB
T6tQyug58aR54TEzPUE0/iH/FNHZMvUjIdhJc5UvxIjkgzxvxiFpdUxJvlOhj1pFFOCPJ+czEjd0
4XxP57DbHqg13bu0uLw6SQJ3gepOAkUJGs/pLg7d6Y7eWCx9MdK8uBgQsxh3M8w/fd+Y5UmLcYLF
hOP8cVn3YyqCoCyvCm3WLRoIW6TH1ZkJRfIVIXu27NuaMAFYxwXMv98Nk+98aN6kBKLeHKmzrQaF
7n25031fY8V6+d44FcsxnSCUqNjwERNWHtJl1Tzq0/SrhrGk87XE6Ywv1yy37nbGTohQ8McoYYBw
cHoabbeV4osK3XB9lnQbNDvMVDvquAJ99ntNfVLB+V9xSR4GpfYyJ5Nc+jOV4mc+uM4e2Xrhga9c
FID+Oa19aQOGEer8YZ7Y4PiBpxMBVfFM+ljzEInuw/TKSJR4hOfwnhpNuCwFjM35LmKe0qy0iCdd
8nrMqafhBOTjhExWFoCLWOKCbhvFlixtkePhYpWTjytYGkkzXTqw9iLsWFf5Ew7rMdbDWP2ey0Yg
pRnf1Zkl+KlR/wb+Bc2FTs0ziFD/3upwVIacBqD1EZCoMfQcWCyuJhZ6ZDAN8jP6MQduusHI9yxq
VvgZjR0xG5pDENJHZyukMcZ3X/XTOUQ0SkFVrZmwKELIMD2ZV5orQd4s3C31XOeU3C3yi95k8Z7B
1fOj0zbrM3US+Mfy/RTYclsdH5DRB71VmVrf3K78j9OphHGl3ap2u9vyZuAvN8wIogL01P5vPF7o
WE9UQh5ZTxf21M0+C+T1jjALYdpPXQQ8f6zzEMmAIRE9+TCxH4KupDtUa+UPajz/TSLoR8v/Z9fh
RmhubSKepsDYvzlOBlCjxuh5ioXgSpowPktKP3fpUBuiNcPUoS98oB9fPJ5LNzCPd2o+OWeAlrEg
vzGJTwmvYPSsO6qpSBmj+VNgdwxR3h6w5OpwI78ZN6oxN5Yqt08UTslVOfot+sDZwu/W/HmMo+1/
cU/mYNDFnbp5dvWDRUvhz29D6ypQzx1Btq3dGkT8LFVgNBgb9oW/BQyY4SXNxqdlZmFm44+FKR9Y
a7XV7ALkifBcGS9EWxt1szq2lywAOdbZZlybptEeOPE+nFKpOR49gy/tjz6fEDT3npa4JuNmKwLa
B1oWBP5fBdTl/ZhJY24z7ZMzQQHwJAtmR/b6DqMoPU1+avVaJ/yjIY7+ZCIUq4j4+Ht5VopoQ1Yh
90W9RkRE2QUCTpzkFYz22wYpOe8ECnoVXDEzc4TXO2Kqdaqvr+bfx1GjfUmZyf9ae/Y9Eh45mEaS
FecwXLu5uZt/Zb1bTsQ2iVeH3TD/4IBANifD/tEuRwFhAA4IoP08g2XVVXUXOCM+RRGswv1YRbuA
ySkbvTB0TeM4IA7/AuE1Py1/vENAZndtw8xv6osNwkoD05BDomd3ADUBCV1QNEpcyhcSQ/kLgazN
T+VWupxncxNCYclGcNDuyO60/UWFfx0oiqN7FBU05uFsLt5zfrZdOpi3c3cbDVizOK1AgydphWtD
oh3ATH8bmIYCSMO4hq4wcwhksCrVa5yrdSuNlXUNpkj2QYP+rajOefKj2wEiYzOlS2dEZ+inWh+s
Hmh81EipvWYt7OccEwxXy5sZ9rKYKhGhF+5dUpLqGdQCugE8XvBfs76dRf9PjhC4Xd4SMngixNc2
R/ZlSiJH3H1kBdEPfANbcJBIYASEarqyKpXyg+m5C0VQqNdFdAWAu9dx5YSwKW60k4O3oABsPXcW
gjZKMHQ/HJpuVishPy6vrEE7h9SYJRP4fTVyhwvwwDjQTQBFSYotPyDC8bxlOWY0tugNzhbGfxww
VbTRhGypcU9JsYzfDawKJRqAe5qjHEc8MI4075QV772Wml9jlSm4AO5D4Z1z3MeghQuDUV+uuGwo
NQD4KOCvW01AFcMHiEbn+YcDGWEGlW0dTaShrd4pCX0KJOYdjASXBwQRQsgWUtDMABHcvH1j8jPX
Oh9Ilt3bAMsmjMQm1kMc2QYNzBu8zY6fn08tU1EiuJ72CzL7e9SuIhh7qrKIvyzh7ZzcbkesxHBA
vy1PcnntyFoIsswa+RM4Wsqe8JKjBDlVwBXGnTTctHWJ62BenP/+Coye0hLlVw5r12m1c2jL+Xnp
TvX4gLygJMptIzeVPRPhk/90BJdAdfqgGWgr9HAHffZmJ1GnI8X6vSLcnc5Rre1f3g8WSHPmXwk1
gexWS3E2BTka7rmmcu/dKjrQMIN4pe79EGIE5u7vJ7v1p+OjDnlEEOTsuqt9cnJZCu/sxLTHxNpu
VZt9Khc6jsu9SdNU0DTy23U/NkA6LFwbFZ7uPxDJtx0vnRrm7kuFvnRrK9tMsGMqEuzTLrR/MTb8
rLngowkiljzI70XvMIC42dRL2RV+AeVmWzU3Ob0t3npIYv909SdmpFUS+kbjCMsdt0gI8IhhEAQv
516MUZtwS+lOeW0827ZRyvFTjyhsD50azYifAzglz6+WOCVXaDA82GEFGdHo+3IbCyIpGU4QzHG8
x17iayrWXvkm7c/cmHca5H+xvOk5hbx+uOYxO/9qirv3vjsYOA0cAUDwkDceP9kozIo2nhG4HZ19
XEpQJNRgyx0LUnXvlrG2PTqriRJKIMkFdbkDNnL+hR9TUjHdsJMx0oqAM3JVQSg5nUh7qorysVNt
+cB/kwIPwEwX5A2OhzX3mdIwRlKBkhMKIBpZVVAvDtOXG+xrADAGGNX9FYS4YtNJnDu3jhJArbjC
8Ds27W2wLoDb1MpSm/GMwLhY4xfR1DPQvZHoe8JsV3PyGp8biq3We8BXr/PUWLuRK0YRd41tfwkI
S6E6hqXb/ouTqyAkoia3G9EaxDw0NfsKWaZQ2HCemnRwgyEKuATilNpY9yE5k2Vfg36831p/BBT7
WHOTOfcSRJfSJH5NDYfdkCfvDDWiYU3AwD8P0OoKZ/yl/7edDkADViT+rJrIXkFAgPMjWVRPpBMe
f+ZrZRrcSWmI9bIJYTvCe24nGxbJ0qhRDeK/o+jaGWhB86LGvI2ygFZxskK3wDOSd6MH21eSNDZK
SQYLgOu48API9UqAJ+evn6PJCdRe1y+vgpy7wkVdg6qVZKBOsve07foowwDpqX4N9yFAP3+mSpWw
dshO8eGeKutS8q1290KDlvIxRDtERnkRnEMOicgPH2TAyIbk9W1XftHgU1E/4eT9PyaMM1LZRVqn
9c3LdrYcWoN1KBhTc1mUsTdhK85OVuqzWVA0ddW1unRnhudUmkQT1drDaO6J0o7Exhq5cJR5385q
y5vRN4Br9GylWwiiI/Ec4Z2Ar4BNMgkgltiz0b3EIkNBaLE3BeoeaFc+q7EDJRLdWUHMDqPfz0Pa
H4tUQ+a0vKVnmXfWZyXXy8uph98sCsHvcHy4xfZwYlDKwy52Lkb9tFO0lFaREQN89xEHMY7hysr7
0wvzHaMUzXyRDOTlzNaXtNvNAjqBjIPxRgOHvNJOmQbYgXD5D96m51ONA7cpVoUyAawTlN1FCymk
t0Ec2vRVkLLlNYXV4EJZSaXjtwFHZmHxdFaWpGjmKrZK1lzmevV9bAN5y4N+dkwyaiV9Afa80y7O
CwIGQfRG+H1iHW1HN9UIe8p0KwhPt50FLnsX2VpQlyseX0dzcGA9ULvNGpoMDRHSeSX1MQ5gh+4h
zTiDM9QTiaOWcFPnRWazPd8NRuXDYrhOAU2ciwnPt8o29Ey4emheMvvrroj/v9EePmd/1ApaVnKp
BZMC0WOMbPHvypRROIiOwzSXCgKpbWDrRREwmLzaoJSZOR333fKjavg1wdfna5KEc6cTl4WlHjkF
i0yiJgGQMSsjuJg2wJg6hcslfMHUHCo/ZIqOcudFG4rj1hN+PTmNte7GG680CDgoHCi5vwR/ma6i
yS28h3hc75KfozNqCIW9GtEXpv08wFfggvc+nCBdCpE0G5mztQIE07iAfA2AJQ60ZMzDhejsVEbE
EJ3/lcNZ7dLKprhlePi75fmMnMMp1Cf0kJjmHE+3KgIvcPk51Cf6wYp8RsULZp2ylQPCNscUWB6c
/x44YAp9i35670GjSyQ/9bzpUeTdmbML7fNXNIiX20lBYGXFfZfUZerwNP6haS6OR9/rK3Ysz8Cg
dBmnzJqT5ZzPgxSA5/7lKMy97OK5KIFfF2CiS2Na5JLkwFCH4CQ4fSUx+jwgIaJmYiqJsnXvSzIC
/ThXm+GeAxCkuZqk8jdMkJcFFq4lccIGGClYqTJur8jaszcvnOslPMbUDF8ilY+Aev9s8FDwF4ew
cnNkB8ncagKM8OXQ4P8+p+j16b8LhHuOilnpEYsNUipOm5IsuR3hrOqehreiUwn4Z6s1HH0M1cER
SaJ+9k09XgjUzNSmF+JmaGbv7k21Bumt1QHtHV6p+v1Gmf8mIPOgslOuWmzC2KxVg5gAjACr9zfF
SI+W0kop5h3yot/CYoH2mRqj0ibl4FbVCZBhOrizTG57vhLnzVkXFcXmNsOsT5ISc/tt0JjWJq0U
UzK5cOLckZgFS2R4MmWXeMHGheDppWkQC+sRFiFSH0oRaJ/kzdSMMl6fHreSqSzd/Rja2PYCePVO
TOvr8VCXbF4LQLf5BHs3H3hVL2t0yjuYKLcv2Gu5Gt84z7RwzMVPoeM6ztQLktc62izB6Klu0Myf
0ehgSe0N1nYPlc4I3KBHTh3EAjEmxZP1juxoagmP1Fe0wH2cXV0r3DK9bz964Bn7c9IWbWGGX3Ex
mNe+64b+qNdMbtZtdO9zW+gYr802d8ZlBoa21mdFQFpH1gfMK7Bu3OeNHtAwKFegPGTHBp0RWMbz
X1Sz6ZBVxQLSanWqgxNobcC/e43WYz2u3JHjjCs5dz84Tsg6PwEVeRd+LwaUSywmexyQrMffchVN
ISxxKGP7Ve0yMmknG9pGwKo42put2zQ4UahE7Y6q2HqYzIBRulfxWPixsmOtcHNAUCw/tVlsR932
uAFCojrrNyDtwG9oht7T4fzs/Gm4T8Sj7J+cS59EdDp+DBGMxMBrxOfNMEizSREehOuqc7uToags
QF3IyuSmroFHR3Vqlihzib5nNkfjZOzHhLlczhhwief2QIE628Zfo7B5nlHrze4pQh765EbxiO2U
sK7XDKYtFbeDJ2hN8siHwDvIUP1QjM5KmjTV8Jod9AbjSiIJw2pySoxhf41BB2LWbLW4AaXGa2ni
ctA4eXjjjtI/zfHP7caKtQW/U6Nu+y5cKgJpg3DFR0TH7yUTg2LRZPZF+dOzOEXDkjQRWJ4mwo/e
NQzOnynGsqJ1h1/PksSlliI+egRn1EmB/W2oRl1pazhciHeMEZoToFEn5geNLpZHjYxuTwhV47On
YjwIVxBJE8KNgUKhkRVoMXGVy0t9lXLqVZRXRyacaiwbqzRS0qrC+iJnoTZN1/UtETWrKnr4n2Vb
0joWfYRs9GL24rd6yQbEumD9FPTTvjQ/lNGnbzy9KN659lquc/ZATVw7vIH9it7BEaHNuchHAMhA
jW6H6Jy8ZViu6DiR0drUlQsNBJM6CKIMicGdxGqxUT/WGXXkqyT6v4sUpCknbRvBbIqOky8W7wEU
hqTKNGs6aApc77KhCLUD8rvbvMyO6B3jvfNVrysLd7/AWiM2a/FRJtwTpxiDmMB6x+tywDycC0fY
u1I2WAzAEsoG6jhfuxt+IN/JZZKZWhawm7dKspOzSzzqbPW8FkFHkJfj+JEGXaBpWPaJZ3tPKlSP
jXuU4GBMbkeOzka7y81UWio70rr7wy47gEVhfGCF5cOyThs1s2ehfTySFdDbbj+8izfJddejVcWO
Raopm/ky/bmi4kRswNxvIGYfbwNsWO3u7Xu5jbQl2ig6avklnXR1dLBn8xLepv2NvT2uJLS2LQf1
F49ThkgUfhgGjy4lJ0FB45wTR181dL6qlgfBmQEnYo5Lx9aAaxHARrYiGO1p5lTSLFAsgGYqcp1R
6AmV0/eBBs+Ms57omjm+uonXKmuH9fLAcXeBrMiuorIs1L7uvlBJjor0wR0jg2mxdJmvnFX366Wh
+J+6bJQzrKy+LDnZ3aSYTISTbOPHowZpMzjLqdEgAN5GoHSwRwIlbheQzkEr3SoCqPmcam5QlIHj
B5qi3CnMx1SlWHzMQhnsM6pTn40/HlyupwHzlvGADble9iV2lCquM7kxKXIQQPyhDWTYouWL/UPV
3KKelbxiRCAN18L1L9AmABrd0Uc/Os2kmdeZhlTWqKPUOicX+c3DWH6hOdjQ/uXF3Ybdm8Mqv/lV
xCBjtwmLhmkyMFxHZWgbETGbKEWgNc2DVcsvAonFwMdxfzl9+86IMjGFsRzeoQ7YUBASDd6kngqG
OlWKIPpXPClqvAW93KGcNHfJ4zna4r75TtBJYN8I4StKLvHp5oF7imnaw2X9Lm7gpvd/UWfko0vr
qZUgbOMdfjMjtXK8Ak0fLTUhLAv6nwBZg7fRvsI2jvZCx0tWeJkzYTTi4vL0aClGLkRAkhEmNKcj
YePv5sdD51qJ7iAdnIcHYy35ez8iGHHyVpVYwPxjbwSIMAazgmGVV/D0GD+V2wHfDPGsWuLHFYmd
7Gor2+fent6/YAXCYihNsC8dI5NwTorXWxl5C8HX2gZDvKDFq8TtfUtjUcBM9gRf0QxV4He/Uz1a
TsbKm2G9+Xm+v3tcAv6RriiTFJa+aHYPseEBg2yh95BQv6WUP61LMDD+mKQWsavMy1WoFxQv43Xv
TId667+s+Q0Kwcs11zijUcZb0XPcpQEXwTt6FL+OKUxE5mKL3GRRVwU5D1NdszPF8to2zlzT1CTr
aqYWTljmZHF7XB1OJ/8O2vZ3ykMIRhmKczcjdpCtvIh4/elridwHg5vqTV/2PWz2oATxz6X7gRTK
2sIt7QWIry+CRrAlyxu5j/5FJyRqlr0sbYnrNxAjupvUGd10hPhsxTHJmABzeXYnHTBXz2ZUlaKw
KAH/7mOOXZ08dsls06Y5bC7i1rZMlKKOYs+yTvTUzsH+NY2/3tKeZ6SRbhlG9BBTgHrUpNSTLick
0ptHH3USw++uIMx6KfmCkGHEaNPQ0TMU2HpwPts3G1lHGWdIASKVMTOVMxRc58D53xdRH0lwvz/7
UXBivDTRQxq6roKParfGRniX1i7aUpRY8NxVqW6I/ZLs7dEYKa04BFdgJBaW3IW2tJfpKBiJnNcl
KxUy/6EKNlOQirlBeJFvFARBOlVKpY3/JG9/Z1OnZ02/cV13Ah16N/j/Opr5zSVEr/X+Dn75TbBy
dVHYQKBb5dXxtz7foBFYI4laf9z8v6dJYwe5n6oN7a6II09qTOmKpFWo1GvkbmDaaa02JhWpNVTe
SCTU2PD82ANEFpFAO/kdepmpgxuaQ5awB95XzDMXHE7+x24bdandY3lJzjGMDh2uQwmyeiJmEcHH
iPfV5LyE3rx1jjuqSBglgDweq/xAjV7CER31d4lG46PoZJJddetfO9XfWy6trEzuMRzmZiABlSiY
OOdtQWILb/rD7V0UsngLmV8OZ6l2MN0nyHAFo8001alqDMWRb4n6kwnPc7iiUmB+mk0OHcVMZdFq
alh2zK9mYufAyaX8y8id37ZP44m5WRNdJS4hX0Az9owLZUzGmM6Hsy7AJi+3g2YUIW1H0pdRcEH8
94Ds5aSKvKOXG+bit5ii256vz7anxB//qtCFMmVzh7Sq53T0hiv+PbWDJ4kxfA3RnlYnkA9Vdek0
Dn5qocJwlNgG0Yvo71hkuLZSzuGbmsmyEvV01XVra7eLQRrsqzZX1lfDW0O56QrCKgJosY3+aScV
JuO98PcqD9Y8eONLRSBCGnAvOUz4QJ95ABUg6hKLnUkGrjm4mWg/DCbqsy+ZwuQE7eGvuHwrYzIm
kPaLjbcMWa94WBqBz+/N09DzpQlq25FUuxP2fCVD/7BCZ3JL6xUZjuCpssa8+vQrF1utPfKERfiQ
WykTc+SmIoutDgaM3lYdgPKG3dadKWoJkHtadD5tL+6TOZS/r00xI8nyczWh4+0oW2FGf96pKOp9
KfCTY6/xsyjIjwYjixMOoTaz8UbjmyMgJj/nXuI8uLTkZug0NrrVaYfS5UK8l/+rzCZDND7jbLzb
CC9blWrWSauCOkVy9drPn2SnFJnPHhf4UrkD6YJTBD+FrUwa4pvFxbVTbI5CDdCHLsrcjKD0gU3/
uhFghQ3aYTRPtG/t4JZRqwi8j5pj4y/n/0J6TZ3IUlUjVK2QO82dcbcXCZTdPipYd/gmEBP9z+hy
18RX5Ol2jAzM5CZd5C0aohHYUzsZMwdFkjAXIDcChgI5oDcEZWoPZ+MXmfrDUEEIKG+/+L16/O0n
M3ZrRRg0XjqbWlhzba0NvDJNLVv9yFunVtxQEQH4UrnuyOdUn0s/4YhuFgr1bI/JkbUzBw/C/9y7
XSFbcLRFN+GUMmHQk4Vilgj40K4OUuFoZGR/qtGIpSjYet6Y0BBwQAOt+YqVcIBsFte/wGaExx1K
xpXy9G0YRozlJZE0zCVZsIZOZTXEr9sYjVC0GG3iQgOrnZo2GaTW/oT/A6NtlgJY/O9eNqzMcU9x
qho6GuQrqbqfihpqdim9ng5M92mapeTOqJua5PfW0skQqHuwWBA9aJ441DVx44rSf+aoFziVYQ5e
t0s4XjNwM2jT1g5jcwfDFWE4+FgqLu3LRRfzNWUMlT3SImsWL48t2GFX5phvclHke2ArbR+A499L
Y/zNqEFYEgPKoObIS5Y9clI9JzWLvj+uUKi6EopGgQeXYgY7nhor5HKcu/i3mMdu24GTsdZ0WWTw
UmomcB/0T5A0VUYkspB2mwUq1Z7A93WO9TbBhZszaOx5m6k26sRmIN4J1CnGGtHusYnZzaMqtILo
BGlwJU8emOfVqm0TCwlidqLBVvam6ETrCe7j9wpd3/BSJO/TnN9u9eugYWnzEPCc5NRimdtIBNXL
DAVUBatsOwGNNEdDycbIOxT+YEskLUPl2UMhJLHf9C1yjKME8WulgDyXzXq28rgxk7C9TbSWOUTM
DdyzEgBhFKWGpJcDtUDHJ7Feb8NEChZNwEgK8cFyzJcRlL3Fmt9UMWqX0N6Q2Pnz8OLpU448kUYI
oFZ2dQLHGrBQMjIB+g5rtwGJFKGA63jld3Xj1m9TgKO9keJMG+imvkKVQVtyWoJmV3o173kTM2J1
NUS/pPabtkD1OO78b/rH1HW9ifPLfGq2K/O3wJV0LOfwn2g61VHw/AvT4RPw89sNjxSdEf7m6M/g
QssZLx/HC0hSziTBFbCkKT42R9CbLPEuSW8bGZZ45VsuJRuybiK00lLcTz35KZl5u4LqGyUjiE/d
0kQ87EMxjXnmnjSYROdvJ4BfuwMBLWc2FO/JY8Kd5mY97t8iKfKH6feHjSBuELM8lfvdQMvQ0qcd
ZHipCoc9pPX2V+vpVzeXwGKdgbu8oSpN7mDjFWC14xLyAyYcSTnmIzMDuk2JsiufgDZN08JyisRx
t7xK+7EhInklL4PyYx+BCDZ6f0l5qevNfvfgPv4HrUBENeJsNNncS7VG1lQ05LgrY6qWQILdBfWG
2XyidhG1tkHRQSQG4d/UzhczcMZXLbIRU8kY/QwcmBddMEjn4xcEGW+VFDSjjNuHkM5HCy5m440h
reXNyXDU707l6e1mhtzfHkL2eGUXmLjc8r9bxvCeojjIf9qIrU4GAwp1sxpv/9TF/kf2mHCvN3Eq
LPCXQTn+nbWohqD59tJNK/i0J0V82cAnjHfWOlfI0oZTA+BIIV4pftxolWQ6oUeKzW8WtM+K/zk/
JazDcCUdJQwswNxhmiAM31mkaU6P1BmCf4+ALPvq8c4YfXV+gtqUV1bMX6aZlQvcwH+rCxKNiacy
EykmLl6JvI0vnLOaFxugirAJXBIqPlJoYK00vvOReoE8R7/YLkrSXriDcyf+LEhQOARuUbR8YHAD
6ETipjOGA9JdTjvr6OLoTA/zNW4Qu74atojd0xZJ+2yRDZu2CmaWtgSQxlHKqQHdbLsJXjnwPIAe
FhamOnOG5HD5J9Fsyg8XivQcfnJiJeZGrgcZmFaolqbMEBajPaOUTePzuXjETmCKzddkaEULPl8Q
+9NKNdlaQi9qBN3FZDDh9HT/q41fzQ6QyQ/dg9toVtPJPn0WiBTw6sSHsGDElqnksPxdd3fR+RnE
I1UbPueEmhzojt9zrSmxphwNeEESkzdwJiCSCE33Iv/JDQK8L3SWNPEDgctmL3zXVe7AilXuTtH5
ea9DMXeMzGB01OEqdMsp+Mgewhhu5gdgrXy2b7fqjpc8QhIgfsoKadeSeiJOTCo0yfsIFcj3vkKX
dTj/Jr5oYMmeknLwaCOYxQ3+HZnCUKLe1RAQqVMDUAgbWD1XtGgzLDkdL4riT1eZ1eJBurwDmBjJ
3ngn3ry2wYbtXXT9jMVwLxMZLoU7qx/ZanWZfkSirI5Bv/8JAiJWRmDwncXldwb6wSCgdL4mB4LZ
bCxyXMzhNr+xKfC4HlhXpLdlNxTihfGaibce8l2w/H6RXOOdMSF3TaAiikUBn/p5TT8JLFtw5dzA
Bn4nT20Ghes7WqYlSAEbExtfiwnDk5F6WgNAzVl43XjtaEf0OAyLb7mWuyVVF3XauFZXAoOun44D
aBD9p4ABBTdTNb+spoKVHjOt0e9R7zX+Zdb8F1xsu3tCP0dQ22EvF4v+g0dCag7iXQ9MmHjeo2jd
kwtQvK9uhTZFS7F2D9Qby/HczBwC9xg+OlQ55GYDGTbEgsGU9wKPSdxpCOarjNy1877gZJbR4w8o
hPtT1Qf+Ch/Rg8qeGKhpFbcuaHtERonF9PhhSQZd3AgS0VGm0JxrzaSSTmAOsM1WctUeofK8FagF
SlVa9HhYwzP6kCVcNJtyulu0t3lOb1QSsOOxJ5BicUXuo3tvuiWt1XbCptCqHt/vDUVYm1ajGzQU
8FZNyBvkauiHoe+EG4DjNZcNYzjvMq1E7mN9A4AXz2CgP+iXcyULZxisOQvbjNv3HV4ya/bYFfxi
/mJaL8zDA6td9ZVA2UcdwRCVZ3TLUrXIndkD8+LTmdMS6idnXmgk/Gkai+KoyiN0XQuWGicaJtsf
PVgkSYrwL14zhQYqv8yj6QRv2kk8tGqDNTOrgaYKoc/72weQ3X3Zt8QaQ69cVhdAuzJiDPKVD8jR
tHWeKGHvrM7kcjduP4e2adBEzxNbL9htZutTT2qsISgwo8OmnhRCyIRU7m1ZGu7T6CrCjTAcbCRp
nqYqApbQf2M8Ee5qf7S1xRDQ5D/29f7jIYltdk2QWIRCKr2o1YdBuGTab0I1mwjR1uj8OrOv03IC
BnUkK0WlAIeICZSHayfmQrhy8YRVzhOdA7w5uPpzSChvzvmiEwbhatBjUiazueRRpViJX7PcSShG
880denrBCvAgacdrZiEeE/uCAs0YzjUHXUPm3luB2ubqg0+XkLxsbspPw2uoqZhxjlY0LAhsBbvB
V3UFOFD9hITdskx4A8AjTx+Pgy9UNe6At/9ITGpCbkx0+AUzjDlH88hAa9G6927FwD7SkAPA0nCt
ZzEYNThZJ0of5NexPcNjvLMYiVxSo+jdMS7/2QXM+7VGQYU1uN79cTmq3u6FsjL7HXv2//lgncwN
Gigo9zZm7EG0CPRH/30rTUsYWztXEVP3gW/JhkGRDxnpF7Sd+LQVgzq932ukcKApwx0kailIGBxm
KjRkxm3BXM/11DXa5z/W8RRe7fp3yuoY02lFKvxRmziSvQcRyvcx+1WW5g0Qlf/epMjJSJ3jKicl
2lP3+Fw4YXYQN4CZrltjb/Hk88LXrFU/KnGjVmvaAmR8zoHr53GGgFbnF3lSUcd8mt17th1t2v2E
AfWEp1N5ct9E8Y5WJec5qGLEkGX14v//2LDqayEx+4iKfPrHcJvQXT2aci45Ox32zfdun7Pr1cHe
nszH8kRUO8e6tpgIkIDgLq7czpZYCAcxmaHao3u2oGiqjuqIqQqnI76jWbedfC9EApzcM6q1GR69
3ko7YIaLu5Jfhz6GQhQuHBddGHdrKB87kiyq2mVM3blpGE3IjhevcMNqENxHo5n2UrnjWQNKHF6w
ga/uij4OLRQT1UBSiMyiXWvinlWuT5a+JxTLeVodlyy8zZD4OCOT+84zfPUUa8rv2IUCmYMBDLIm
bdzRT/mUqT5Onfc1yENEB6U/71bR0Ca1HuEfdyf+ymIhK6D9F4euThDdQ5iFpJls09S3MFJnwqmI
K1t3ctkicw7gbVt8UMzP4x47Fw7ytCFOuQ7CV5c1W7MsNQa03MiBM5fPXWK3BVFS7IE647YIO6Ts
cNzsIPD0vFHzOmOGMDwqM+IW6ixMPSI832Tje/LtTMxzwOap5oXuA3b6z2aIo+Hk7x+if45rAGzj
d5xMSODx0n4BGdCAQOlB6nddUKo9tX9FMAQB15PFYHj2lUIjOyXjPko7CHHyAHPWjad2v7YZcD1U
jR/mOOKOHjXAHpWRscoMPUydI3NXtKXLIuJE67yfYY3M5OPtqjrSO+1Fq+WptTQqkQ8om20tuhMh
03uPL0Vc9jOXDI3TIWFkyaJuxvBmRpnv2r//yxyEpvwQtebKikDMIjcdX66LKeKYrN7TZHG/0EE1
P9K3IBLEcIjhPxnYw5rWW8/UgoIuz8fYAWVY0WA0+hF389ucQh+YyU7qk458PjRuChA094DELh+I
kCs2/loOsW3GwQH2u6C9ILAyuU1hhmP3edgXT+dxPmpkJ70BT71PFzQ52xMjQLLM7ODr9hWiCDdA
1a3FL37++4dxL7CHUZ5Gq5jKTUICz2mNieFXkEz85yaKqV8nUcTmIDGF4rDFpNmSfygF7kSmXv9V
+l5IQ7U/NbAIo9K2Nlsrl+IHOCkhPjzBqROdt6JSzVLDfOF/4N85YlYYh3Ybk75h10tXwUGxrvY4
JtD8aQGTAVvxrx2HnkXsYNp9H580e/qscHxnrD2s2rz4sxXOeN+IimISN86HDtjloP/IIsA+RKpR
2ER6+oBoeyqhvVcImi0u/f1RN5exlAVq8xuyzA9RkQbsKj5xjXXv2HFqSdQWhxGIi+5BvKdP8XrG
sKTi17y4WOFGTMTSa+xKCoz+wmvA4+RxvixM/6NMpeK8JDZ04ceD1ITHKBLhtgTnI4QRf81C3Hgr
fohRbm+wNuHrIzrRV43Zy0V7KfRwDdpW+nKIn1Er/2opCB1sUM0ziKsrNuZ6VUhsprQtzVmjy99f
R5OktGRtCyXHVlcFTzrMOydJ0JwC4CHzSG8Ph/mXr8UHYj9zGCkZddZszPc5EYRW8PavnkTvuHTp
7Vt8tIiUN67ELaH+PshRnGLAP2LGPSHCipyGL7PjmPAxDjs+jyliw/+0uZoYg029L4RSnqFMauws
0jlCkqOHXmcRIkbcXQt9WJCzVDCtsQZDAigxc9HAHSbTPC7AYLckD5EQwQV6ineC2AZ6cWCet/Nb
iqEAJfRvLkall9ZBP7MCcDZeV3Ov8Mv9E2NIfP0zKtNadQ/5FvcthDL6vAmi6UEXl2JP9Hb0QtAj
YJkphB+w0acyPV6sc+mkYFSYX4pL4OjQ3HMcTImUWUBe1DqBs7TRo7TWdQaYTErfaVuZ1L5YQ7ao
Dx5kKeHyj22njjXP+fLzaRcDh2lX5hPQvlflaQIHP7id8dPuN+kHsdOBLbxTL9deXpexotm7/YCw
oXilsL2Q7E4scm25s15KoIdVd1eQPdxfucnO3D1ww/5tXGmtarOTRm+/3FDWY/kPr0Rp5DZNUZdr
HtxK6/KSIAbgRppI7o+iIJ6RPa59lYEq7mzddzfMrgPs4RFM/VmdM67/i8wNRvAGiRBQGueZ9iZW
cgYoIfasdvzM6Jej0m9+gCA4ws09qMNKRLKc1OR5++t/PUnyRQTawrEvtRs8HqFPt5COSE4m0KFH
9hSPjUHHC84irL1aZEwTVlpGas5BRfoRqJVPmyB6BdSHm95gTRTj5gyZgfq20rHPnGAsgMq8OXqP
mTST6dY/L4JS6ej+5CTUxBE5kmaLfNbXQcZMYzlT6g+H3GwyLyDG8i73jdXwBks8lJo6geBAZUns
TzdRXChh0DbJHXbKV7UfI8xVuutoHeYceZKFKCG3ZZ6+A23mX/3i5c9gXjALPVhtBa0Cvc8nZozh
/nTBiHFtJ3XIleH2MK/aWpDzBR1l0tuz35s9ajCKCqxfEQ4TYIUBRaR4Lx08+Gg1iBS0+YnJA583
4GZh6QboMMAGwNDs3rPDJRY96ht4cpqrULH0woYx0Y1nY2JoLURRlmKfL+QV0WA+k1GqjTaxiVCh
UmTOPGabZSNtAhbfxk2OdH47XJLfdHHFJAndiA9kWgoNMNWyetuc5St0r/yaxG5khnAaRbGcO31i
rFU/nAeJgPyAEP+/0I03gHNarBV5ccLxjwGmHbLx4r9AExOmgASf2Dtq3DVW3zkNpftqn6S9wLpu
WIARiYoXx05BqSRv7KbGry/gohd2btMQ/zANt/aNX5DtcH5fvS6Hy3/kgS2DZbMoQ+gvyoj/mDYt
i63NR3DcQcwhnlGcqFnkWyVx65yQprsgH5+B8YOyWyUTgwL8MAejxHHsPL3iYnOLSTFJfwpVUxHF
Lpajl6Gq0Xig+/GVuuI0ABllN4lc24heqAGsxr1sBoG/mQMCQBBAeL7IabP5s5uFVC40z77c8wIR
R7FUhcYuMBcNs353tKc/OiSJk9bNA4mK1BIoRIYwZFVtfe8b3wRkkr80hJJzCS43vl8L6u3ynhbA
E8SI4g7BiB++1GcBFXXTCwKVCz/Xr5QkmNKyS7DSh/Kn7jg+1G8+BotFRihKFU3v9VM2AMhCsVMt
LYjQ00jiyOPK+IyDKAUufPjDISE1ykQKxC7a5hRByJEHpbf2Qdu8+Gydy5x2xOnnOduHocQiHBCA
yLeViEMoCGgYbRdiVzRNaqzOE+QbczrWzLP7dbo+7neqYztIuRg87FCQ4r/4OfQMDxGLB8wtR+SS
lnBgbdPt9S9Wj39CFuFSV7AxEWoE6FeiGGu9RE1YuhgPFPkGFIZbcRrWsrs6oQ9RusIah/FEsnxm
uc0hu9Wi1BgEqIFJSUUk1UtlmWW6fOuqcGJBkcZZbgf1CWZIdOioP8qXnWJtFRqnjSzA06pMdp0y
x+HkNTyRT+Xo+bnR1SNbQqYrHplaqKYnVmKBhFVhoLj4yCi4o0Lu4KxxREz+PQoctvHr/wfasV5O
IVFtvgRl4w+x9jvysIKimpP7ePMA5KlwlSw0fN5Ht6As8uQ9LUOcZztOoyoZVWPwsULkSy0h2jW8
BTFKu0lgMgNpQkpG+n6QrToyfhdyvYSM0hxQuw9VowfoULn7cR12qtIgD0F2qxdi9dG9eZ6RcItZ
pX3w+506W1/WJpixqam6LXckmaeKeEKhF1yMAFl73bnn9xKOhXhZhayBdfRqSLYNnk3lHdaHsj4N
r9ZLpo+F2viVBoyu6NaLuq/LDZ4m+5CA0ERp2ZmALqqs6a62PpQLfUkRHobSa8r7mkUgxyMoc0Gl
ne2jKG4o0diJDrQVNz4zVr6dbhK7tUZXMkBsCfLwsIVd7925Y9Thh22o88l2sbtEbc2MaPXT0jPq
RVfyzffNCxpe7fC6/psBWOzbVYWun03innFg9PiGvoUWtGdyrNQGFE/NPO22lhmH09l7e9LDTI0x
VjB4+4yJLlWAadlnGHq7zb/wKzseT78xhl4Vd2xxyLBpNqoVzy6ty62P7yqUJ0oGFeZXn+LQn7SX
tCjfke/aVzAGlKZvssUN+pVq6l2feEnuZH7+hqMdNqyYLcLi4x3zvsPXyUtB81v/UJ4P1R+w1Yv7
wA4tfEOQySWgcKn9oabGk8/wbbhrOQ1zWkiieEWcfvB6WeaIgyLcSfqINcrQMfZiFWkylQLu7Unb
i4dpUM2wQVjsyBxBQ3xppcXU7KtEeNWtKsOQTSBm9puTDfIZl0GK6xWquevBerb3vK/song+bF1q
weBt5lwpWKXuVayYTWrJAo2x6EalpLDZyJuWcQzvOKYtemmDqA0p3J6trUpBoQm4sppIrTFN0cS/
EBLl6VcufxM/isCBEqbbz8ww6ilFONsaQVytSdtYV7tpD/394pNPzGK8O848k4t8EX2zIMjOgkxJ
uR0mxnVlHXa4lm1Wqw9NEft/+OOaVOp3v7Mhu8k2c8rUvyYHExQc63/60Y1T0fL3+pS11MJoHTEn
yjahWtlG/O7p6hM7JMi88YNkXdPOejvuunlg8gH8MSUHZnMbfmCSHolRX5XGEjnw7MadsxDYt4sT
OI5NtUSgxZO5GcZogQfvehC81RbVIoZWAcut7WXzXaIOnM2TCcrmgx91VkmexLAy6K8AWez6Dt7F
b+jcfbAyO6VFe19tDiXwvnS+M+SH9BuaO2t9eh1/Ycj3CkxaosFdv7DFT1VfaCtDxZBWrb5T8C+h
ndh36caRF+eZMJADxE/8Lghbuadbptgzmkucnqoude8aks0fgwy6hnunQGP9hqMHajNxuALwPPGP
ADdzlCKrOL2eM+LPmB3/sAjcJCz5xgKtRjAoX1kGIFM1/RsnOUGFaoVkPcF/rJ4KbbhJ4pa883py
EviomWJacW7QgeIIvpC3yzyvD68cJEuC3DL77cR3o4VCrbBSG9S7AGVdI7slRt7U23kQNBY+7tI7
KNgFy9pqxGY+uPCCD/VoP/+ztMmbbAxfFispHz6iTOcQU1G8zxu1shTsKdEgmvMYuEnrLgBogJuy
cz/0EqhZYio6eUfB5rgBqhnDQFT/BpWvP5mA93b73FeG8af9umepe7ywAqqiLG/V8Yrcb5+s61de
mU200zsieC+Br9/CvI9SQS187Bc0nX14Z5o8OPopYFpj/WIOPWgCH3P5YPJmM9lqErwPzqb/SAj9
P/PS+jC/0BXICBcCRwHo6MLWfFhClbOr9obEmUpN4cvPDvTecb/ZdgF807PCcS9ER94oJiNrvIr3
ThvD9WxXhw3kCWhBL41kShAJh/iD8Ue+AKFC76gMdJiW3VMl6ZMhLWJ1SFTrVQdrQFoQjtg15k2A
tq0vACjC2DEi7PsnEgj3qjDMyECPcwrjDzP3Z0QbpEha8+H1vRuPPOUI0yFn+dRYCPtn0OzXimMH
xx1nPhl2ZUqDJU5NjtUIMe7vD+0vt9z0zsEC/MKG9VOdOFvvyiTqKgi8gVjB6dAYyxg+BH1FAHTF
HtNxR4/yze9i6ImGoziWSYYgRhepS+Q853WK+D5zHpit0P/VJkXXFHmXECl1KWf0mo3PyF7Al10G
KAQ8x0XQCbQhwwAmcSYNfdIA0gRyXA4gw8ACbaT1oWJHFAlbMuBC4HSWroFGENvvjJRIHRMrCBxJ
pDdnvG8WOP2sRkDG4dgwGbER1QMYFQ8m3rPaJsHDJpHI8qJ81EsZHqhpsdjRHli/ADUPwDHxV9S9
Km4Nrd0HMCowPeOu5hq7liy9N3hzgFukvBM00IYEPzLLnhTWrnV5lxbUdpIlJCNbTG+IpJ8DjxEB
4th0L1wnis6cXgH0Y0yXncZRlUUKebIBIsb0s8QsTic5oyz92JuhbzBCDV6PgdHIwerBfceHptBu
fy3dRv+sfrV7SStRbbAvfmSV105UwMTFTpfEvZb9hETg5LOGIJXkUGp30mTZH6BWlkANQovQ7VYM
VBDrZcSNNMxHjDb2xS/FQbtZNuSWFUq3SeZL/W/n575PKxOyW/H2hbJGnI5pB4yYSccUOwg8P2Aa
yhX1wHPJYMC1tQpTW+XDMtYsAl86Bp7CqGQri+He7sS373JNwFKfqPBpco1HdzcS2mhtL+AmWNgT
qOZxViWhiwFWw0r6KsbOsOoas4jtIzTV3EWJtSktWUn7MjcrZKspJ3H//XfL7tEobbJ9ECesF1s8
whWSBomwqtpGi+HZ/1LnnksXjFRLDi5OBowI2STn1Ob65SN1poObpEs+AFsRkKxUUxu6ypA2ktvn
Nad5qEdpE8X/KaA/7pK/fGGZJnfbdtCiMGjVrNekteGbfOQAOtwHgvGgezMu52fZcrqi5riqy0Ro
DgEHHlheww3dmF4gHxQQn19nlxs/WjI3TKqXkeqeo/PIA6FHq+vkCfSl6+T+IlNMWu9Ziiyf0wX0
h2Nv4yfHS4WZr26aKN4qL23S7JmC0knLY3B6QYaCwnyhKiKY2PYnEb5HSgmTLQNsCbr64+oWwRYx
+Y2RrmbJH1thv5/dfjmKAuYvPuXX/bJMiwP+v4KNCV3ExVTVXLVU+px1rhUnwcE/JBHDAkYbdfef
qIlDnMKA9Kdi6TdpePO+2bPvZGlAR4vY42pTSYqHFRxhzIjDUQOTwjq1uz5QxovwV4IMicgOb1El
bnsjuuRw2IkkE9FmkowrK7RAkt9/4vQZimuDs6GQZhc3Rl2e4JOXe+b1AJDVWqHL9m4GY76iVVFS
x0Jso7WE5r+M/qNa4/0lmUobAlXOfFN/QduEsjuK7Ze25+TqBzTXqYtHOeVY82Bdct56HbiisRzf
ml+QTszC/lTSw+QidMYAzA2WD1q5Yeli/TXb65gS6gSkNC/n8XcPeI78pWMk+FwhWX5RVNIvYgQ1
oj1Kp1VivEqa+AWcee59aNYmeC2iomjbgETU4OovolguUSbK+ozP7RZKiUnSRiaBbw38kiVl68cU
X3KJFgbABM/g4CCGIdHBK7M6ExG371ZspT8R3foRrj/N91HbOLY8G3iM2t8RbBdfMz+A4UPs5PQP
L+1BsezOzy03T4A+m0NIza+tkoXl4U/tE/Tb9dztLPk2gX+Xga+Dg4H5OL0FvrK+qGAnv1u2fSQS
lQeeycW300nrFOnuaV1CjRShXrxXoQwQp0dyTY+tH3DD3lA+UedCA0cuAXMYVW3AmHCFa9EMJoef
0LfQhW2+/l/bRKHtfMgxZlF4rZ2+F/K6XYS67XG54lYMO5lTvIMTMI717n7e8r4nErGQd0cDcAUz
DquZDDnsMkLPTPkO75cubNMYvyyL29wiqBmuINeskMzYGsydk0B9387mb8bn7od5U1xI2ePxcXMf
SG5ntbB7PEktcwrCVLQcCSPd4/nfD9W/wa6oqIy0/J0pTfflP1PHh2tY7WBuMBFIveKCbqcTUcaN
CeuoNThztx178UPXUjkhljzxTxZzWPMV+SpsW1UNyr3f8JjjubXcVHBjeWmzZu37cJHTuykPYT5f
9F4eYyMkmICMchlw96gZ/ObtaQ77Vn1YxT5mpE81T26U8z6XJr2fXBOsuyjx8Wqq7D1+lr799pYj
NjEnUVC5RouZ8WdWvsfp3wNf5yswl7gNINUhqzOzNP9UVecBrxqN0KUjLRvdfYre1XMyaWNGZIus
pYskLfc8fdFMJL9bK23S5q/k8b/Jc4vUNysBU8oNUOjhNhnm5qFOpCbYRKdfNWQ6Dn4q3xXVg8He
gRFTsf4kM+oHhUkBQE8UrdVjG5CcUcG7t1e8t4bfJqmAbSoJatvR7bYThKpyw4YaaR7QzmI1iik+
cjNCLB5zqH3DRiwMMAGyBxDaafMwYpOexPTqfigN/pLN9Et410/SS8RuR5+j+bWmYmwE2xZw/4SA
shml2cZDk7bI8IWb1806SFE2Fr8POb1morKZXIu6jTYWIdVf9DewpeMPcZpgFwRkacixA+kBvyoA
w/O7SafBDv22SUyazTjj6fuATFfQXLTq18jsPXApMaoI3tnTzFka3bLlS6kTVJ0hlJiU3XaPOJmX
V3zAIUjsl4U/R8WCaK6urBAg2eME2tlfHsBuV6XUg+j/XNJC2aNpN8MFga3IaBhVwNU2Z5P5MiVf
6Vupm7RDyBWo+BLmpmChh5CY4aIHsUEZfmf4B97S4M18kH6SbLaMb17Z4NOm7FkTZB3DZThP6YPZ
/WoDBjGtBY5mZgyoM7TtGAbYkCDmJMsYHGIZQtv0FZlmHkrl7H8zJBZ7Fk89jeW3ni20WPIwgtkp
lPsJyUxOjfPiu3DjEzEl5kMinevGSzqSYa539YXluLUjRVnmrubK2Ve3jjvdPJydbS1Lse2gyae1
2Bk28o7nsYcayaAaazGWB9rN113tnfn4kO/0U+D/xoYz/3P25Wz9zO3wX/lRpix1oWo0fDZbNhcP
4jyYTWrMBCw1/OWvCaYnp2NrFPwo6fUNppkytx1dFbG/QhOTbVzq7qKjbs0jt7hp+5m5s+k4v4VP
k0pVlMz2aR0eJZQKKg/0RKGKCq/Esp2XaDoJGPDl5jn3Y8hnzsE4/g5iPNCF4Bd/3QK4LZjzCZ8H
dWmqxdry8QJQSZGN2hJYWaatxvx3mwE4HZNFPRZKC4JXWKkK509S3z2xM4EJUtm1SWYTi1YMDPb1
Qnsnl4aJupbN1caNm7cW9MyeBPEVXeviP/ZGeHfVdfRVussjWxKpHK8ew9lyjbDi2eOpr2/CtTQw
fGu7YxB9ripR+LlClCZ0VnxsHOj0QpdD6zl7UDNLjgtypgIKLv/xHF0vx3kEzywF9jJN/gGDrVc/
YRjEwMEAs4IbKHwB2RI51/lMbtXDM84llsRhbQv52tRMoOK9d2a+J4/dkQMql/gaf6QePc7cFon9
AK8EIutuSJPj7otWrOgg+IFLMPW/u1wdRkIG9U4yXc5Zd7Do7sZgmodWC/1iK49P9m33Jh7NA04H
Blplhg7SA3KAJD++x8zFOWC1wBR8xLbpLoNUY+LcK16mi2Qfz3Qt2vegQobuYO3tcAsvDXpFmgQB
m75Us9N1Zw9JzCCqTUXzmn4tuLVQgDVABbfDgjQ/q2NDaIrNmr/SLjo8QK+qpiUwUnZ82v1Adj8H
Pd+JQMQBmpiMi4JXYlyD0/TvRlbUuQaprjUkvozn7EOgZw+u1VwjhSQZwZCHnqvEMz+MRGdgN/2U
xYLnpTJIy/QLJgdGygvyVhIlVhHQCItara04vSq1qwQvjOW251Q14yDzymn+adPun38Xu8fMvGmw
OolytMiYxPwksfwux/IraYU3CvPMera9GJmv9nKFUMgBh3kbm79vCzgyP8Jr5cXcYxBp0DH0aYnE
5liexw+iVnmcbtv/gtvPFLe7518SED9BE6xN6wntfh+ZGzBm8jz8UA10yFPbRECVnaxe23Duf4zs
MwyCi7GmePLwSoNj+SzqoIsBupvWNvex1iGtol9khTKF2MyNzsEsr3GhgLXJWLj7rEpdzzBMW0V7
vFytlX6Hk9TkVfKKCii6jT4/cfKOtYvznPyKtxP7jkxny44shgQ+3tOeg04PGc0RUCxV85ud5n2s
v3VhUZiO3qW6RvRZzx8yPoLVKBNkDwsrxF79wVKj8P6kAuWCE11/2CM6NwrEV87eLHXmBK4JKWok
kjSblpJIdh7pO67liz2mumdZ0LLrNJAa+ezitfCrDzwKrO/l3O/Q+oXyAB2awu9WaduvT/T2aLAu
I855UHit+24xdHk4iFRSfBUvYFvnWnC40dqiOfDr/yrw/WyergfQKYv3lwWvvt8fC4KykGV0cXz7
mP9ZmlYoKHKFXE2EYnl6MWxfD4z6ZYMSaO2c9QvbpoNh+2z12sjSibXLXcsKYDqbMmRy3U5ONFv8
3PrJGbNij+H1lRfaYB11YJtMz6W6NoV/swcw88htQ98lbW750eUBpjZYByZKr8ly8k/Ztzg0TIU9
o4V4dVKS9a0FxpUADZymoQLxz4ofA8X/SFXJxiWP6a5eQIwuA+lprjWOrOicoQe2Y7/4oe4Ys/hO
S3FP3uehRK3Fx4UMtzIJz5cB/5Z3RYmX/lK8oYS4UmUs6rNw/vV14RZoYG4Dtmxn6by6xBF+E9Q7
CwUMaBTfQHfm71dfW7kj7Qb9K3A+LLjFR2hnj5plgX0ZODT3oO1ur5SGoFwZ8yOxvEjuUJmXSw/H
pETf/4YjBBrJpyKdQdf4T75Sz7wCn+q31pw+BLwOdEj4jX+LkdZLv1jhsze+T6LhxBgHzIhx9zGa
8MJWoIIcMeJx/VUogAeMW0XxBSuqEt3nzpkVSNHWdyBGkeijLPx0LOyfaHZyv+M8fTgoEWPEa7Ex
QoQ+YzKUXdsrGch4ecodeyopIrGGa3HNRpHemE5ArXmzHEc/79rL13EOH4d4C107M6Uf6yyPb9zI
o66qCTDCBnJllqZ6jDS65x7yV1J+ND4npDwBMCUF+uukCXfsWpeZ0nd/AK+xS9AHHKoww3HqIIXL
3HUynXL8YT+tZ4aj/3DAkuszFIsQVrjg4HKkTQ8OtdXB74V4ppsWV2VbXURbQFy7ZHcC5gvRu2Gh
tiOP6sp7yYBzQYYibkwGqn928AobqsxO6sQr2igWXhSTmuCcPdzejONDHEdKq6qh+E60fb3desJn
ywc7Y/gnw5TVHGu6muUiHIPny9mxj6QKT1O4wuQO1mEmYkCfXCStqYBpBuBJUIFDxE95E5IGTEIu
vR1GHh1QlInCXUNEZq6D+2comEkP7nCAH8vszSxSuzfnuvTbGwnbPYCIGM4LQL3rDOOUCDHEV/tE
uK7d8zHTHXzyXkFsjhMNru66rnov4PsKcYNF0S4bkylw34gaMOu0i5+/eyarzc2gFv/5xrse/EqS
ipdS9CN43VjT/v/q3DCRFo85jVeiFm4rcDC/kfL9dlNkwUGjo2szhkMOU5qzuU7SCA/725/2kMzP
+8x1DNTa3WlzQhT9Nx7JTnxv7nnkgCT3xeQRkX9JpeIkggoQgDBTxXzfBqdekv5t9eeAD/f9ia8W
dKsPAvAzVbl7Gq21sK9qxLQ/cabmXoDUie9g5h7ua2+L5S1FU/E3xFFzHh2wPybGkKBWwYmi6XQe
go7DnpjNY3cHAfOgK5HEx9OlbvTxnpOwEhi+Np278IEtQ4EYq6Ir5AhUhtv6edEYvNHzSwJBjjd/
KPDpFn09Ko9o+g+/LVOo3gECiLy4YeyEup2AudXD8AyKY6Hr4Cg/qbjnRrCwSawKezjUa8N7P4cH
UdPPg2Eq0bo9Wr08zX40bA3UAGflo5OMt+MOZQjLQwv0HUmQpzYcVCzQmRirOtRWo9RwAdE5Ts03
EjnznMweCkORCmOZDIaU8nWAx4Zf/9JEcsbegGzG5cseQ4hgAUmUy/QOB7aU9bwvY+vJa44PWdCO
Sb/DgOwEt6QlMUsSH6RLS0cjIFYvFFC44Mqgkho4iZyRNFCUOiv9v44KPhBK6o8iHFBBBzhFARLO
otwPljmlcYoIeLkrp/aKlX1e9DLcTS3UhM3U3SNPjUBhufCKVA5g9rkuPnwwPG1pHEmCOXTi1Gg3
xaENxrE6hFs88Ds8m4LHKxmdFqoAgxdvOtIxKbBhNdUMUFpcsixo6KFAXcmiG9Ozl0tOfnkHYtq7
weE07Yvxsl2wC5cwIPHFZXGv6Qe4ftJnRn/9nKoiSKpXNYcdQRfbzBEXfks5ooGMApx6tEA/nUJd
uRMwKlydUfccLEsBrRbGe7gnm8DSiZuSUG022meGU/Qch8LbaXEN9ynQqGxW2SOgQpGzKYttuBzM
S0T5JjWjbtNK8GNbAr8F64+7r+Kyq2uOp2JT7SdTGzsoL8JjgDzdQKjdpZp4qik2sLqzkDBMMoN4
Lydn6iRTJjMVBl9iA5Pf7gQ2uUFAj9n+Ao/01Dn2bA+volClhjawnp880ZR2t2Dq3oAjRWG2l1um
0ULti2cc5sBkXhuBwZE2u/Pl45Fk3TBTo0DduiENbxpOtVYotATRAclRW52fDRDsto/5qZ48Wn8+
ZqY9zFGbR16pQO4hlXb9/xXenR8PLii1wLO4zQ4jXB1V/5+wblR+KwLPOFiKvIMOycZzB6SUFiFW
akt1D9xXa0cda/ZhTncC0kTAcoVtHssqa/w1X3/H3ZAjvu6qGNQTkZqpYnbNcs5eIVXpfLGpQNI3
G2XSH7YwY79I3NWwRow9XmxcUi4pbfMrxcgmxCBYwSL1ZF2A1FVEl0v501Z5jylSSv+xfTyjdjdi
6C72vM0j0FQxiQrsYcVrGoKWCyKbbWS+493mocAGaWtsCLErzFyd3l3sNzVcrdy7jG0Tnc2sag1w
5At/Zd2AcKImMqD44poF0qIcpBQlcNTJ8LW2aNzViC9zjpZri4hG1IVHHhSgigmZGB7yBXiGOnwl
x62pcT4YAYUrIVC0ej1geaLjaDUrJIdMwWeudvljceawWBKz1hjO38F9sQJNSZLJT3gzmIJvpnOW
JrDTnNHSdnyw2496TS9XXJQScG/mktRwS6fJ3iWqkrW7xrqMet9+NLi4eWkm7VK5m4oX51vQCAI5
B4Y79hj/tCE5Ku71U34gwJRn8i9KViKoZ+3xsnEC0eSv+QYBGUdNrBbo4n0gpWADcSydxcv0YNAp
r307g2frk9L+5aT/SlD+uvYxTJvPZKjaJhR8ZMe8XEgePvjIQ67/iZscvtXf/LLwO70/rTb+VrQo
F/Mzu3Rf4A8AsCo0wGxrcVZgIxwW9/qllKBRy1Q/n29mUnn3cxkFj03nT5CzF+U87krq2wyXmpTY
eQZUAnvs675fdqhGVvx8xVhMPUNXuTd9UXFiw66x+XjtQIXQBySTt8WInM3d8svWywmm9/5IMn1f
g5GnGUD7qPYTK+OEszwVv1esf1KvtZghj79TXpgvsm9Sls5UpOjb7IxbZ0sic7c4vHyODUcmWMbI
uab/xpcxLheF7qZZE1ATwL0ioiyxNtY1BO9bOwuZz6fQAg4I4OuASnTKjjDQwo8w9mffQgEQz1U+
2NutfHmY6l8WEKumwQ+7xPuRlI5ncVd2gdXdwYOjE+hcxwc1yFgINHnk+44KnBGE72c6XCPxNZTy
B+Iv0c9/9Bsg56TjbeoeKjD0nQu4PQw1Gp5fNF5OiSAhMSCDsSkA/UHvGL3pTDc7eisSfpm9jx/R
qc4jRddLfkw1C4Pss6bYTObEYtk9Hdy87nwzuMeEHvDGmPfmuZqyN6LZ3srkaOrVg2whdigJ35P+
zrWK84PN9nMAGTvupF8dA9PXbpKpsS/Ywou37gpwKJYipbxImduXah6zFO3i+UZP4mpmekTY3ufC
1AqkPhcq/XyAY1lkq3JaRB9EUZ5XF6d65/OMtBpq/F9EHpOqQFFYjtqJR8Y4AGwcX+XwCCGOBH/J
7wjZxcyzdbk4AWSSKCL/L8Nm1iloRfkVvxgpFe1UR3aLEGXdO8W5IXGk5BHWqJLHnj0mTckBwuw6
sXbt7NFAbnAn7l7nBpjZBw9s0kcPtXHmkFU5HyHMfJtzGfw/jNF2LwU0DOiuJVDSmL5Ayou3O6g8
sd8gzUBp1MAUGV6+GUq+ohG33yZGN3zdAt2XyXEUxYV53o1f2Ty7/MO7F1HzUDU07sp2Jfo3Qya0
AU+95JN5gt/EbGDkOmCHIoruapEK3AveGVOG94fsWv2QdDexipk/lHsgGVpRWrL+E4AT95sx1ia0
c/kb5CKaPHADwsdm3xEbnhcnp7nwo7lM3DYyXtFBI3zwP/f1z2LtYZ1gYtDa5NXGNiE9NuCvJk2M
2o4yC4D1j/wFQmQC/7LzZVimpbHtz7+tUCQb3sZ/pz0HabqAgeWB2Mh3jiKTjpqHUJvxAUloa4lv
J5Hqo62vkZ4ijqexADh9XdouDfE287AhHweajAjm1HxSX+ebe0PPOT5uFlmRli5IxWxBiRtdBH9E
cTAm9Db8NewfKrEnLYWZXYzlrg3cPfBxSShph9CWtHnU2AFiSwDDnzFAIYC6EDWQMkVAgLhOnL2z
XRUvZOq1LdmwIvUvpI2DG/B6HfYAmWenOB+ALYxLZbbOeWkuRXCfgsbfTkXapOWankAx4LnbGXv6
WF5juYSi6BqXcwqRR+B8y/r78zOy8V8Ms2f3/BcW/6cXZ+m7ReEhyIO31blt6r+zVnxQHPlOktNA
l28DwE4n3KyY6ga1xe8FNTFkv3mBqoO8bvFzGZc93TrKRHXISqIj8Qw7z0rShwAIfEB6xe8kEAdF
S8VutHj45i5idbQIWAUdaAVMxVktd4ho2qZPW5tHy8hEpzkoc87UkId+JnbPzpx4sVbvDfO9487W
kxEpOdON/lNQRVHUaj+hIX1SQ0wGuRDFVNAkqKQmlfIu7Wg0EF53wWj+RyavVVjIs35rFJJaFUlE
JTM1egWb65aZfj0dw0z4Zeswcmk2WtJg1izIbmiwJ8TVXxHSUYoXWvK2KcRoEH9aJZ5HG5/MGT6B
/lzSw9Lb52mjYItZQa5EGX+nbHpPcGG5rPR/WVoKQqTMj1fyYA5AtH0Upaed69WRPAtieOzwWSCg
uPQAD/a9TygLl1ZZOlqy7TCDiAbtLDfZDzaukymewlvptR/W/wXL8utS179fRdFyXO/1VrSx4/7o
9ybzjpYTOG+5YvNyL2Lv02D0mA8AqmFR2Z9Yxct75Un+M05az4c9l20YYvWtimYOfACMKTap95WF
0sUh9V2BS8HnDRXQAJMoD5vGAECd2twpsrSnnoFDUrB8SEhK0EQ3hsupUt0LWnefRcYhGz+fzZcI
K8+srlTQqI+pgYHfobTs6rhpinnCThDiDEIBr+lkKrfsyGhCjAwXAoGMDqsnrDP7vGNGwe+ozDVP
aueEhVszKKYW1i98PS78zMiPcQZxYuYBsaUs41W6dH8IoX6fMtm4CKn8a/pIrYyFExkCxG5xRVVJ
+6gOxZ3hyp1lKJmuQcL15cvFzVEWDLOzhGGPYayGzEFLR+gHXLPNM5CVwFleU+dWZaiXlf96Bd/G
bAe7mYuRHeSxwQv1xYsOgI+OBs/p3PHJkSzwYIRQmYy076kh4l0kCdSFD9xJx5k1mnQdHXarqRpu
hoOb3GdonPkbnY/STOS7GEdStI4g54AbNajFvw9hr3ZZBtJn549balPob12Nz3HbF4cgtt2JwKjG
/QiAxsZBQrUE+NTGyo6P7kKQOY4+TMqps9vAGpS3G1QDf1mCTj0lOsdz7FkvlE9vfuK48T6uM1Q0
HQAgCZmrA4dYr0D8NPopALqUcDV3OmSKDY/vUZ52aBH+bnzGbVk9IQsVV0w9G9+DkCiEXnXbw7cc
X2YTIYcL4B2yGAVSnzjsk/i8JK7PcX2IPaE+YuCoG6JEc8WwZQjodEvkMo0OrJVC043QEKu2E9gz
kSkpLZZQohQniKxcVgr9/NfGcYMeDlzkyXgmHv5oBc6j6g576GE/Y5K+cln6SipO3aHY2/Z3eMKY
nAvLmSYqGUQoickNeDV0dpLzeOfC3hCAdTQTTHTdAYqLpVDGSd7mqrp6URPiBoWeILXNE/HV3B3E
YiEv3InQS7IgqxGmToIjIW5Y8HNbVh3o0UjlsR7QKAb6UowHX34GPTg4dMC6QPtgXO8NKTgsYpig
igAo1QmtBhSS8tcZJIUeJ/NXL2H8CFNTdTkp1rbZFl1fUp5TDnwP4yecGDgmj1l3mMyOAbNbuM3B
DprPug/4HtmWEOLqrlS59B9zoyPCCynDOwR3J9aPZcAIiqt54+cLr5PfurK1XgtohpUFoEUfZ1Wu
9MfW0swsYIaFvgcNY9hwI50f71hUIrsSWoPD3PiB5WaIjqf9qoSi93ZEG5K4J+lMyPOWWDipgjSi
/lGLCeW7jsLYyYocP9N0n7dU+SiRxdz1yYyFqgl2yVZFjj4nxhaSFKs1pbnps21v2M0oYJx4IzpP
yXTkW047h8vpz1Zk60HcP2CjTbHQj6SjnxLxTkP3prIk4Pl5W//rSqjw939g08FCd30HgsWD9qvT
n2fge7QSN6WI1LmAHm7GnU/ss3sMKdzzxI5qZOYv1rCBPlbKJHzVWSN7gtaEqvz5Uf7+IPNtjAQ+
6zIrukLjS7UyBm/6AZmaf50jbtDOiSiKP724BpsdaNPYRkpZixWc7g7EFCZupOFRKCjH9pNvTxOA
++rf1nNK88WEnMlzQfTLH7MFUoPxf7fVL6oqrrJcASlUFFKxjo9iVGFMkfjg1tdbEVQ/m280M0nV
Vfd8cV3kX0/byBBPdmqIYKJH5rwQebVik2j2pny2nX2Kg5dCw9uoaYz6NhfNlm8VM2DZZAIn4TwB
jtkCcVarjehkbnHRN5v+WeZG5JdQnsohnxOpl5O5JEH6L7mHotRAw+w9IIEVSTj4xbsgczxLCqLA
0XJcXssh5X01d3edi+tdDZ5bb4OEDmVwaOPvSRQkL+hUoi0ccPP6y/auiOWHsFvV/IMg6U29MQqG
UQ1jnmrI+ZJRCJ0mlRAluDQQqHpoVkdmIYqkJXdnSayDgTnQ6rS3Xk40FJqZZtqptN/4GfdaOK19
O+KgCanf0dthmQWuU432CDLeLowdm7YCK9waxXkRc7yHfT3+64O3gbkMIWXXoPqrll8IO1MGwNRA
Z0iMHT1cepNb73EKj1U7KkmqMf4vEOyG/jnjg6AgWG361HsJ+E+cn0J8ZP8G/+00kNN9YyA7deAR
6H2KKcBKr0Gjt0VfXt2MUQck6aXBH56KPYcNZQUVLmGR2yK97w9SHN2lR7BSvafQXFTETIoNINN/
uTncB1VRSwvyyl6gBtPPS/h/6fo/rk6xhBXUw+/EgNq/3WN9cf7N5l7M9QsD5y9iTtEgEit5TeIs
t4S1YnilT+TE+wEtVxfmQ/2zd/tVnguirXGpAyA3KUHz4Sbnd6dZncpPTk9NKc2kYtarwAONBHRu
A2NrpZvGn3MG4ZH6wVW5PoXM3lTZp8aftUODhG7yv8io/N3G8cTj6wrk0y5tABRXEVkr6ug3vdj4
I81cqlVx/z3OBowrUf5lWh/v4ww0g1r6+2+Wq6+g6YTMeZG2mhsvTlWZGz5zo3AjnyLZcOjriVh8
Gxhy69/pfhjmNd5IVYXXwOPWhlFa8xdzo3OeK2KcGyui5SCurkNcWwnuC8z2Ns+89GDXS3HLW9yE
Ai1RKPkeoDVbvxKnwewPgX6aHeM+fIgVX5gSPHc8SJWIhtai+Ot6TPC6BO82f/HcLaw5vBksunA9
3IDzOsfOpKLQGgX8SjjNl7JOJC+3eT1+fUFM9cCqiLjCWyaS7TzidKqsjQ0hd/3LTcpuvTEt8st0
5VDapJNN23BvCgWlR1OxjTv0DKCZA/UrsGn/zyb2EZe79IHMEN7SgbrzL2dfevLhkSm0jeJmmUQN
UFfK9+fmGDut+e+yAIEb894bQRhHughvCr/ZjcjUe27I9UDqcY/2xnb2uCSbJCar9ey0UWH5zC42
vJG1+EeGIsL4g/HQVUtBkHgNN0yMrDLV91Xacdp8oiMMEakxhKAgWL5po0dDm9U1mRDwkR1yMVL+
jkQBz8bEhohx+Qf5myqM8XqP/ez5RoO5tEBvNPtlo+uRxVz43dILSPhfWRH1dXSkYBWMaiHdY0Nq
2yqHGXbWqYKqTAmiG9X1fZCrleWRNtfUIlEU7Uhft4VD9VqVjl2i+0FBDa0XRCa4jdGm62fiAfWc
+sN4vhg95VnCWofQydrA69Z41NgQWkHGYhmYKOkPtSSvNAbNc2nljqTuDz0wVUWpkcmIhjIVosoz
9kGwzWQ21m61dc73J5WGL0wfm7Zs11FB/hstzG7kERCm5PnmvJvbY+YiAL3QgaOvn2JkJtwv6akD
q40BPMrleCtXqtYp9EkQeUU//w+P1psJZTHLjLN16iQqEpdwsryE3WE7R4O1n105ovjQgpqFVabF
Et7jIChEYijwC9DGAlhBqij6d+BwiRChALe7xNUx+gzZnz8p9HoJLXUjFIbLyMfwo/Mul2z9dATn
TOVvHdNkEWMhNGahWkAeuJ6y5ViR7aryXzrxmkBVfqDbchUtCSV0oymIr/dVOYV0V9qNjnoPUQie
KDrZ+CKApfehSwEjdQsTW+MYanfYKdqEg2Jud1qI6uF7G3lgFnH25anxHJ3e3I5AdAQRD61vRNZQ
TPQNCBXKUCEnPIkdzOwAm0p/4GL+nXJZEZgDtyTvdNhmoRk3/v62mLaa4IftakBffZfDuOSXZcVl
3qrTaC4Gd7vHOJWYuVhYTrKJN1lSVdP815eGRaeujBytz1HryOZkhDFRirbgak6LQ9HTxezdw5oO
Ju/uxRTpZPpK4o7R6m2b9ytjTHQNiQNsqxubOkiZutTvgqEGtzGLc12qp28DuE+8fPFSsfDW4t9W
h7wj9s33N1kWSHhbW4ngjDLwvcKYcZf5jSJ+kBrOGvQVMnQnSs47WgX57h8mbCX6FEZsbMKu6nD1
BhdpOEVxnvGLthgnTaEgu+Ey3B42aWJP4I0wlvYivz/nuMw27Q3iCz90zKY4fBBDghs+Eyy3ffYr
RkWEU71pKJA8FqypaZlJjAaaBwwF6x450kWSUeqVPmOAJyC15YT/i1zPSaJJvV3Bt89wiF6DA5nL
z7d7zOAZIoXQ4kCI2OBpWgQnPQAPdHTDvUwBAUlbJMVeQw0Oco+Pb9snoi41Tk98E7FfEfJQNCcX
s3tPxYQKPY3vc95XtgCt8tKjjT+rmfOpZx1LEYsBK6Vsm1qQwPiV6J/amn27I9tdK/91sufy+/Lh
72vv2XFCSjyse+K+ct+Z1BV21aCDAuLNQixEdUSUJ9NzDirZeP8btj/Pw1vnfHQd9LCOKJc4v7EB
j+YF6tIbfrPfH2Pb9aKKz6yzxzyJm0yQ7EdxhLf51uaj7zXIUFqAJJp1wstK/SkWEIt6tYFN8r8j
ibM22cxonmOKWMPlqbwQ2UerFgKRW+GtTTwHmMmB1/DwvuhIxoawcf3xJ8DPqdlhstwmqHaK88VP
bLmNFqKImjOcAxunbJhRVMKbRL5sjgoY0jpsxLBW+GVKaSrfDcVrzigPM+1SYVNEplSh4q/II1hm
f/6zg810NlXL9cB/5vgsp81H5sbq/XX6e7z9ZtOqDBBOv3gbOawUSm0VVlnNxuQoVlOwvFJRD9SB
gXXyVJNvrgXfG9cs75knyBAh/RZFnAqErjWWNcu87VWkja5NEHBiizt0bKs5taFFwpKuXWl8k7Pl
1YomVeujtrSMoCGjjZ9qc0qB/lCbBVbukTYS1bFIF/56uIOhhXERkWmlVgnxvCkZADlMtVtNlv9p
fJx9nS2aTZKolykd19uIs/I65HpDvv0D7X33bHueiXWRHXBcVz4JXtxOgRqCSNg2DOXTQTw1Xibr
WsHx0JgcxbpKwunxXC0FTtwtnKWbwKlXS4KvHRyrjZ3UKU/XiRnxH6YhSD8ysq3PnmgaN6idrd2h
BC0IUVhaRaryQYbDCww6Ls55CnPL6DtJg8pAmqDw//525c862N7mmVj9Kmir0Qbzh+Ep/lGJ5Vda
2N9Q6WGYK/LBUbbUJh3opaecDn8UkPnbAaTVuFSMEgxmCW7T0GiWUKmXHidWkiBO95uhuQ+R1TSV
9cvSEptgLb6fRjMz05bqs+oXBTUaD0m2gsByvElrR048fH0Xc6rX7BpO4maYKiHQMU1Z7nff2r2G
oY306Txxq4FnvJQX+6X4YvI+4eswjyxNMcHQNWfNr8ic/t4pF2zEwv7Yi9VXGq1qu5e43FWEdJUy
isy3lsdpFdPYLJ024lUPJ8o+k0pCUh+Ipr+O6N/Qkv+UcUE5laD59lM82ub3I2siG1WUYXCUQAUF
05NhUsDaxbHSOIO8E9ETxwKm14kw34efjCkM9xqY8BG+xX0IcYVo5R3lDDM0PrGejfCCNXKqVXfI
hvd7UFZcw7uSV8YNWgcCYwS1VJ7EhLQ5mKbcfhQfm5svRVXEJHkG8sFIMvBBI4ZBczpEieKMTJ/Y
yv65DBK3YcHeyLSiNVN/gOKL0r5TB80+293YHOZNaXxNJJGOjqwxmVtHDhefsttLjkuuFfrtK26M
juM841z03/tJ/98rp1GScjSApKcB2RG+qTujGn32CfBBbM/qPhwK67zi59OIwfsK++d2qpcL0DGK
qquQChFMMgNo6TVs9od2GLc1c/h5kzUbIdprK+M7mnozTR6Yj7LCV+pYAbHMLsZgRG1NEhqDUKxC
Ea6iUBXcdcIG7VGoAvOZC5TjDeOgrWJh1hxweMF+vuIyEs94MyDAl+aEIvdgoYJjmNFge5W+76t0
UBQ6b4IWWVGhfNo4TAsyi9yJoIuDXvgWDpJ27WK18xJXpCgGAXMaIfVkCcThXhNXcprJXgcYioZ3
TJUGsvDL7LZ+xjV5rLVm/bFzJ/ge3kIm7YBA9p+gK6zSznNZy7VD55Y3HRDGnpaQTAW4IPX79ZT5
uOZAD3g7uOqWqVVLDXjUzGPooCMBokAyP49S90EAWr46oahjcx+QiDtEdNd5561DFsoARnKGWA65
sMZ8guGiIqtiuCLhOxE16nfGf3s88I0FCHATOhIcRhFoPgNrwPBW7P01GRlPh1bA0cQCL7rZ/ZKa
1mbQlXpIz65S+hCefm33WmInANEyRGpHpH0Vk4WRCFqNWFWGzEt0xdXoyhR5zV1dLHgq8wA00HQ3
Wob/DEtLijKyzEj6cZUR3ZTjx1Gr5b+r/8w2varmE3Y9XwCEUqj6JaQ67YyOcp7RLYey0AJx0hNI
pUr2Vy4cSL5/sBQCyVWjpHb1JmtfH6JkPxsBJVr8yfaznbTzqwEmwsgcXADh3uGfZThdEwrndZDw
i4Q29Sl3y+myLNrz+bNMe3WF0aPSLHAlv5FY6uUHzgQbjvI6oDloQ/Rzlp/8jicd6GpBys72eo+b
VSXWDbJ40lAl9oOdiEI5R6g8NO34Nrf4f687r4zGequ4SJEA2BZbP1dhVSN2dkib+4uH4oNVgWLb
0+joMCnvnVuctdJ2C8wVJVd0lhkuaYLJI6MtZQiS6UDMj31QxoE7gyWA0VFkr3C0/TcffpSGA3JF
gqyQKK3hwd5dd1L7SfqcVGt4Cd8IzujvwAbXw4j/e2LJiK/i6R+Fq50R4lRI7NU+sAQBncUJ5A6O
OlSgboW6cbDwVTa/54VkCLlO99vYCsJpL0TDTteuEAv0R5/wtaNAiRXUaFLyqPVr47QfvVyqBMp+
r60H9B7LztoLdxOEfViGof+Sl6T+tpwry4X01Mi1dJmreL0pZ1kA+p+kgUx/2PJApeU6HixVJhNB
tV2/GhnIuX7PF71q2BMJ1y3G5eKMrLRcvV1CLCRYPr5rViovavstXtlx4RuCgy/yup/VfyESVpDQ
PhoAwB9mzKeG0BUssDNBIkw5kEFINwhoMwCffjVQIJjD3CrYIWZu9pJ+zv7PsJQ7c0fUodjo1As2
dHRO7awqooawJ05SVKOWalACgEBQteg54VK6nQL9aj60UgY8Ipd6/O0cjX7ERh7dswKZ2tXCLuka
KMXL/MyUyhPzsRgKE7lsNZ1MCuuuL9Y+ejiLt7UWc0EKRdffNEBEVcx2E6cSinFb5ogy42/rdR94
wIQE1cfF+VSofy2hFvbHT+ZcHTAr3hk+blBwEL1mdyu7yHVuscw8UUaucGV/T8Wwqw1FRSZrmY6/
R+s1158DhcvgR+KxKlsY4Q8iVa0qPEd8dLW7H/p0XAAcSJoqM/gFXxVwyPZrvbUHBTSLlFFWt0lp
ijCbuhGi7bW+T76Q8A4XRZR/oTcgesCLi8nF+eOYQTUTuoguQUsxzeH3//XXJeqr7l5s4n1WPPxi
rpj9SNYCunGAleD7hTQRzk/QW/TuVAM2tvMOaA2WEGREM4fLLLjanDx38J8Xd9DMFDJHlN54TFxT
/S+wLVTgQEaebU7tO4aa0VX/vDyXq1VeR5sKqiSrgCuljMCXZ5cIN8u7jUMC4jyNDaMTRqrc0ufe
N7xdGRezofZUBDwlx9TceloeFoWfT2Fm0+r2undvHHRdr3F4AeCytO8KGtvWv80nThRY58DzSKt4
w/G3yVFFP1i8Gt/ijDZesewuOjUKwBFu4S4z4rxdUOQVigV6qMk2oHxjd8+nmzS5btgVy4Etq6Tl
0Yt/hL/BorU3ugYCUI4C80mrlEYL1BLZFJKEb+VZyLjZu0fMgA/zfJ5hKe3t0BNxvUTzsPFDxJqL
Ssnmc67awP9Q2Y7hStnf90Mm2Jn9L5oZHJc+IbEffNPv3rVHXSWzDaMgvCDTO3IWCgVRiJ48rLU+
UNNoMiMa93xkVIwhaaoeNIX54LLJqxPz/5fYVS6EV6qLhAB+3CXSFydh45V+HXP6xmmmZ3o2fJ+7
4N7Sz5Wf+v7a/gad8pnTnuAKuJgqGxfY7fyNexHricvRM9Bwfl8ifJczc/KN1ixqnAKFr/5F3+dl
8jyEEG7GQdukdtZRx1QwNME84Wd9mIA8vofDdmdHwF9Y0xNVmb55Rdz6o+H7fFvfz7Dzu/0BFx1I
dynR9qSBrAs6V7TF2FAAh5SveSVSaftx8v4dbDirWZ4Cbhaqm90ZAmbA0pbSSwgIWH1zTW1mNmKi
mS2MqDrt9SxMgoM7jjjf/T5zA9q6KeSliY8ov/QPDwKHupn3bvRQqu9T1W0x1Y7L710EiVFRu2Xo
RfKlkbZZ2KPZRaUuHzFamJN3T3XGlpFaNq2t1hV6jbwsEVG5RmNZr+h9URNnV9Uf2ZgGZ9/HFG6K
sVCmWv3qfn26O6KcheVPi15NFNMD6vjYoa+GpZ6XkhqTKSh0XG6lrEgOoQ6qKcdizYaGW7PzXlIB
HBDyGcYcTtHG4WVIB9FpImAHhA6fs/dYtoRj3HbKEYz4R0vPEMZSv8hPjWzIvHox6PT+FLaxKUV5
0K4FvSQgy1pdYnoNeLiBWJcDixlICPT8+JXzTH0a3uDCwgGV0Jf+EjUb935jnJdV/RBqO0T2T3S2
P8EKOyWV6aID8OwR0Dv13/PXUB/ShgbNzkJe/oQJVE7stjCoHeDWVMpl1Vl94FHDNlsnN11whgZX
jscVELSTkP294sTFdYyewm6/UVxa4DZ93i6lhXevnAav2TxfiKVZpQymat9Lc1mNFDzAamz8BMwa
uZcvyEh9VKPIE11KzhbDYgKbdeThYCVqe0EavCYulU6wN6UvOdcKl5YFLyvTzJnKTykg8hYbU5BO
xJB2P77U7eoooqkmKRGYd0H3ABYEg+1xlo6SjKSNixSwIxcJzpelWWa8kO+pUlgkcK4J4MYBpbNM
uwCeoiKIGDjXuQd7UYvjFX+aZm9/bxNuK0viK0q5zjNsxGzRkd9/e3Ed35WfoGtd//W1IRecKx2D
5PM4mZK9pw0KJfm16zVM04tm4ShWSV4KOwWoj+h0/+HXh5hy8T6KhoXIX7n0nFZknPFRNvLW2FG9
XPmJWFlVlrxcgM+KqoDw+FKy0HgMDBfWADbeWbYHRBRm4sSiutqFrHCgvn49RZVcFLPWOqSWV9nN
AL/33IRKSgOEcEuBcjFSug6x4SDozf/IyOmT6CRueDMGoDm0/dHpmNoqa3frRe0w8e9revQqDa6H
BVRd1Ooo23PPL/CuhhcRC3eMjI/0q8fYsuBYrKttOz83bN4CuPr5SegUM/hYOUenjshZrf0bvfPJ
wZKAv5XGy7BOxNGg3+7ROhD7+0ODtoOYzjNaWzg1htqa4wNwPF4wtBj7Qqu+hTEqGf3siptHLra2
xUsgBrYXictTDPCclNCRagXjAt3Fa9apGyfwFlfX1X/LXut56b0i7dGOgPja08w6jjjQl8KJ259O
b4Fo+gqyN/VsciwAaNNbYBeOwRPpKc8p8kFJ18zeN/b4BvwgioyjFxoNva3iGOdqxjcvQ+D2SUX/
lF0Oy/c0vaSarOJR1yWZscv6MjYlPq93DB69wC/orrThMk2VKOArm9v0/sA7BQ7XQ0JINlS4Gmvo
yDMhFWyiexYpHfN/RvJ82/OjsE4shErX9It4YMcQLG89vtZB659cEHDhO4BHVuO9UT/wcX0ahVDp
CkFhMi9jWd/h4dVSisKkiXxH1Qtad9mSnJjgqmn/TlBg7AGnP7OHMIiA54kA37YDA5Gp3o3ZFbD8
VCwpVl8UQC17+1nQuhvdyeouQtzdjOGQKgd/KjbzT0igPYBq45bgon8EPX1mvLGGl9c7WQtqHdwG
rf9X344aFrUuAI+4RNOpQVQ8/ScY8OvtC4F91hcFFzm4z3fNNqKM0uphL/IFX5JDmwX6iqC+894d
NKgnibeL4H39+/he0A5MtRt73h0rJrRXZK6lOejEHjXPrxh3Rnwr4AKYkh7mbr5zMXi+ybXhyzcI
O23uH5fpyBhwcAN1AvLQH3oxc2NQY9QB56ZAZWnrTFEfMMHgA/HoOhtWgZxbYn703GjZbI3XP4Xr
7OJ40tip6xKVBpM/3Xz1IhNTrQyPYQy4Q1544VwfUZpEMIK50oJ0ZnUlN7PkDLW6OJ6vz6+5lPaL
MP0uoqGNxxFB+YphM5IKR3xpeEFUZFyOebpWcqXz0B8DEtKpy7mpD9NJpKF6ZtQJH83jH8KWAdWf
8yu2zchIctgEvUIlHRXOcuaq+SoVShZEwkq7Abc37zFYKcCYuz4xj/eXOc+652Hm4y1uo5d3LAjd
GajBTDfOb8oWKLiVbYDlScu8Iiw0WwA9l+aLD5keMpZRwQejBLH2Z+FFxBCgvDOFAahsot/EKzet
DFXXsy8YbMgVcLADfDc4iNPZ+ipkCwb3GnFeAF4S/ehE+qmcMnb/iRZHmk3xldjfZmVakHCC1nM+
nR25mlWfcPSvUzzaMhGTLVHlWucP+N+HdDfN24XSbXT2tZHmMnoKLFqP6UaEzIc+HmYZgs6Trz7j
TPHFR3lcxNSXbyUddODMzhqk2NKbyU2P609g8LYqp/vl33U+RFeckiS957sYxriuvb7WmH1P1rLt
PSyxE6RiW76Boq3MtnEXChLaIKu4+HUypniJfJaAoYD1DvFnJOKJneQF3RqgDlUuHJpDo6S8xk3g
qa2vBTPM8NFJ2bDEN38IoMihqqTAloG3ZlWJtRu+2nD4GOufuzLdnIu1BZMj4uKADPZVDIUafw6y
CajAMcKMAzsNNUgsGD5f3/I9i1VfUc0e7YucVHgx+Z3IcFLOgG8LtOkIj8/vjvLv8ySmemN7bu7v
IP8f0Jk59mYB+G6aIl1QSfzo+LXSbWhOIB2+725/v21W2cm70HXWidh5Pte4P0KJRZ5dVINTbHo+
tMlM70CQJY7jAta9KzoAOYE09j0NXUMwD/hOFwWOhSPvyK4XmLCI9Lvg3EcyJvIhNZPGw16ZR2FZ
hf8iFsK6tYkvjcaHCeXDKyXqcR/Lj/Iq0Jvz8pSrIlRGHe7khZw+GOy24kgUEqHbRPrp4HglY+7z
CsTT+uVy7s1QKJgWFdr/GfYLqyoIvXYO1SwusIPj/4zlF5NytXLGO/0LZKl7XEHdOG8c0V73NqZl
wvcGjbC/YAsDXd2d3BCAucKmbSitZjZRltwTl+n+RPZC0o4h2fK93d6cQRTy1jxMNem7+csBCKt0
1fiBAp0+lBQhzdHgs//Noh3r5xmE6nMSl+7nAiMdPSx2aeC+968qCdsBgdWyac9zFwKF+qW9G17/
HrTkx7LtdUHjrtHC3wmUSo2SQkix6fBz3yO7sabMRYrEhRojkF88RpbEjtuXt5gozMsNDOrAXANe
eRO6BrGsIUxoDRvDa1UCG0OtDhEnjP0Jq8YdSEy27SflmeiSHtwWfC1Gz7aMRLE/R4uE4veqG9Hg
fQz1D7xmv0OzIXk/UiNh19YZiNdmFx/88peMnZ5IZAAuzR+RyOEnwEhXpgt+L1iHSw6MqcVmhVkJ
lRCgz6wG6ZzSr7Oe8OSmRC9wK2ZysandB7dnjM96jYSMo1zoW5VMQ4Z3kJjyz0vu35UFS1LeQXmp
PTnilhHlRmhYdK0wCEnJDz0lv4glzYS61MBNedKZKdHVi4XHUQTXva/wh+8R4mkXn2Sf3bF+oAbH
huNNVF8b44U/JuKg4LDZcsd5C97BaadhsUyMirXDWhEz8FairscKSIMl+zDWSIQwFe7upChfgt7t
6VEYESYNuAWX4/oeLtescA7eNK9HCoPuE3A96/DGZBo8UgWWpOGB1DuSZphve8ZKDkRBlG2/KWt4
AXXIrvBYTt5P83EUlTSzvD1959+UkRrf/hRKgipjSWsAFMPCzGsx8+O4scsxbC4XgwFL04+xTeXg
Gq7jCRWmNuFBbzPpOgDqZgdVv+u4rShz3HH1/0UCAHZ7DOBQyr1MMl9uvYygWN0+0bHsLp9V+Aoa
O0uXiNTflV6XfRo9NPFaFX9iKETsy455Ya9bystJxLkosDNXDIlIJeLALGd9RdebUeoG6+EFXqSp
hijrO/etS8vKa4LKsEj7frn2NIE0Nx1senrixSTw/44ZT9B2iGg6k00j56YiLuOo0mBx6pebBjbW
H+/Use4ryVzqKYO+3wn0EsPPhS9P7WMLX6EdfZ1NyAvMp/Ed5v6ofqAx21jGnlo3KsvflnyYc74P
zz05KyOpWKeCTDefHYaxfimkUd4Cbghn9sV1AJeFJXbslmLe5xF6pYFkdOmJHiy3BxTSRtkg6SEo
CeJglsLaIpqxDzWGMvIH2JcHZwQPobHKUeDH57OuNq4Z4IN0ncDRlsjthy4VWb+6LucHgyivhO7x
uddmLJdOnEX+ueP0ZNu7AidLDniTmo+cULjc3TkVL6qnPtiP656lEm1CZoazQKfNhwQbiPNvcgct
6mhdF2SSWxrRqveSDZGWbCoT1xeLBf6itQScxz8+45wJxNyxoPccZb9xKJPXHUM3Lo1L57c+OLqY
o82T7MarP8cXHJ4V81fEAAU5THKPz1NEGRx7wTVsgMX32U3u2Vo2IbakS2k9KYD/Mz0W1RgdGMuC
nj1iEO2yStMN+VVH7XqMsx80u8zGvE758mzS9qkLDkFjAKSSjWQKwE1vtriVnGCjrJ2M1DvzLN8N
QTf39bS3T7xBt/oaAG/FQahtT3L3JYUKsCXQtMCQHdANpw/LPTBJkjDkCliiS3hRhpFV6zHAaFJo
m3k9faFHjx9MQIHYcMXsi8pV3owz/XVuO26y0hk1ycqVivY/VjE9vF1iyCm2T1YsIdLAFyHS2tI8
a4oeaccFRhXMICcNGEUOqUHRfRvYOpravFO/UXkIJffDi9FZhJuk+zYhYzFe6NaaKrj7DCwhy5iS
wwQHxsJTIsbuLYuNuKtJ4nGKviZGF7KBprehtsA8xCbHr4QsAJrt/TbHdw5lr42v1ZFQC428AMl0
kXWrhtkxMZ+NOw1Ymjg4+yyL/5AskP+COqvVUS+1UFQMJrG9+gtqkKI3RW71+GOWH2OdSnHfn0HP
r2eqg1rTqkOa7yFbyYoipvPswBDoX/Z8yO/ETSSc8R8z7n8gEuedvbeUD9VN6KhDNykXRlWtg221
oicXiPxQqMR7nCbD3p2IKN5hDwS58ogYDT1jZCpOav9TwSZv8CPJOIW2MySd4Aan/O3Vz3d/Qg3J
edADXqBCzPobyw5xKA+JjDEzze3P5/dO8mTQ5kvhORkec30a9ugp0TL3l1D0hgMWgoqxfsY5gICZ
jIpXrMrEaQ+1TCOB4h0s/4oVR3y6P+eQ+pj6pgJL14/jkJaGCdroC1d72s3m3qb9OOmaowKZvyUy
UevZmz89X/3lDk/DW8m2kR+kHMav+qZR4vxUHIuNyZdcYItx398x+Qv+2QrD0+co/8ryw8lMjQgt
9dM0gZlzgF9UnH3OlNxZYeI7JzIpBgMPkuKyCCmlkt8TdgHAEQ6Oj1eSfU/Km6hG6opJgwqwxFRF
96+svXvkjn/QyeY5m+F5LuZaLREovk3daHGAjJxgoz++Q0jpjclGGQN9gCLcPHhTEvXQQ4HYsg/J
L7w2KUrmP5ZgBlmTkb1leQJtPpnF06pO8BU8sj0Xli5zXi2JXx87CZwSKm2thblV0fvKyCsbhl5B
d1Co2Kz+w40LoX6rvsYZojpRX6CNwbKIHpJ3W8I8V7rrYlBZKg7jqKg1vcVmy5HqM+BYhv7ARacL
51FuFntRZbqn4sDpdpH87QFus1sbXQzF5YtAcNsbHXX3gfQcGL8sa/W8Z+9j79GSdMNkTtSIUpOI
OvbUcyCVpUyV6Ph1ou3pdgCn2JUtjraEyfUUO3tBhdShNajoc0qUz7Ax/Hp/V00wxduuJ6ICR9/0
el6n8axjPGPZA5MatBxcukaD8oRZq1lsjSG016xLgUl8O+hTkd44q4Orbrv9M8uEC7J6I3S/L9xt
tOxrGW0k3AB0gaxwFnqKrWHpSeyZS3jEaecq4jFEvMB5Egf/UUEWimKSuuCSjAo5I7uUTe5DK5p5
Y72a1LFqA4+YRQrvkOA28bNFvqQl7ufQT8wOrVZg5wzPx02/+5COgniI79VMfgfrRfbnDDWiuIVa
8iIdFow9FukJPjJ3+LBnYZ6EVUQ1t+er/LVpZ6sYJSZHpeD7zRIujGAIv+aaUyxriNMVl86M6daS
Z59wzvOaDA623eRx4OnGTdnLPuZx7WozOz/OwNsX2GVfyX8Nar5GxT+2KnR2emCoYMUFBausFpzj
ICsHhTcg3bU6NGTpgQcOcWVsFwfqujslQeopvSLnKkDYwirVGJh49Mlo7KSj/ZjE7UrDIyBWWVIH
wkYNXPhDYynn/8jm3zx6CxRyw8rOO/bZn5DUfY5hQKAi+UG/2xQChWYsiIz5TjwCx+B3uqP+aVES
nlfsRz795Y7YeSUyDEZwI3NKneoi5+eTbZ/gW2sCMJujduK1m3myCgXAUqaeToNSnsFGdqHV1SyD
34q7lg+zy0VAcrNZkGQEWCJyady9DWz7eO5f9XodtUxeFs64mqGX0zvHqr8wTrLSSYuROzLcuqfQ
uUFWzFr2YwlHKfh401jTX0VXvH4WsgEfnBmVZU1WIRfChMnDT/erY9QMsC5WCRq0QMZBeG+p1Ew9
e40gWXHguIyMVkjCxph02c6vqTafeyJ1xp8l3ToHQG/E3d6GGxSgDq6IcKswv3MK9htr9miDe8u+
JQiBwIjtHxVUmxurPxUfs+tGzsYh1IoVf1v2ihxEDTR7qMnB+rOHqDjO0OoKETwDOZ64q+6j8d//
BSjAUjk8bl1U4J3AXSd0tDlu5vjDHFG5YajyOEMAso/N0R/3OxAjCGpzSx4A9qm2jv8XqqMT7c+8
TUYmWysqqcELDlim1meFMOVGXq2X+J5DGLuT+VerR1mnLPaO9aWC8H4iPGIKlrdZYLtRwnvuS3O4
i0KD2ughfdwSlCl+uXvEXdLWIrqXlC2fKH2lafUIOx92zlOdFJOKkUGH3ICxM7i3Yunudk5mt+ID
7gxN52fhAtkrJ2se/eWx3+hXtVk35zGoSw427431YJ2V6Pw4GoigqrbtYFtU9TYEKxILUGDV3DS6
PgDsdSoK3PWCWenL5u1LVUNRUlGHklZGkouy2ucV4CB4PG+skl7RHoTAZY2Q5rjrWx2E/83j+3Ui
umsJhCUwoE2e/ceFzRR30gQw8JF7a80cPfdAQn6dnW7ayr5IQHahAW/NZVDiuSTXwef8d473oGM9
YIcGBj+CPf3YWTjUnSWX60fEdmt/T3q2cRy+/xjM0UZCME8hIxFBmT2EsCjs6GSi0GT7fzL3VgMV
Z7inrUtydi1cHWTxCmVwen+Oqzh5oLz7DQsYnnAUG8biYYAi6AJI+AwJzUM9r2NKrKnCbUUi9v7y
uxsr/ADH+FdJkBub0xqSxYkdgE9LJwlP6tqh5nyfPixoJPNQuE324jEBM0Am6lHQ4txH9/eSABxU
r3Yr/hPnBAot7/G21Twx+NQxG8eVA+0TukwHTsaaUxYLUsVQ/nnSaDPi8jud1v8EjXqPmznIWy1D
GZCF6TmRaZBtCeyeoOYOh/jMoLkLvaad38qpvvCHmjbZQbsPnwhMKrOMm0oll8WQuqDCql9Udt5C
rkpd1bA2iaxRAXTRZJqC+Zw4ji5No+ozW5JiJX8ZJ4aL8P8k8FsPuox48qIrmi5SKT2CgAU0sMDC
00Sj6FaNgITHkVjAg2pNir6oGCTfc7qWtcGvqU/8URoSPdZliIT6ghUS/YfZgwtBRNGsSf4OYvMz
UvJQFQ2ktCF4R4qdETyned2pNQEaT68J5jn9u8m35oB/dSqE3MQtRf8gdUgLYIm0njDk8InxaWXu
WI75phmoI9rufGvuS2lQMf7bCCNc9pa0FvGVQaR0m26fYQ2c8hwm5s05vcuPxgqNaRW9+nwu3z+L
y+Ktzu2y2RVdy8N+1f611AKDQ+sLOyeLiWpBroCCW5chTgouIXgesZRWbM0jqAlrQfQh61/a0iXk
B0ExNNy4bTtWrRPsBa4DMVL6G85q6NapEkucDAXP5q4dJNnYZtWCl5+81qmTp2FXVUYes+Ufle8F
kb6dP313NVmWOUgwj8VE80pAvgrafhvn0/Y1P3ozU5c/oeJrMkRaudk64TKzTqFITQOlAJJt5BeI
tTqvjgavLkCkvA3i0fmXqFKOD+/IEX1Q+uZ+a83j9GjdPBdoXzSu41oKv6GOohfYF5mZdvWNMSHB
z4auof/FmLAz4B2L0Ts8jCDVvHakqHJAsGb/7VWgIltlI5VBm5oF2xHjiyy1mOxW1vLyAb3lO1JZ
BSsbZ5wkPGFq+hbFm2ZIMwvlUoqsnTdWbjIOvjHmbVesvppW8lStSBt8qQh7bcc3Xt1ygCmbkvpz
tBMYlYaZhklUy4XjLIUfut0E6uOA8yOArvFPZpKiR3zhWN5Lg4HAVB+5KD7MqdUhjidIVjKqflto
vFJ//xZC0HvfPZqwWNjXV49SKmci0ePIVOsTZpt5PiuBaQko+et+woeAbIMdeo2gRTKd9CoC94SL
jyq+ivB0VoTXyTqGf8TyOauaPrSlziyaSdsaFHdwCC8x+XjDUATcsJBWOpgGy1gKAEobM8fkJrru
+k3j7ejrsh4K1KXNcdHffPcPmbxJ5xhXeo6WacrA4eWl+KBAbcGrC03NBS78au2JP1YSM/+YveK+
taIaclY2DVpWlcXmOPcUEiyqXpLqQkBlQB7JkUzmnMKSiABTFqjbqQUnqSu+N6VduU5NXNHfkcx7
C2iRaHXC+8DoRtxv+006B5/PeXOfpGfFW08roNbhC8fAlFd+qfS6+ruMqaBnJ4VW27kPWjP3QWlZ
r8zhnro19v1YKx2iMcRrJCptpMmNTAQxoL/uhJHqSxO/CzRUdJSSdymnBbKbIkD6Qr5ogltW5UsJ
fEaKjyE8vlWiG7DNTt1ujNmS7T+6MMkS0FeeyUmpfd8IgCbeI4qJ2KZF18XGujzMzu9XnWn50NY7
ZUPO7tzVyTmPgoLXz07yRHxqKTU9WKstroS1bLRRW/LSXkTyWpwPjJolj7nly+qumLcJu9ifnfpe
4shfoIVpaZMsZBwyqQa5Tk36fn2jYNoU+mk1j93Brb+YGG/NDv3jOMJ7+DSdjc6QaPX7WOQGrT30
2dGYn+Rps62gcKYxKq3OA47eBOzRma43FS8XlClNeBMeUXoT5xqf/Xqc6ussdt56HN9DtojasOXn
YXvsSMGFLNvMHoKUTLzVk2RqIZoynLNAdhhuvGdfol6h9dxAYENUFb+PpVEmbkcrw2c8L1IwVHKl
Dd1JwoSHvMpiEhexUcI2M58uS46DUGfGIChLmP0hE/vWQQCgOmj0D3BpYj0sd1RukGMXTwET8b/S
mC5DntiOGkhe0Z4bR1Z9/hhmfRthmritdwqaVaxl8oy+QdKp8P69s6du3hRxgS6zTQ4B59omAut2
ApRWhpk+m91OxA9iCsMMZR6rWTWJ5yVM37HtTaUPVV2dVzf271JAVjiKLuN5Lnv8bdkQKlM+vZ6a
KRvxVpbUDWnUG1TnsrGZvnOrZ4mjekjMtTungvKXjTbe6ld6F2vbfLwWe7bESpxsbmbOaDODjWWm
L9D24971qg/szzOYEbI7BfrvdRAWUyLC4kLWeLEtmTpOLftkz6NTZ5Jz564jyu8rilaagCkhC+RN
oZDa7wtL/v9MS7mUKlQeZJmndhowBOysl0DXnvzlSCWd13RBRqcYx8njo1I8wHzzZiv1crSOcs+R
rdeAyrYWbvpGiucuTLxUUBaetMcBYN/C2qE0i9yziPaG5huxb6Omh8f6CNFR3SZMOGQZjvVH5O1j
Un/8aT883OqiOliv6BpahTKjl+7P3LNUOQ7s7dHz+pHKTfTBjPkQmkH3Z0gDspmCluGKfGg6cvyx
HRcy8Gm0v1vsJH/gt74SosnbGdu16akxHaqFHCmt02RANXHWjGRaeTIdi84UW04LrFLznJ0Xp6Qv
Ku0ceVVCLpXUdjOhOfvne9Vo/IY+e+GxiN9vWtMjQBjHzW+utiOPfcnBnPQa0Y8vTxoPDbpwgrnB
+hf3HX3ae+urWbmYCpkpPfWuDG3QDDK11cTbW+ewEyfavFWdt3Omk8QOr8RhA0UV/HkyZSvKIjAT
cz1eZ7dwR3mJyTaHhrQUUlve23jjGOmJH0W5mPuf6AFmhtaat4kZfuQKfL+kCw3aysYPCdrOZljf
sluhWMiO/WiyD8Aat7BBxXNrMiVMH1+kCtmUlAnp4/T7mKbiBhq/BN2GheFg0xWdG5ghSpfHNQ0m
r1gXn4ft39XMcVQ9L1yC+7H2TFpyln0P6MRDQ1n4LqguKapPC73HwVbZIMtDFCth/+kc3s+P1ujx
GX5M81jczsyhl5CWnbfs70lkDptHkuORkskcgl5Zb98vN+t1e6ZFIgNASv3NnVIFgU0yUYF2tVmS
i1b2IDRB2PMGlNj6j4tSqv4opPAgMGTn6p22L9OQ6JNzWKubnbQCOVXAtV/Zcaq7AP0uZ5lIzWOv
881Ps9HpaXaU2+d2YxJRZFbriQW5Gh2bX8s76bpbJntSmBrlRf5r9/kO88W0zcJzMCmEBsgLrZaE
6PnsSYcS9GAkZ6ti0t7BovbQgnfdZ8pBAN06zvWEkUGQG80JLpxfwS31OsMttKUkYF/3KB7nRDFf
S3haMxCinBwkr0siB+U9Su8MV8mmzdtiNYeUag5uhpzA0A9JQy49ewIIjIFgRkPEdloIgU2l9Wsh
3wCazgw+wDRtHnFOcG0Ao5NTtyk/YFwreajuxERlQOBnbgJtNJ0Mb12BQqhFU4f2t9C+SpkIIaY8
OpPhBMJU+8R/1QKA22xWRtrpAceXLBzgkgoJHqXmcRG3veG60CPEngm7m7LknEegSLWCm+abwpX2
fsaMhyul+I2S16PCnYv46pWpDgG7bUaQi7J+TEKPJw8RNIyfO9ddXmHBmN3Y68D5+v+Wt9KL3l01
Z3GbzfObK221M3zjRBWHT6bXfqGauNQUWvKmy1enKWeBmsfvdFFNNf05ZvMu2e+Blsm7gESc8K1h
kuNHIvhxjKDZP4QCAIdmNsRNfmh/ZBtGzOnFMjeici8s4wnIdUBrjNDmRwwLNRiMxsyS8dqekLjS
6/ZEN3qojJfKWkdL/THOZumagJQlQ5/5ijxjHjWIv3cgyHjSQBvr4Uexf1vzPfGFWC0zvpcAurC3
pmZMHhoE/UkSfxUj91pp4ur4kt2OkKBeWT9hfV+TW/AUoSLqQcc2nq2Qmr2CxVgCqYy/1/2w9jSx
KLmswNZ+0C4NpQSAiNpHmuRYwc1FTru7VlHSGZaBd0LfjlgKb8Z/Tu8rQ0z/Cb/2rnW+fmFVcaHA
kHdnd3106j1DyVC2nPft/uz3bcsq4IDmdACdpvyY1pVJ0/Gmp8UpebQdJopCwSb2+WdvmF2V22dD
Ul8LeeoB2WQWsLbfV880M0hbyRP9YeD2YsvIBJR28t8nPysfCan8N9VZKiYZTEzZsfd9KhT1g8+F
wW9yyqhX74EJmbi3C8meG3jCRttsRLbsSkXcIi7p1ZB25AiyT+/UteZZksPu/UwBnDO11/odZy5J
lMhXVN8ijy9aI7Bf1ZMyrc3jvHcPX9q0k+GZga4259RlFb7ixCN4HY07/t+bwPzzUZF6/4tFfOpR
GLGxj5Vp5LX4oh4Ok+UgZDRWnqYdk9YezCG0jlznkGQ11lKoivI0p/yXbFCTTmcDnpTeXn/kpCQl
0BK0Bl1eOt2Qq0qhfVBPLL7NiRsufEjJ5b47X40rw9cuXewAAHNLmW8eCy4VIT0xjn+S9T08j0N5
x4W+DSfyCua1dyjZt2Zx3PU+SxhplFdZfa5N6CctIOLFN1cw5qsnsYKeBJ+sbky5sRtKczqtaoa1
uygIqp+XjAmL1gVxiY6OIpDhPhKyZ6cZBVxGVq1XOyN02S1Yg9WYt4kiPDXdldDwNQicUQYm4Kwx
86yi/VChRBmJym1epL8APVdqhWTcf2oARZkjUv+Xnks2YzebcDUngqPVjpze5mQtgaL3mSLWABwv
pIaMn4MDJl5sSrznOY1rYdiIfuxbrhpQyGqkaWPDqr2Rki+J2czLf0vPnBmq4ngITFlVM6IZi2Rz
Z7W6ICL1Hv+ArnODzLKj0F3bc4w1wRk7vqvmcyVL7COp6x4PjIDUuqXPyWVzxWw2ma0BUbKxHPU+
iRBA9vS8EWzAiwP430vNyP/mmJhQSltr8dD/GCwtpvCJ2Gfv4Er0Q4TqcZvqHD5PimCoY54pTaiS
XPZUWpOb6IjKKLku/Whgv0RvAmCI3z0WmmPI549AXPxaHsUZPqMB4m6tqMH2tbn+HkK1wQLLVHXG
emyGwUxe44VhLO/i1BqweFxj3nir9z4w/q6Fk8O392RZ+ANDSXw7X9jZbkKnMttlbHtyWsSkSYfj
qisB+NXGwW9NpR4os9V4Xp1FadQcuOg8yBQXcF0BxhbFTTkc0AfAuIzCP7VPzaXKAqhAtxPA85M9
lNk5q0wxtDE/ljogRt0pSYnvwZBlT69/TCGRwy0G6rBhruxRYmgVpab6sgHy78Gr5YTv30I3XDfo
zfmMli1lOJmSJEBTyQOLxcSn0/tUiSFEG2puU2Nkjr2b9anaMK0h/RGBBEGXEqGE1UXhaA6EA1Ge
wN4StesKUDRhn83yR6BG+B7Y3Ka+J1WI2P0K5f70x4nNaJEZMDDVcfV7A2PE9jndTiGCvfZjU5yx
GHShh+RYVj6XwuaYPsBRE3zDQibrL/Zj22tvGMJyOge4A8BQsif8wOyfzsPOTfNhQUK054ZnHzVy
3pFFognTG79lj7aZzsnQlySsKX+EXHnrFykFUb9Czf+x7PTR6oHA1uEDYE9/pOsRvp7p0IDIo/UF
B5AE3oAdIp4dbs2+FSMvzcOACPxibUdZXXJtfbC9dZGIJg0UXb5nZAp+j1yiygaD2GIwBnmXtGy1
CuJatSpHTAWSZHnSBw2tD9H/X71PUxdQ6Cl71k2SI91ttGRsqZwGiDQkae7tZinTHC+IL97A3L9n
9D8LU5VFPYztbFUDBIMCMlyyG1D3oZocRKf03NLik0VWD89aDpCuL4mic5gqFy/VwoZPtIit+Zaq
XfJRqzimUpQbJdtt8jEX8+da6dyVjulIq6Xl7bM7TfCrupMb/OuKItPIT0pKSxj1BvIi99Y97dQt
+SfoAxD9coyh+/K5odjo3PKObcpYwiFpxtFZ0G2BZo7gytfPQ7eunXqbRW/IH+bLVsuFUEh0fnJ/
N++fWf/BKt88N6QwMvXIvSkMLZJkj2UgNNaeSNlul8rlPwRk1gNb0CXrNfOLifMgMK4RCrXSsMN/
2bCYLyg+Va9c5mSlVJ8Q2lbybzewRrazV7Y9fO6RT5eQuub7h897DYxuqhetnCHEiZtfkDPI57Ix
I3iKbgQ4fRwdgws97aWx2L1jSYui1KJ6yF3CSrjo/jX25GRsKzoUxmAKYaXqC+dmmLGwtzfxwcTz
smGd2EVrHUQg2oEHuU3pUc//scIBoK6/zXGIHAJ0vtMXMPMLkSPvKSztc/Z/B7vKnbiX7Z0tK8Lk
myBpqJHS1hOA6Ujev+KpZr4BIcJ6hcJPfFem60GnAINjGsRWeQtmcz5M0w3j/nt6q+dHwPepKFRd
qcTdRjTX1kUKwzuwHEk4cD3vZEvC6nRAWn3gFz6uRc54ssu8/0bHM9xpJybxiRYRw8r6lkKTum4a
EJihbP+M3KMgexDSw0r9adlUUpbgdAUyYQ4zJvUXLgzX2FXM6l04SE2gOiuud/EtYYsJFDgJtWxV
52x5B2qxa8JiXbFBd99rBp0a0JRWh7M1FclSmukWtnVC1vGD+7Ekvj2LvBp2X7aPsP49hLVjhOcn
5iRn3HCCEJQvduPwNU92rzGFlMLECwJVcIe8M9DLOnEcv2vCp7VfSQOfwGVmaxCWnAQYGHEcULOl
VqbOec8Wdx4hVvMnxURBpYS2hqfQkcmnUCUNqHzpFSGLw+hwWZ1cFjkSRJaNPo9Usti8k5PdF1rq
N5KrFmhCF+2iUG+nYs2RMXX91fyYXfudYCeZEVSBU15jc5qm+RUw7w2qTFysJ9yrItWiasVyBA5l
atNkIaKaB4u7j/bRoleLmmUKifnOvqzYyQmhxnM/I7ozX+NeFAN8HBYmyi2f0IU7Z1MdM4flRX3B
Ijgq73Fkj8Zor2tdqg4ExuykewPQUt53W2d0igA/ZYeyJ4TIDd7AWlRs1H459IKdw8MQR8FWsqDP
lmErZ5xoqqETVjThTYgnCIvQaFtzL8GuU49baFVSjHYmHjArHOBy9gbjEcGAo9dgx0H3YNr8cBhw
kasyH7fe/H1eNoJbyUM9ZErpgg2Zo3Fq7k3Zaq6pvsbAmNr0vABx4vSr/TP3512IGr0kmuuKHHNY
L3tqBYjeUEZnCgXk4lRmyEf9CJIqAWj1/1gwbK2oP/6dWmlRQp81g7xQGOzLLuKM59FWC5+VkD2z
aaNuIbOXNV3KVHoBbIEnt/BRBpGpIJ1hgbQr3LDhnmsDgugW0aYNcmwUtbBOmXu+Hn8dTovX1PFA
X4fmq2+te3DyFIwSfbnCGOhAen+lyll2XqZ5Yb3iMy+cGRrp2/EcS8o1HWZzZFbrVbdL6sVb5rY7
6OlYOyoVIxAUxGxXDNohltHQBWOvgHKGgSnRLShA0lflbcAlA0H8H/AfhmMBgjCz+Xg2GPltJsV8
VsNJc5RG6p0an3rROgfaPVRvl2obDQQTsumB0JfW3fO+UvJ/l9yQxpe/KimMJyk2GnVm/E+bayxS
h7F9G99FvvTcAEG4rJjwnrguQeP5aZZBQZppevxJPQb8ZKCVS/D7fKYsWiz6kq+d6cSokafw5imo
Ge5D55W7XoEJDfaiKQ0fRLZ3Bf7g9HbuYF86m4sJW89jaqtZRgx+TIUI13Rf4BW2A2yJzFz187YV
rhJfsSssOGiWC+AmPbw1N++/FGg7LD66X7HW4fosWQhm1buV1Fhm57dTPwsto7uXrFKWlpSduhkl
jr1IfLMUaBg2GqjQ8qdHViCJOXBNe1i6GkhjsPv/3n3odb0ZO2PP9OkhDwYSgvySn8S69ofRzWZQ
t396T++iG0N4kzY7qf+S3AHdbZYOSdEbvmUZTGqZjV1h+uhqpCUFxhSZ95tynyIwX1YgA9SXlHEB
dCy4KkNUCWUw8RdYREwCjixBA32jtACfSQJXr5QgBu99A3zFd9G7sNbhV0Q80S465DsC/I02w2wW
WAathSaJn7saeAvG5R9U9yUVqGbo8Rb6rHP/iKC02Ume+cP8tMov9iTV7HIf/jFqJagb89DYD5jM
mEMEu/azk+/fntRI7fWJPXDqc2uc26FMkgFfpatTlf+YMbVBwEwIjzDMmtqKnidm7PjKjZy8yQwu
m50TghJR6LfAIj/QaJ2w8OmKeC3rdkIxyDUmv+oLLM5ck/zxRoCpg4U6cvDhBLIMk389x+OWvm2J
VY7Oln14FIYDvoFG6Qu7pOy81V3I1mv4Q+F3cDrTdq4MHDBEPIAUnBHugzTvMEFy1GZBRSC0/VLK
NDQlysf81hANFQUqDtMB1nypiCmG3wly7KMWuTXE5fpUq0k8jHnKPZ26rl7QVJsPoPGc+e7kcoRi
ruIYemRcEuZUJN3p+7++AXoQxGYKHau/TwLBkcYKkeFvOkS1TOFczHhqVYbjf1LNYxzzWCQg7w4L
XQCXiemZBRYpky1CZpRUopYEICZljsXfMDyMgNlmD1COUaSJ3jHtrmSMjhNsk5XjGyTgKrH99ubd
sK/FQO1ovmLzSDA8kR8XDHK0eFqGQT4I0ZNm2j18IXBjLBH7OKgaqUrd2dVEASlFo2LfIXLYvi+4
9LR10w0mD9R/SNuozHCGpDNCZWi9CuYpaQtcHUCyq9chDFDqGvMw0lyH6UiyUCTds+u4Uu2ZLam+
YBbpRNjWrBSqFjS/ktiOFgzTYaFsdHYSdjNOGnHXcjHODAaW5gRn/d5tQND1MtU+6fD9BKLv+GbE
DYZM99/pmdEjnVKHIvJNnCb56fCoWGMJfHxqsGLL5vFWLRK9tMq521jZK4bnmdL9z6/3DE5Wk9+I
KvWm41x+q6kr2xUs3tUryRtYAwYfeF0+gBEmFiQHm94oYmxh7LldbNLgKSIb0w6HFVZ7cf8CskED
cdhGCgZcCwTUQK7mFyWnQVwELnDKb6AU74ZpYRYun/Elh2reshYbZcdNRNvA73gupemBuLxh41+w
9kKjl0qIkaejg3KvUJ2tk3qguLfvfW/vdrT/vMB+kWZO6xHUJMZT5pAIW/fngeVoeHA9Ji4PJ49d
mLx3/iVmfcQ2Do7chx4m7VR9awMrfL6lMeuKC1spN6ATaaIkvr1mKtgPfb5AE9ThN1Mxpznqtxgn
founAC0If3Eh6POzRQnXa72HV8gFClM2w6cglPOe9CRtEExQFsoupG8fAWfy0CiUiF4gMjQNRD4B
D00S1epsPu2Qvge/4vXRE49FLE1eolrvODQWTlpJHwckqvvQqS39syrYsbPwCeKuEtXzWDdR6jWi
6qtKvyjaYVsraWSdscnAWwj0ah7tYxBUREeQvdfC5y/ZNbdgykijJIvephC8mmLvs1WnkyKYL971
10B04g2bxj8LPPK0kgeMWpfAOv1D+yaupuWw8hak3dg1bGfLcnOigniWq4L5oWlMo9YoxxmaN9YH
WyxNgeUJUXtc7X6CH38EoPvxi2KibF5WzlTfYIeA7FXygJaC8+oQ/+Pa/MQXyKzJOzErZGDnR6fr
E3y0DkmwMoIi8Hg71E45ABhM8rSEuqep2gGJGVHN9wH/JPOkOZ4Rs7yOrOkCUkhteZusZQrR/jxB
ywUvnO0hi7+DcSttZcUhqMxm2A6JSneBJvIZ9rRLn92+ytG8srMhYUozikmtXn24n+ROD3TBnneU
P6f/uJoyvaMpBut8P2lh3UZePUPOslLz1PrnZecPBhZL6/D9yEsFgWwokQTeXxrzZP+KaFZ2eWiP
9QwQi/EZPBgnsRo4b34hYV/Bd79NEjvFXEWWtKok34hSO9qW/slYzGC1AxaZxt8zeprDRibO6KlM
KqM601qlFVHxG8dnhPREHCqjyYA6kM8hq8vb2XTBLBKsjSG+yrAqEJysPrp9zzG6ZMdp81C/0fAF
htDfABhn8+FaEbXpsnt8/IismblHpz95oWMm1QBrXzjef7BeHtDhenKS2O1H4DlCb1HUC5VjDiGL
f0RpdXz0uET6Nd9ZBMB9/N8QuNd1mIQwxwfzedE+C6MwBdg6hQvgxOBXGwdUxtOwOlwOSB21kCBH
SwmPRHzZ6GNPILcCLNWqBPC1lSUIxieJFQFUw43/L+8z7rkP1oQwBYjkhnthPJYcrkmH/fFIa5Za
GjwmtSdYUOohDDRTKTClpcsqcCSq4Wyw26K3gBigZgwL3ZYfvwDaqQZ7nOyv0cAD680Js6Hmtxai
H5iOblj++3oNwQBfopdEBh156rpAf1WUbpf0xKRool3KA3hVi9POODLssXDsTYKlzbw5SjuEiUWe
MxA3r2r8wH93/S25z6O+yTMkLlAmMmKZ6vF3WyIlSkOpXkM76hSzgxJ4KGORADyX/ClBgj/xi5J9
8zw9w6699Uq0zrJRp8Mg5VnLeUPc/X0FS5dm3QBmC95i5b73PheKFa6F5HfLYmzBNOGqQuY8t+3g
Pya8hzOE19ehJ0IIj9o9+ACUDKrA2tboktaz1LGh1wAqbrDyqmCsjRCGtja3JDFqmqGnnJipnAy5
+bg/sMKNyFSv7bwSi5UCa/J7ZIlwWN3NOdr84Ss4lFExginvf3q/LU0wpew610pREB2lr6N6PKE0
N/PWPKJX36aLNq4WRCNIXeXcbWmQXdj3/7luOhO//NVxdR6UXWPcyyzRv36jJAVn1wPMvX0MZ5YK
mjGlPGrqYACeFZJf0d8xTNIKwpzEftunvVWjLJ+Ch23dpZWi1P9QN2Q5Z7INqn/iIct5iGrnmEyP
O7zHgLcXwB1OdOOqxCP6N7UMtJeVuAD8Fl1kwVf7kb5NiGeSwJf/5DRpzg+c8zBn/qa2UsHk631e
d3dHSjOfhDcUH0eNnGb7owlMrw1HVX55IdKsnbzsSbkli9GXYL5XwK4tUBnN/PpvrGF6uFhOlUkb
RrshebkReDXKvIjrnGgrFiKMtGk5yy1+xiInT33bN/0T4zfHRjFTyaNjQV17Fn+inoxMVlsUhf/9
St5M29h50OCOu9HJfdF7K0cN3DbT/wBK1Gr2+l1rxAJfMAqo30+8VnIbE7eqD2mlH7vpH3DhKx7W
4xxRtwJBzp0jKov6/WSbDMQvxHsl9ctLE5pENj+7qbAJmNl8F8L7hrJu1nXxHUYafbXgCJS+sCSs
ER/L6P++WTj0B4eurRNZNrdixZCFU4xGjyFfOjMKm+wyVOUa5SGeNx2K0IzuvhNAJpe75THq5Q2K
jyi1hcsBjCiZovo7cv6if7aKf+rZdwnrulNYJujHyym0PfbaqXrQnZFBKcJjCRuLafL1mJBH315D
vvP4dv3RVXrtTUE1NiSLE35RN7dbnCwQVaIdXkC8jZIldY4AIMWUnVlN/oVW/KS4XAgA3kF9PIv/
hGVruAGQuZhF+awjDfOFdfnTH+hy195OHwQoAP1FcrMsgRq3Zvjh9/lVw4wvOpT/2ToF9UFy+EUV
H3pWekHrbk5bV0+bSqk24H9WY8c0JcQbXeT6PWm0KfcwKT/zLEi1E9Qplj8J30U/2jvH2psI12GR
rcav7NNRLeswpoXV61a6hJs0y3c+pwyRyRuSfgsKLKRb4CI3fzz9H87CHlH5mFpnLHaZPReggXhC
vaE7F4Pbpae6PYQU3RCz3RzFtFzoO7TZgtiOAmZqZ/KE2nrkms/sJScawQit2N5dxsoS5sjduhNX
eTHgbWP36zAp/SAzkUmQdubFZ+dl9WUAygIM1q0ocb3ilgz8K9E2bb2eWqQr+SlePnCLu0iobJlu
hD/pmCf8s3gkQJadLCHtfZrwh4D6I9C93Ukm6UZYgsrKapv5jKUlCJGw9shiMFHuBmU22xDRqeWs
BNKFYueNddQE346OGRs/yV73sG3L3Wa3DIc6g/G/S/p9bpZXsdv6Lt/2Aij+gWKighqOjBeryT3y
j5+fKyqbtwS9l0WDb7mttFJ6phZ96NP45COk2WstAaVc4bhMxPSIazIoS5gFfgIPREtC7sQxJmMK
A33TP98DdrzJ+wCwEHAT+vIvSpDtdr9DY4ziUwlA0awYiKibf5rqKceY/gLma52sFBJO0Z1iPKJv
kLL4TPR6ZqFftxw0OUwJVjt5NVF4u16ybf+til3jmO6uMQdEuXeBAQq8BiINmzPz1BOm0cq5oxFA
92KHcCvjfnQHiu032mRy2sZ11sr3G/Iv3UuY6KpQeccwi2aedr9yC1BOpk8XVc6w3O5SJxgLJ1Ig
943RZ5icnq7o5C8MwM8xRu8EEQhDIM6h4yxdf1XfVOQJ2Bp13SWgcEykmrUe4+xh2a5ZBIM8r14Z
nj0DOWuCtC/l/+I2y433B2ditoksxSWywBOVbD2paY4koQ4pZorTthFY/vgX5lFO7BO+Z35Qahyj
bzldT1YC3lr9BH6mXr2anxnz8GT/DDb6WECxxz4gktuP1SNxg5y0+N8P2euUFSdRXx4y8YZ4acFe
ZiBq6FXEVMbtCr8cUpSmjBSa8jFDzhpGAnsJXICKpcQrKsmlwrs9Dbc95XLksaBwd6gajv9tuH6B
RFiQuz/XUsU0xvAKtA5WhT8Zxz5I+c6Amz4ZlpwwtXbphDRrT1arcSJ0Q/X8Q1xjitQTfgskeYQr
VQu7jn50QMIUggzl/b35qvONxvbfdgD1/ew0EqOZvR01KlXdOXltf+K8l3VOlXIZ+Y4lSUgnaoNu
zVV78g1zN973mhwE3N24TAbGZtKxLvtVq/4N8gIcElOEWB1EtRP2I7PAeS5GjQ15kMznXsOdujBl
DiUCcdXJMQ1YE4E3nArShSnFiNZbQMgdD9RYHwMaxEwLMLsWpKhejyePNZJTTmVGG3n3BOK/Fxym
VytoeG37XhNzIkIlmtM4ieeD3IZ0YoKNtqFnJH6Aya1Dt7zObstNn9IA1YyThjs2jsXiblJuUvUg
dVUOG/jXNfUjsUhrnt5BoPn456Uso9S4rwAn5cTc4/dBq8YrlronzUZh48zXsaJjWPjqZyyWrhy4
ZZiDA4WxHhM4ci73p14uskXqTgRU+Yl6HqlCEw+ljTS8ZWVlnMh7Oqll66uF/+OFCiv7HiT7guFt
vjIa+p6lh1r/nozp5YJqXKUR0kVUEKCe80WCMJxQlTK8qACrYjQnMWo4m8oIxTnY5esz1mc5Lz/w
IDgB1F0BbxOVlmWFFDXs5iZi/+pdYvtlCY3EAF+Zu7xjS2qGyz91DIw7PAnNV2wmKVfwwWTjGaaZ
YeM9Bxk0xG1ZSQiw30+QJ9iSXbnabehf1TPKHoDKbRwTsZJYbFiMPWv67WSKNWHh/0vvQ3VJLrtQ
wpGtZ5x7Msh5Bz8UP3AdqS5OSK+4MKM5Tnx4VEakt2j+Ff6RcpOB9G8qfl04ecRdcY4JaIda+LzH
v2vmArULdMpTaWHrGOkN7jGE2fYDOqC7Fcc/sYknd2B7M6C4N/EFUudTa00BHxeaNYLv9qssM/zT
zuDj5K32rrdwMUlzhka2qRddLo1Vz7G91t7FvjCA67nvNf8hJamdx9qBiZ/MEswfSICgF0k5V+ue
DFc9xsVV5IT0iIwX9rvlpevjSNRBIGJOntD/vxoGTEde8HpzZf8zDuxoHVmdU0IzvPpE3q0RhxNq
JQmalcufBgUNzPvqCG7DK1u78sVFhiHLhGvBHxUKHZFZwyAgJc34BYs/mibGyQ4rrqCYAV5yX16z
GLbabbng3BTl7O9EObK4ECl5Nz3Bp4Mv9HkPt3d2gG/6ZpNi90fWQgnDx2XuPh7WdijBzFoyCQ5y
xhkWjF886bgbR7j9oXLsuFMXsP8Yk9XDTPp0RfBnBHIa1DHAVFlTsWuar3o0q6fKsM2qGRalC8C/
Py1T6OwGvN8ZKCEfockDrZdYcppyotAB30khlGo5e7iZG2s6M+9ANjyBj2t6/pF59mhNThk6m5dW
O3gXTqaZphXZ195hbGuUG08a36GKtixGFgvupadlSwymUGSNdqMlpdg4KH+2j2pFFfp1XIPYYOBI
DATdzCqm4ZF2BbPRIzRBhzOVYRgn650ANWeIzB4uKo3cy51RG0ao08LUa4uvDD32v9cBSuiiTTUq
rKhiL5C16llUizU1ziIy9LUojadT/SwoXD3NDKEBVu1Dn48Js6efuwxa965+mdrbpFb8CasKMHnH
xzMHco/ndltHIvFt+kE/WNQ+Hr54gbi9NFdjdgONdwro+5spyCDzha3sMyd6ArXhdMcfhf7xAZFN
S64cczDkxZAR99L6fU8dwJREOavo7svWhBSuB1qhF3T/OLpQgSTcm3MFMSwuoi429U63MwLe9q9k
9gdcToQMeAyQ9IA284N0DunxcOlfEwOr4kiH0QWPJtGb4BsxEMUKYlp/CVBGZ9xWhtnveYFW0y7G
JeQEy0pb+IhO3PKlePmxGAuDRNg2Tq+GJILyM891ekpB5HCdhUpwkrABFTdzd8cVoiZB4E/dTTsd
Iu8VtpIKZ2IKOe31rmkBWatnAY+aBSxhGu0z4M4G9hABEINFjzY7qS0UWuzum83miM84JVnA4Mtl
x0ObfXePrDu0ygrNnXjypzk+UEveAlOhvkmQxMwfQKKVcGc29HJmDMEA4Rs7xYsgFi1KpoBEREG5
42377uPKLosMnwcXYqeNgiIr1oK1uxW5252ojZLAovB5nptrJoYIqpLVdOIyRP5qcC0msTRnatCw
gvSwXrJMImSafhwKIiE0cTMq1wv4XZFsk0JL6qYSKFNB/lObHCLnNgBk+qrirzl2G9D+Xqm0Uf9z
VMsOaQd2v9b5CFEIZc1PgpnpeMhHNZO1VbNn7dUHDtPjfBN4ZRTlAUCaamZZMgsyN1KAZhp4YO9q
XrjHuGL+Ih+0D3Ef+e0EFeXtxOzg6rxsOGgV9SA8JOG0XxWbw3Dv5Y8Mq9Gs3fzt/P2AUGKDa7Uv
6HUuLAQlE2gvcDkfcuYOLS59BZTDCef5Mun/IeyR6gXYkZjthgA88UpujrxFxZtQ1maugphlQG06
ETQG8ieLnrwtUZWirhQnKrOOnk3i6p37S0xSGUrW8htuLW1Srt3MAlEyn1yLbgeKP5Ws8MR/iek4
gWInksMIbg8HdeNikv3fRKjzTd9Aw6/a9K7734t6gZDBz9b/F0tCj6q47P6nGKOxdtLD/qKojOIJ
TJ1dx6iTsM18z6dfIEKg4PptKUtVgUBmCbvIKTc8Ik4bKQKm1C2JCN2ha1viO1hubY+dcnmg7f0j
XpWvYIlL2rvRuDANTi/fULmB+VsnzG1UaSfGVIbGR04biPUtP1XYAfM5JUay6GEvmBX8y7Xzn6MY
PlYxHkPicnZNy5MrsSPjTItRE9e0jnTyUeIo5Ob0KvN2K2xMRkxd+Bs1wwRSV1t5fK1K3rCQJQdv
+SlC0uqPSe7ESwqI04DkSxltVs2ufXUWqHwFZL0sqeKmwcLBC9RCe8/Gfl0lkTV5XTc05aH987uV
kXHltgBi7/OqEpUFOYDQePN1RzcZoGghbH/Hz0Wp9DkUTmoI0w022faTXV/8zqR05DsxPdWfL+us
XkcAiQTITkfESrODAfrqDaXtpYSS4vrhafHKHFUbDwBMDW9jWKHoBryQTFqV6AxWvRAUj3QUNsZx
BwusPzCPOhSObthy0PkO+YsibYzMtiN7Zt8SpSDc52lSvGHFWFN7wM6A78j8bPQab5zizjUircgE
wvE5BoctEx2AtG2HnyttDmJXWW4ul+MVm/5nhY8IJwwlbkCBSuP/LLmkZFrNkxXgNg3rdmzxtg3J
xcerXfuWbn6PfamqalL2+gQ1ddILClBtr9LccR+ZPmAWzysh8MiTB5LMC/lJR1/zC7NcXcUdsjau
qEY+Td9TDkyTRGQ9j4Sx9viyH20tvl8v0Loy50u2XasMNfycXOW5h7jmdl0HHqSI/s+xRQvx6AL/
Kh4/rN828rsbcs9WwQwH/KuLQbjtgngdmfTYKSlw2O8xQ3W1WNCAZVEXUKOXAqrdYfvBhYU+cZoi
Yu8L5u4SoiKBlkkO7ZR+WTCdghBBGh6H7lGvvK0o6tIQbGIUXsZqpZP4CUTXEsBhXjJ04fbiWTCW
T195I3a+ilKEm5QumYboD/OvsPGAPMEWY7P3m8sbbIV7nFZ/lSFVaNAmlEsqkfGUcB8R1h6Ziqv9
PM10KP0e+0vmRZeXD+0XXjoON6d+V5elZgHU1/mzwNizxiW799mCpKcnPSugDamgTAeOhD94IGBN
9hz0yZ8RIULf6osuj2/skGybiWNypgS+w3Fj+f54+8TdwwpUKl0+HqzzRt3x4u04RmV8e5pYSuTo
/RCoSqLsOAiJkS0zcDz3QqM35/CdINZaL0YuN+jFF6EyWCZ/6vfqM+3rM9yF89Qthi8Pc9eDQ341
DOjYbTFkzyLc6JItFu1ofQCsgCxuf/UCid5JIRgZxXd2ZrlfNzqvs64+QbDLW32JMte8x9oAHmVU
auL3jRUJSfMHCEcrwT8zPs0TRkROOIhCU5VhpwVmnghRB9ZjuemlDAQE3hjInYQP3xZvEjspEzIm
+7oXqhhTDjfCdUghK57oCgiLT0QDqOngkCS7/BcOKnKSySxbYGPeWhYuT0n9Ij6An4vW41ZhF6wh
1h7x6CXFYbL9YSefnsU1OLourJo1z6kQ66qMKLD8/elhDai8jBjKGZDYLlqq1Qd6XVa7oq4Z6RKF
n4FBeJl6aZjjJG6AOzAtQq0EpJ+9Juj0Az5Zuq2ZCIOK6pyz4e+h9Y5/F81csbWzymM61y8Z50H/
/6MYmfd+wARmy9CUZMBGUH3uwo8qrTCGtbgimaarOhDqew4HL1s8u4/qt8mJnYjwnYV5LeOaDEh1
ATOyzisN74wp5JHmHgPmgJSVGOafT1DMgNsaCXHbKPXnQ9/5KESGrpquh5mzTD1G7A5W6K8uvSlP
Q/e9Mv3x65Ak6a7JMYKGWLze11brRUhmGLSLBfqL/JCZqvLF2Ob9TL0ip7GpMtBc14rK9EVUfWaP
x45pu6D8AbIZEu5K3BFawO7xh38gch5XvvG419E7oJ+Cktcr2VpY4o84+VDam3PjB5zWMzksaxyt
iZDSHuklcb6ziutLqmXD4imyNCBdu+5q5W6p3ffGvJt/OkA+DRGOk95p6ncWzytDOVshGJvwEoVH
NXdRMDMvVl1kJGb3PnRCJJWWAKkekVQvalLx+Bd3pLINs3LUziD1FdN0hLCQtTEz3WcNOBGEcMBd
LvkV0skAHf9gzED8bxWQTvFCREQmNQCbEubTktk2rlS7RNH7ghmKXBigTGsU+vh81L9u8VmsjrLY
8pSmfBe+2pMIWKIxU0SMGvgal4tA/ui1XkhiqpJ9D3iKbwK5Yv7l0tcwvsVHt/m/iEmWMJ4su9h0
JhLe4uok0QkZt/fgr8YyQACiOOAXmiwugvXPZyUTTWp/rHq8zWs3w+lUDRL77M3Y3dSDq0VSMeBp
tPp1UI7YcIN2nndfqO1ic9CxoyPVrCnVTU82tbe+Pk+E9M3QUQjM1c87ASB7VRPPeBA4se+iNDPd
oCwG6vmfM8yj4UW95f5VTA3M0L/DM4lfODLCiGKTxUvfhIoufO73UgPnMhkAp7eMUIk0yXuX6zPG
gksZ+W8cxqIQKWBSzryH6o3kMo+1axIY6RK/SNFF0uDQyrXde/UqSb9rTUehCzwiXeQ9tp5yKFAJ
lfBylXaXn/xYS7OLpnGdNj+nklEJ6tdDq3RFiyAM6yWIdAmJG6k1OXr6JxnvUGk5z53udJNQvlDo
I++VE1VqJUgKG3666ogjVO8TUL4r/wMIiZEByraNSwENkvR43Fm/cD6BrnOkZeP/VQ4c0G4YEDL8
th+lydQ1mt70dudKxRyCM5WfjkRK8hWKS6pkHVNqWXVtYLQsXV2ilcQN/TmnkHSGGVKbo80BHNrK
v68dpy05NEg7WAB/z6vHUPy3mY1GcKUwz5EOgLNP6dgtTBlZ7oRe/h8oeo6ZXc/h4LOahO47Ztso
Nn4WcjeIoj5gnJtXtl+/wROTp90rmYCk+bPagH/sge0frsLrwX45+iJ/J3GJWcUkbH7P+wpmbw5B
u3imnT7rVxFB6rds48/InmyHucar25NjqRcwU8ouivydtMzexg+/KvgQRfwBTDdLstQtiyCb0RuX
iSodNLM3HGZ+kp9fEiZytV9ja1Co9dDvyOt7QcWL14fmMxXhUW8TgpekUKnr8+FKQjqs0vL+lYNV
6XQpNk9meUQHr9EAKKozkhpLAq6HzUSrivKCCJTpNv8RD3C/1yoTEe2tLrF7FKHRaNPjooIXY00I
M8hQRvTT6e8EA+23LgQCVftezAFPEfrzmsAfUMT3uEHh2lm+y/ir3U/s4tsVzsmbVnZEPlwNyz5r
O726nTV1RI7OSFw0ojZEI3V8HVGE+3af1aZjEowMaCvABYIUHhSi+sz0RqwboC/ZysPIu6+QSkJY
kWD1d1+Ecz0rtjReqa5C2p8Fr9ShqHRp8sKz1VS6u0L37bSeoOLbqsfPGqzcAx+0W0DiTjntTV6e
ofyXy9WGpMThen7M4WA748v/JaxFPIsZoj8g1Vi0sJx0CmZ9b6iutJ9krP5F3YnTcQFaMfgWAPd1
Uxq7MbgSOKlolcAJ061DsJElz5PY1Okj1McKkx3Y18wA4PB8hH3+rN/Q6ZNSiYiePtRnYsNE30ri
+Xjm7WDPB9rg0KPUb+3mlL2OG1hozZcVNeLm+JLF2jV0tlPnvdZbTl2/XHIT6vtpllBe8PzAv7eF
OA/thi6yHJR+dhwblHM2oW9xkS82hi9qYm1wyTLaKnEESRcTgxKeyaLwW6hKqNMsdxZP8sLbwTNh
dWNt7J5HUiGThuheqyr0PfjR71u2vD2j6MLt0/R6Lu737Nl+40Nh9VF6im+sl16Iun6tEUgR1v5y
yYg0SOl9nFbDjJV+YhQ2mWgoRDQXqCbt/rhPKTgtyaghbRyF4TaT8deacvFqq5ptXQzu1i2m7xz9
1uOrkiz9cBIsbFxGeltvTwn04W/b7W0e4XezycwiN8/TMVwQeinxsc4GU9IKyNxyrOlpXUz1KcGY
yzIybBZyYFbMpd0K5qvsw0vg+SCSLU5PC0PVdxRjclaNuJDD5SvRhnWwuyzfryqD814mTPIdDWOS
5+lWFC3FU/kuH8AvtLR+YwWACzCttLnaZYbsIR0Fw+oEJ5Qzaskf48EuEySa1YvMJ2oFLUm++NOj
y2tuNZzWGLQ0W3ZUxf3A79CBOAiJgwNkJiNpAljBJo5tKwupIsnpof4mXrYu9LjVI7n4nZylk8OJ
0f9lZHvbBCtZe7jfHLM5fAnJq0zEoOxJI1n1EPpSs5ipWPdPEx12Exblhfn+nptMcXbz8kGbX/Fl
ZyZYAXCu83jk6lUhX5S233sTyk6s/LrZiZYGKa4SyMPNXFqaJcLcRxL9MEsqdfK5zminf53GW5KX
fUZ0snlmnMS0K0krGxGFvQMW8KJIFGf+5gje0RYvUXaJi0naFy7jdpCvKzVpJdoFdoYbfaRiS0Dt
CG4WAw4CjHM2784z1AAg8hBetytwc08qPSKSSiI+JO2nLHz9T6bXP2ZZlaC249d/0gxiY2Mmmky/
Y7TpCvCweWmnka8/olUQ4JncKt1QbUNBgdVMjjSrHiuXbPo3lxNDyJ8Ym+Qc65J7L3JuG+Wk7My6
t3+PQM3pbe4AjPqiyBkb5Esh8UkIcmBPXSIvKIQ2gWOq71Zro1Yt9G0nbbnciS2UKsVNlqxii9jS
4ZZCpTMoxs/CiRdWO777ZtS8agpt4t5HXCU3s7MlZfrD+QmBbjt7DbFI+AX+jFl2Cr8i18Rw5S/j
0eblpftgZSnMKRDXoXOWMRnbYa5aLSLbHch5SwFjBvLmKkb1k9lG88rEIiVvNMOTJtvPFI3BZQTj
15ZkSkKLre3rCeNu/5WCEROp2rRQKt3NZbr7XL5SUbkMNEOfZWB/69PNCtZS3uzA0AlF3bwesYgx
OToTTSGFb1+bAvZ870xT0YlOhM/MOJ9sS1M3PQrexnUh0KwdjIjyd/WsLo0BZWQCpVyioyHsGGSh
p6/gkP6OxzNx8dbeEM9/mRXNGR0s/Zci7g7Hf2E0YAA7cuuF9FP1VHlleQwNUzwCSgDqxFK8UKhS
jI3C9K+rCRplEHHCmXrOj9guIKEy8Yq+xfHP3Ahr4YiYtzukXwDGanrpLIS4KT1Z6A0ynVMhABNn
Hmg1RyocF64ng3DqGyFIJn3FgAqczsu/+yDOfSfu9WAP/F3mxRcmVlP6L3zoza2jfHXma+m1S1HL
FGZu/DW3QNJWYsLiRW0GmtlIqezpMrzBkBTwKTLg+Fr1W47VDD1o94NF6jHPjS5N+Z9ULHyJOZn1
D0P3TLWOIHsqRXQhQvWxv/H/iIEzkNgJDF9tzFRd/oY7Jx5Wk0L2c1efSdyC29wUUmmWtgzUiSGB
etK1H/bS2qq/3zpDTaET7b7i68LetycwrEDm2OkIo1oHAWIfg2YzUUyaVggQmoRNJBjSp7eZdNdG
w4DHzQNd3hD2YzkBNAxZjhRXVAzevUBla5zv4AF5Y63F7vB9IaHmpavyqXXQZh9HcNYyWKvYLxvZ
DmNjYxqKPpMV7Ex7ugC5S3jphG4+xn0n/4FD2OXZzLtR4sIsvTLoG2Z49H7BMEckWQbg/PNOcyU5
No91IpK7hU73p2XLdaH56PvwRscS+sXXj0K8npse8dKLHy89cmr3vQMJmrtyJCJdwU3TgAvkfifD
vTN522iAsY66j+0XeW6XMG2iSY+KZIwKnPv00Fpdq5Ulh5GL9VAYsRC/Pb4S0jYwVPKlSo0eIdPe
sKWWrqqpIlZalDXrm7hbtsH1K/9XdxElxhy8DBw1giEV45yOCJzBt0MK5unINjxt/H3TGTnw2JsX
UilpUYBwm3Xvl5K2sx1kO5mSQ566OkcUtjQ6FPzXuEMxOWY9YxZS2XX8qbdklHkqM6TdQHiwvFw1
BpH7IhPENDXLPIkXW2MhkKnwhbDaDOEvQk5lZ8SMZOrww5UI3sFejkjKbGLgXL0n1ygTubBTKqwS
oE/bAWRn1iJ2UnEY9NzNZJ4gj4rjVxri8EfDS6F2xVDvZ4Ejk3M8hF/NGfdt0OLRq4J0POPM3vxH
GSy6wpwKduY0mI4sTjtN8czcIuOSldJerRpXTsfZQwah4bS4YrSP/Iz6ZdoAYOqPsnHZRH5dZGEo
mPNGWUREZT2kTSCQJyY2e4NIVw51vpImSrAqCqCx8NTGJU3ctMMRvd7GyoGpgdqo6eOlP/rT3FHF
+pGBZ7ZA/Fg8FZGu5lNkxkR/yIx7zNttE6QtIWQb08QSqNloYhpgQvuyU+44yqRb9i9BJburCoNm
Izz/TnUD7CVaqJ15WB2JDlBTwnW9CrO6J9JgJI7gQ5mkcKPspVqYZoorDh6yHKDkBkz4AW9lO0WT
Hax5tWCzILsFy2HcTxzDHWVb+SBmtRiZLHvtIKDtwZ1eeiFEvU3HfTf1+SKS6ISxQuvNyXIYmkEx
J2pK4DUbVRpbA0I7IAj5dSgDh1CHAik7+JIrdAfHsQSGuaiZ1ze22BNiXGHGtUEHmCNuICd9llQK
WGzLAH9E26XSkHk5pYByAgIQIdY96tJTXUeWTufIlPR4of3IDUhf9fR1fs7ywsgHwHQfxtw8Htr7
f6YDic5Rk7wkfhZ5VFMFJj+WecSvBXksRyVKulbD+szyaEWQ/yPYNR6TrtKV6QLC0hPxhh9BkvP+
LGsHEsIVSSNy2wtZ94v5msyp64FYsF1yCimF9jB9M+EUfwdG9lISijEDSWwvYwWlHUdgQdq/4YRT
KUxoFQtm6ytedVNIRKYVxljo6Dwo47HJLiV5B0NRjvbjPlds8f/CTHURUNHOqU2zSBR+hQpy9rZZ
I72jlTV/g5NodsoD+X6oRDiRHL08hW2BPmO80YQzcMuVgaMl3oFKKnnwXHGLTbxqfb5yIFrId1uE
Qa2IE31P/Ex4rEoLuWPI3VITr2H3r3eJYpgxN5Ivs9JO34MJrZNTMSh9pyoEuryJzPVXwyZzu10i
jWYvJEZwNaLzZEnoKLZRp7lBo/4KeLZyoDFvIn9S5Hfzw04m6tCw6nyUkpj9PPIp9qhcrYaAygre
E9Z7/7z5KWjJ01C0K1sbXcxsc6MGlVm++oSe9vVFc0+qUu+9LGnvFCPYdx3CqGAP0yd7LUA6Uba9
7GpQS3LbnqEqAHWO6e6Qcrv7fxOuYH5bPITYXBiQr4HChF7j6BiF/IVvFFHl3L2eVcRhF7sfyWtF
cWEE2IkcyppRYKKaEc660zNbGSlJM0Ubqmj40/XDmmktsnE+ntIKVik8RTg8dz8T1GstYG5BCOaN
QBLzN5ogjyaHhdpMNYDZcnyUGS3QuIWgmKFGPggRH6KSjesIqCodx4hVuC4bMJUuOnk9QLsyaX4W
hHF+UXaOYP2E/+ao4vIhE0VurgxqMKPqTOLM9kbUPAuio/rfY3ZzBIV1bi1BjgIhUfOhWYJK5q/J
sTsL1oxKnljrfYqYE3KwKZPmRY7clZ3m2Y2yOua7ni9o2N7RZldmEY+Ci+W/acqWvUx7nb0+O5hP
zvwg7yoLI3jOD+lNfaC0pGPeyiEFkGB2KO/hW8ccvzEDkSoWRMsM8FrFOdMDjb+1GZhgJZCa4n33
0lMAkLb7YA7riG+QOz/3Y/mNVMltJm0UwqA8GxZig7vnR1AHtoRRk6+smK3qBZSsJCH3eRAywpRz
2xukL/3WgP7aTwirsA3gNhDhXpLDZOiYorU5dK9krQRdI9QreyUCZEtOTVQXFdAUCTME7gx1Oe4r
eQGol2GEJgylziWuJA86eMlClEl/EyoTWBgGjs6zr3sW22rBjvOzCEqNtbRltInB0fP5kWLYA/v3
IADPAF75YDN15VYbPzT4tnAThf8s0qbz88HZ24KsazX8vcR2z0+k3TF4qxywqZ7EUNnzxJH80nLz
AeAlvMVLfcurdtAnl8aC1qlZC49ZyETwLpkGgxYzHZzOqLz7vGoiU97ezVJqPF9dZPZmQtoblYtS
r5ynNQ9I5sxK70YyvEUPYqdcGf30JGEKYkQBRwgS1zHiiG9L8FgCHvJ6pnO+8uPaRJi6NFvOFmrh
HZH/ghpsJAOg7bRAcgvapjnUAXia5aOpWRenVyDqemfK4veguyS5k2wXNl4wD7KvE31uMP70fMzu
yLysa150h5dVvpKpWPRmpHDaRqnxuLyuBAzhbzEoXhv8zNTYddF8Jlejhg+7djKaaz67Li5p9Veb
73NqwP7ODqSHSzszlzrxnauaCdSxCfIk4dJNY3yv8+p8IfLdn3MDRAM2HZIcqkn44l7aH1RYThht
LMolkiEaAj3cJH/CbJcRfDD4ZX2JlE/hQeOplRcyAu66q9ZZzTDKJDLmST2bXpA15NdMP25b132e
wzI2fxoJXMfk2c5SFuCtfAHUCEy1jVK4js59Efc2QBvuVIW/mNl5K+uctkCinauGrt6EYF47l4EE
YtnhuIxIMZ0Dkm3lyIWsZzbnUAXRREZll+njbN717Wm38Tu4wQ6lmLMaIHBnof9YIkaXai4dDSQ3
fedaV7GFKw7xeu+S6K8ISIsW8lGR6Ys3EouU5UG7E1P3RwClkjPF73/g9ESlfua13i7Ew6tdELBK
7Rwc8g0kaGSkCZrGGeAYC/EJLHN7OLpUYeZnNvkM3Uq/VFfS6yAmI+skD2C35w4P3KFSjBOo/jI2
czVCSA6xarYScHh4swmnF9dceE2On837VrB8ltVI8qkRTrOnfSuL/ezbc1euePJNhj5Lh0AuUO3w
AiQ3sxKsUq7c3jiae/sNdwUjN7l69klt8BQmWgAKZdQXR8+5dhPpTbTErLLA9WRs1k1Fq674EFna
eCV9Go2T0dBp4NzUzPjBzG3uJkMXv2PXmx+CMZhn5LWPULM6oAnZ9sxXrSqTPvQkC99RUTklrlEt
dDthLAH4+Y2oRLXQkgL+KANGbfZSYt2pD1W7KPB45wwWEGZgHH3zqmTrlCBEeVziY7NC04qapu8m
klPswfb2B7ECAMsBpWl39vG5QxK6Cclxt76Hg/04+ZO11nVpKD9goKNW937ZYpo73/bYibcQQval
w5q/oCoHetT+Zpuh3+olwKGkL1Hv8K2a14tigwz3EICkSK5YW+RzMcGf2B8n8dX8DIb+ClBa4PHg
J6avF1J9ICIEbHLjDRVXOeDlslL7fBc51fKGzLx4jHFZxlybEng1sLFtiFhASgEPNlfpXSWk7vdZ
/ypDMk4OuXel44RVYPv+DNfsFkCYXiSY3IpXIzjvjc+RCaDlgQKBkMk5Cs68Z8zOV5wCEImK9Lc/
YYM5cbefx9GbwH2Tze0AIlM3OMo664DK7Hoc+sy0nZy9aONz0jXUwzQT09Sna7PY6SouueoYSSkj
axieJS/x1JVPIslgO4Xb6/yCAtWwvv9+ATsv+y1IKe+cDl97S6IbgbHjyUX0Les2jZ2+Itc/h7Wv
2IuXf2+RY/hT1RMA4q6irS5RCsBBE1TuSfiHfMpoflyoXbujclnXEyfpJZZTOOvFvoXBBrzNRuK+
qkjP0Rb54mj+SMrpWiqztVSzu0XLfgtYqiHaW5goZPzCd5UVnbB5ke8LM4Xrl42HBsCIqBlwLphk
i8c8EnY/hMFmWiJWh3BvTqUnowu83RfE4LfqI1WT5dnwbClbVfBonuuEWFeg/eRXf/tOHG0ID5NN
4wTPZLESyuFsO5w1WbY7v5cUHAdbQcFjACKZzKo9OqpZjtw/xSXBAH/cvg/O/X62gUPHMK8KEsUx
m2X0ShfILtISOMBqbPA89Yyhkicewz0gwXR+qUplJWfrwJOsKdi2CpmaJUKBiODpB87FRimRMHgx
OnMCARqiUQS+PZRhlldtL5ihZ/nqvKZpmBr6CDdPDICOaxsxr6ER1PfrYj8dGYnroVb7s3j6l6J4
3WtwWpBtPGQ7a4F/xK3mwkxK5szK3/PZwrgoyhp7Hdp3M/W0BqjrOmUtexA45egXiOv7K9xNfJ1d
gLtU+cfM/ZuH1PvJi/ZNAfsTuMU/7OJqWayqcZIRszPOCN213Au81GVb6PAY22AIdI2RLoDpO7F6
dHFTW9u/jajqiOBOhm111Cm2eREKWwNufy7rmH/y372rqEOGNCYhSzyRZOc2hd9epxU3FG6MDCLl
vX5NoxpkLdYxxJv2sTm9BIYKURS5CNBuuV+U37JSr0H3fXGsM65zZpwXiZyI4Lz62EOx+u6bcPpv
LaQ9RdBPzyyoJIWHUadlrTsRt/9JMiVUxE6u3LMVzFB+hUu0XEbUE9wpYb9ArPIDCkZPAePdlDcM
UI5EDOw3QXkX3keewYbKKhXQf0bJDjRvFJmmsiUAlqdQBxB1CxlblkejIrM3QuP5lgg4Ohm8gI6X
0G2Kk041VekcGW+b7oasPDqjtbhxEXx1KoPPA//hC41R5Hxfhhg0qpRim8rtM6CVqfojuwrcWiXl
v+xUvjvGHNHkwYpB3gjy1x704o+Y6u5JDAQzdfptq+i7oEiVH0TwI7qlcQbB/LSUcYZiUOrgP1NO
yJBsTZvx/A7/gxhQxbi7/6xroiNCVGQHcWnTsSMgJ0UqoR76kEwIbFZX4v/qCDQytbfg9aBtP6fP
5BBg4/3e3HxnCtcDb1B7vTvB7COSykk3KtaOfdSQl2G/m+lCxRz3V0X28hWwf2gUlAHETpYJMANT
NL6azkdxdyikgWdzSAJ4XGPdoM3SilW3NHjJbKCaWElNaWRthhVFXt8F0UrioNR06j9PRjnGM7bN
cEtNwPq0ekMySH0jylqxPeFbUSOJMlPO4szKPHWwLFSpwEtPK65NgqVdCtqI7g0c+ECKYJtMDqY5
U/KbDb2C2ku/Em537yrIzJFh1fUhRfEjXiJPKdURTRciDg72nJyyIeL1/nBU6NHNSaNLDoxGMKdr
JXn5IoFCs3vyUa2BTyJwBR2jSwWe8y0BrCziujOHFG/KzRcuMjNcuWFOE1xUc9LdCs2aQSYLtZH6
Jb/DnHP0YiC5pJWuFIj0t5CoIV1+/KEcxt1IoIaVr85uDpVx+p4hEh/diELRpwS8B9R/NHdN4lDW
W/tMpg+7XnMczCWkTblEI2LdRxsFlebw2Z7bjFcemQ3W9HCTekfLb0IE8GspL24vnXK78Ix/4bg2
S9OgpJfKU9RVrWhoTYoGtMOD1rAIoNZoUiDuu548wDpi+tB/4gd1kxtiHdvb/JssEaKG+FKm6V3t
e53eA5YMWl0wVl0zs7OlXgg3NhaItqEbQ+dpYNToXxzo2Wc8Ho2d47kpLuHC9XDlaCxQpyzsUUWg
8zOqZkn7BUTwch94oDDUySrFJ2ICa7QUS0U4Li5k5CVtJR6CzdWAgsj0Oe1037l+VWZPcd20eb58
SgL2wOTm6ZqqUVq7SQO8ioO6JS9zVupVOeD7RRnCQXYBK4R9erifK78QYfZ8X2zdn/oniLkuqeP7
hwcXQTsiMFiTMuFavxOHIdjrAY3kgSjtzQJSKqh3pg7d2RTq9YmNWWoNQaS2WQFu4dtem0dCokUn
xSl3kXFm6ZYomMfCRFaSXlVjanCvZYktYLJxgY3hqMWymqV4kDCVkJBJ/qa11swhYCR8+Av7Jb+K
32Nl5LO1DfXUz2Q/qDXQYHeL1T36KL3jcckWzGQ6NYrDDfEHJwnDTgMSfU3HtSBFj0H7wu7G/7t2
dg2VWm+6u8SYXZsamVJBWRw6K02mCzJf+ALw1g08aVh3Tfbvf/pQTeiaZdPPogiOfB0xb3ALHWEc
TeIHejOnADPjgCvz1X0okhE+AIYPrbNtgFVnpv+jlv9jrIJlQD9YH+jaoRgejKBchxkVMY4396qK
ZIvXR61tKmvuDdLSoy3vkb10fls2HIYtE6tfLkGGQ2/dw1OHHDdPrmQf2d/klSDzbu+epsHkdvwQ
3cxEnHkb6CZq4aNzZYMInOM5e/n4k0e7Bp3GgcoagykPZzLATYDwxl7kPlrfA+AQTuzm2nps5GJg
5hn2sCcJWG9lYwOxxdGnXgkVEVT3vXwuiJgHl9GqFpqGyZXDPmffQw/pP9erRHyLMAkxgHa2ogo9
m5BKLlZvMUgKVzMjj8b/ImZFcyKk8TZ4asX0VIvk7eyQWlYrznqND14hgVlEtkJL33YChRuKliX5
buKQejw/fpprzca5rbqWyA8Uky/TJQ7H0Gip2Apk4CMGPey01pCS9+7KXc4q2uehLvyoRb1TmMpx
IDbj8ljfyL52z1OXWYQ0Ib/zWImt46yRxsxAYAiF2kxDgoKj4ZT+2qhZBA8AcbENxFrnE+KqQyuN
Ajw4hipIF26AbqDmW2ayy4cgbcQWlEiMZOhyHu3JfUiumSbdcoE2ykv2cAODzaQjqXOt6ju0nKoT
xCJ+iHvGehrAVKAeDDGKSPfNBBe2zH3sONBOc3jhnu/BIAM5QRY0ri84V6brv+voqspeuu+TDlow
GrVQrQlBNk67U11osT1+GQwPsWqkqye7zHBkvRyguSJvc2n/FpbU2N51Pn2UMr0cw713Tffyn1Wv
MyGoCJi1zQC7V9azQlVeZVFuP4/JR4JQV7A0jkTjt6BDimrFAgjCPmUA7GJZ8EldDHN1ylXOcHdd
AYmX4Wa3fengx7qzWXTqrJxNqBSzuWkZdGCZ3ke9RSqU6lA7loBDeRuyHzevOd/WGftCUowdlINW
RY+IElGK/aqtA2u2dFM83pu4fekPolxfkqv/SqbsyIK5Qgd3NaJy7Ub8ZKzCqYDM3bMZk+cJfG+W
S0jojN/lcvZ5u4HAc8skSF4ZNu6TpD4Qu3UOvLPsnRDn3FJFDs7cvM1VDFczVAeiFKBKC1Bp1FTR
7cmymWpueqCpmX3/19Qtk1eTWuIjGnYIZW/27NbHt6F+3jou27pND48j7LbLTNGgPRsyI9ETTZQX
VJHa76VvWuEGb8hlRIMikHBfDNcEQEwXNccb1YXmm12C7x3mCDEvElqvihmDqiw3fbg7AVQtLIoB
+swFtxhACrDqWjP0LKaQvNCtFvIaAJeSYnPia1LJQ+F7R1guqDqJ5eb7hdx9mLfRyC54qrWrj4HT
7uOsTrWEt5NgO0iUk1bwfyvtRq+FiNQ2QN8k1J7WpJT3pBk/LnFDEkKkOTDJRULfYTBUf7Ss9nyh
7uM/QzOWppGJG9PWhPjthJX75Am30JqspcSKeXYPhkXPiErm/kyB6j8PNHze+gbKtPCOrp+6+ztf
JvVRK+6VDeUWYd7ZiMHt/4EQcYdrZsjbkhPRKr4A+OrgzqIRNyQhshB4wlpyOwJC/mt6onkc0yWi
Z00mXCpP1c64BDrhBf549L0WvodL6nV8C7YSPoXSxl3tEvGZKB3lljhi7BUGSm86fgoMJ3A9vKaa
RlQZVXvYWBX/6BH70PWfX9wwMAvxQPViR5tAjd2yFPyNY5j2DHjo9U1UdcryCzExEBIqIkh097kh
rmgu5K5VUArc+ve3BC6wDBVjUcwNPQUEYV6VXXWv1Wb36CfqQ/JrClysMvr/OnbhGPcmqCtwpIp1
YyQSnQXQUIqn7tf7YtRj/Hh9mWAzaOLeduSvrA903N3AgMoUDQZXWACLf9fHmnbT0QMPMWWqGBRV
bIBKqwkMfNdOPKtY2d3QinDYtYcw+QEB9WJidCE0zjQ9GjrGhNoCzWSD3agZjAylFhrP/lCqluGZ
iO8J2IkmlPt+exYglHxMvTKBTg9WFBHGvQAj9ARGKno+3JtcpOEJ6uGGTnHqfzlBaE5Qt7aesyTm
mk/qovvcbOPdxLaEif7xJH1lm+KrWcMqex9wEhYsYwBUmNbwZzZxo/W/7RuthH/0ZmN+sWo11k6j
tAdR3P/BXvalquKSegd8xVBx7hvw9b2CNVEA/niDe1hLVS5EEWwH2UHfPLpJVXdIGG5Iuqgyzadx
dMxreh4OBi70JQ5sOGSaZa3KgfOTE2WBVVCSzWNCmzwNhJc1El+9e3wR3ziyHFERY5VdJmlnIOlW
38LcclElndWKNPFiqrcCczcybwQXenxiul5M8xC6aB+HDMXHJ+zl6aeDsWHjXtG2wusAWx3iKI+V
8P0QIuoQ8SuQv4ZuA3d/EbfsEy1CFYiLiqBjqN5CQFCQz64gfQ1RtxgKDR/cvU3/L+2/+Knv1raO
DGH6e0dWBFknFoDE3adwGsK1bFOiYC+05LcH+PD3HbWQ5ou5iqRCG95G+B66teGx/VHCJgdcRGJU
WrwHWGvSwQfHPyyMsTZx7cPwI3Vp6m79uVKiOwGtQlyNL0/+pO9xaWOjEYjwn12CF0wYXN60OM5/
lz0UEAqSbPo1Q4bhegnuY0/y+zEfOjSn0Ejcz4FJXGcdAQAlcMubqz3wipYuvqrIpA91kmAS+Axa
f1KTqb0HFHRiE+IHOTQkIRFzpTjL5C8DHThHQCVdGjMDaOQM33Q6IDbYBbHMxyKu24mcCzi5FIo1
a3olMQQzEM7M0U8ThWAqteERKr/lO62+5usOJpFtT7ApVM0tYMgwtkkKFDN2d4hv97EeafjKJux/
IF/lM9ypg6PTmcibNteNJi5THFdHdmA1V1XecrfQx50RbjlqPRu08ZiWQzCUR7AumLAEoaiV1w9w
xZPeqPgxIjO1KEz5tlvvGE2sP11L03ytB/vlD23RZ3R/5wakzs1fOgJdctqd+gmLE2NV01eI8h8D
TuDBDGzl/gW8ENOQS4Ls1rqtV7wcmm/JGToNuKsWjHa5UJXs0n/qzhn/wCN/+JntZuu8mZ9LeCX7
Q/GbNSbDDYx+Xv6Md0TcpiOHHkPdW9d7rnkhOHyTo9DDLSC0AmadHJCVMq4dahF2AOPLdaRl9Bn2
LIAEF1IHH1M6LqJ83ayIBpLOtwX/CxMgJQgLwAeWeZ6bZOlT4wQ4CU36D8T+eiKOObVCGm/mj1MF
XvMSAnK6Ly9mRgAyjU8/bTaM1lvM8ycT/IDg0xvSAQqVzlBosQq2f6Z/TXwKPPNBEBhnjARSM9Vb
cSrqASRFKRi+fBwHpmyYrf4fOwCv1L8NKuKccSOFbJKbGBSGMt3LQ8Ljpuv0aplfDMQj2ZSAtOvu
lFXz2nUjVunE6M3q99XpmZmEea5A43jnZR5Y2XOt/9xAcUwZAsIa/pd1proDCguUcCjWpdeTSRC3
EGS1gdC8Ze4GQybz9c8pjfnMNr8KOCwcDu6ulbsJE6Mrppq762HPJcR3daTlhnf+PKgfrJ0qCXNH
jv557QkcIsiShFLMnOLXDTueSemYLQfT2IJ6Qkm9atFk0n+3Keq2XB7E9GZcmjQ7HD9j0Yd2OqtG
3DZfTQwzd6c2j7M263b8Nk1GbRYtBmxqhGQfHhD1/8wqhyG/m09PhtY2TptIJSaudRdrHPge0iwx
TTyM1AYxZd6kStFR0wRGqyiYQ5rixbIopjAR+PzjQcSiE5cnoocDQlYcWcYs9XVKj+OaNwwNoajQ
vLVm772XFnxrEBAWeXjSjjyGZivvWCANeOWrv60x/XY1NbIpw3PPmga6mM/dunsFQt6ROS9G2Tk1
5ISpeboH/+2vwTQbxh57vwBUuwz2YcqgoPunUBlV3pCgG4V59WJJFdFFI97WISsDO10Rx03Rp2Yd
53GNRlyyygijwFpjcOWI5Jji0sauqYXoAW57ZmXSeITN9ROvflM8BtHGhXWPX/48GeXgU+Hlz+PG
cwSBycNHncxHo0myBKwfJehtlkEktY5n5SpK4pLjrcKL0rMXFqjJGWrWtnzfEDtL5TQWauDbZqBQ
NLWyeagcMmVroAEMG9YLnbPAXDd7EbXzQZygya6FqjzqYBg1e4MsF5MSdh3svzLo9SCpL+aXkFru
32Zejx/okiXzPtL261ayRtec0BCun8imD0yn2h3AH22vxfxTPAQaiIr1CYiDKW7jll5YNXN8DrSw
OzU5R3NT/LsgfhrByr5/cDte+W/70CyYmCJ8/gj/clsYqQhzpO3MOUVKLE+j/TeOyOFAXV8jK02h
D0usHXub1JTsRkgMB3oo4/I3oiN5jV1ywU1DYkZ7NA3wEokLv1z3OQUGHOySsDbLBzEpAe9vinxJ
/EJwulzd3GEtq2svpp/NNCY6T9UmOKgAQVCHq6Qidxflt2F+XMnLHt+iAOOBsr4rNHfz+vW2wlY7
jtYaGNCWdHXcrOLxOKCrHhSzvUk+l0ETqQ0dhDIETQ/zNqdZ42T63CJpeMo5nMC9tztpX5AMqCPs
+Rb9SEkib+foMzsqCdYx2PEc+lcEc3J/cChi8HAJ3ZsZTDJGTW6kT2+C50bg/yp9zlLZKN2H4LI+
m8cBMeTHZuln6hYkFmrNaQfsaoW8Xa7bjVCM9sqOb44lD7cGxlBrBpGUuJlMQRxlFa2GomKnG6hI
j/i4An8U1T0ea2lKCS24562s+yyp54ejkoZC039nU4LuS1zDANQo/q+rwUx/hK+YWkFbvfDlNCAS
z0LyWsCu7fnZPZOazahECPVMMNa/abD2StT7Rz5vqetFIphjQ/C+L9hY0nCXD5me5u767HHg9Qv7
L0s6VzxE8u6SEk4HADB20SsAXHw74ke1xJ5rt6jS8uLRhSVN2tcmTytm1wt8+oKlqt8P2vyUpY61
amOAydc65PuPtqf3DVN/hpnAvGC0Q04GmggtgFWtudXe3KZyrRruLfCAVO+BXwjY6MXXqD7MXexx
q4HYFJYWQ4eWu52PYOd6PDIPoXJ5WJDHNXALYvNPel+QaeRD5U8zuPM0ceVZU7JN+VCReBDTxqQr
476/u6JnfGaGbhV9A9aydtpkOeGHShS2+3T+u+0wGxNFQSAnT+tP/zim8fO7qLayvWCkqd5fPd7h
U96hkuGbZ4JKI6f9jKYXHCaZiEPto6v8WEfZsFh6aLHk1Saw+3eksG3bxQ8Bb0orjnuzsNWzCxA7
jOnUBN0PNUMOrjDpmDmyz/WHaA7JGCu9j4yv1e4X8cssMKZO96Y3g3uEl8Nj0MSH8R2zPTWeqKsO
b4jLP7Ik7wB9yJM0Xcuz+6pW/U1jQFVjYjG9A08BHc5PldTT6nC6TSA538mZfCjJOIVtPQLaBTbn
XANKRUCGbYOV35UutOrlOGOBzqi41lFUaNQ4KzTuyX15YrUpBXsLqwgU5KkkGmyGvCQFTiIgnrBv
JZf1Un9Kj77uTK+t7sSmlVq9mvsOee85rPuupCNQyv7kiLZILXjtbbs7US871q85j07pi4JWt+az
CVfetWJ7JYsJIb8PYdNJqkdmYJLHBWhX/3p5S40K09CoNFl0eMZE2vMPdRshUMqgJKWJNYxH5J0R
H/cGbPS82bpobZ47OJojONYcHLC4IKGhAO4PjA6k/N/3B2KKDt8qGSZtXsi38AeTiuMpEqvgjUDq
zJqYbp3WyEA7cHBeYUCRSqaTmODp2wy4A4XrvZ5sFknAXWfWuEAwQ4Dn/gHrLL681ZVoIM2VRkk8
E96W1Bt3eeiQDLfeyCT6MOnMG5zYuFd8D9Lx3XvQzNpMKxrxkV+yAzSLz0Od1v3et0TzzfUDNHHG
ddlFwlxbMU/6B3kYI+OOmn10oapaBDvy0J2Ip/2oqT1J2V7klphwE4btPrqVQMSDNqKVFkWkCe5c
2HJ0L9lIWRU3s4cke3MSU23St4PJK3xfP2WBPleq7inwcDqnW3dewkh2Lj6HqtFT7KL9WsJwd4Wx
Uhl0dqtdwoGFt+wRuAIRmUhqRdY9tr//PYt9LJRpeGsMVgUnEaSZ5JxVw1fDepCbF58M1Li6inib
BdpjlTd8HjdTW18zGY5yzz7rYTDOhJhp+o7K/uD4UXKb/bhRd4Mq34mRJo5PKVbQLfMT8xjgkNNd
oRk4Po5mZAwT0O7D5XgVcUAym0O8kwGFuSlEq04i5zw1ADsHNkkGK/Kw3BjOQGsG0sWteWzpxvdF
X8sSseeXontToSq5yCEsjH8c3LHGkfvZfPBL8muLFZHVB1wjurPHV9L6bduQGTMkkR4ZDXPLcCiY
hI5fdEbl76HxCG45ivXwlEIFhy4P2kpXtGiCK6YbbJCbmsFZqIZVkS5RqO/WWU+IKuGLX/8GCSrH
NIScX4KlNMfI8y3EAFDkfyZvRhb3agt67mKB2kPN9E1Yy7pnb3973HFHeTqeQFqshSehLK4XZllL
1lWKbeQCV511+XRJVkJI+vy/24L5qw5ZEGV37pK17lfueO4wsGwj42U2e3HJwCIk0Wt71dPcmJlR
rUIwqHn2DIXEQQPzXuhnyxKllcKajJTfY3ugvY07d0t/IG8Sp6/b4M8j86d7n5RScZcks7YEopz6
vvvYx8Hdlars1KbhX1YvxK/+MmfAlfFpUrlM6KpGjeAUxNC4oRpg/oK1azvItz/yVhVumHSEGu6t
/khXaI+gi3UVhPWOO9iYvOIa9zjBgKaXcYE1KF0aTuVagTxWH8aQ4ysQzyb98pv6X7IcNiiJx8/E
rsttqGkqCqPG4B4Z5PTASk+/Oh8DWzyvoq6ysfvQWddtBbuTvZ7M7E9EQlpguaXG+wQU7zrRoYbr
ZIcmYyeufFkFq0hf/uT+c4rOF45PtokRy/+3FiU8TnqoEuWeLXO6cy3bbzLcC1aFqtprmCjX9upu
pdzVFBaQSoCb6wzTzc2x8KhtVpUGJtP7XxShBHt35Ee1cV9IODIxMK900ScfUa/he0ZajyJYKZS9
HfsrjduROf4XtRJ1AJVOa3Udv5TanZvQV8kxI0OuHGXWn4Sp8xKev3qysBi0GBhky/VeoV1jo03e
Nw8ViqG2uSTasJNgB6ye96w2MpyyjXodj129OzdKeX2piS44XviVyeVT+OSa5bO7GcqjZaX7p4aH
vI2V8p3yb9a4pP1Z4EH3slpcM29H/bsu2oKcsnUvB90H1ZjkXh2ggu2MMC9s6bswsaLdj/zNj6UP
gSTA+0cNWOEBvKiaPvPWs/bOS6MeHOL4M+IrfQbYd6QO7D9rQBg3o+yTtd0ue/WJdFw94kY5nH3t
HV2ru2oZzJ0UiJ5zcqiZNB6sYv4Hz33r72SMCIVA/2FBdCKNv2rRxOYoYIg4qKu4CjBd9X2fC/4m
1RElRkGgvdp8th0VD4LxO4m2bJwdkUM9iuEbU6+PDmRQvOgvbcY9tgj3MnFZRoBrebNMq/3iaIMy
e71IFLdko0RtzASZ7pA0NOPNEC14Z92c8NFV8mlMQJzmJMclaQZhUYGGjbqBuDyoV4yg/XC9sliu
N7Yrxm6qrJQPZ4+Wmq5CT7nwn6t4c9UDQxJ3xCwau/oSMXLdioJl2yKk4sSPcfkj44nCceL9y+/e
BjskUNfAdOi3sFQjNSjgS+jYBF/Ne+ThdXGZJ6z5T5S8md8lPWExQbYQ4wAVuKthXsqxwi0+PBUN
3B/JMFAiX11rZJG4dOBmzSaQuD+9z0wd6e9W9opb9eLrWIReemrlStnRwCYQ7bqitmq6p/WPawkG
xU4iguaEOoXo+sh5DlC2TxpD/uFMceJrapGsDTxyPhoPQ09U4vHMaR1FX+3i2BugfmMOw6JAmCxW
C2MQ6moez4XaosIocCf7DuwKsYcN56MzQtq/Aa+bq32Mn16dsDC3RA7JZ5LvUs3Q/TF9sZL5gdb5
VNaCwpamZzreOVQUwAyQNucwMLFZ3MltqqA+0r6vaHN9rLXUMCeb7jNzaN0iVXW9GWpHu1G7Z43h
SSy1a/CDCuLFLpk8tDNjG4gDRIC/ak4kQD2h67QnR2Tj979435xv/WFHTU0gu2KeTq3sbRUdi4oQ
nRhxInivlD0Dsfn+dtd210YEpVpqUxMVTPOhoOIXn7/SRWmg+sXypjH1Sb+tqCee5X4fUlgfbY8q
nenUdgr3fdaHryLlLYitFJVSE1+GOFrFnNEJ6kJNVVYZ5W+toi5BiuXQPV5S9GUrVS7eodYn+8Yq
torIGmn3peNLOlN4nKPrCtoqJ2VyyizDmw9biwWyWqgZ69TknfswfnjoE4Huds3zwlLIJI7K3zN7
zE/jh7OH/xqylZ6kQP7ircAX/6kW/TJqi84Geivn91jVq+1tCY5+zB65X/ftWmdxAF6zZbLUax0i
ocsl7zJEG5/1VLxi0HzCEv4bC3NXSxkfRhWcKEoBpS20fWm4KjI3CQ7ziptdyGhvjohX6+XGhgLk
bGERl/o3NF++pAf1dCliUHSNbjTw8fBaTZQRFD3xottPwdRxsrJoFo9mfg20Hh2zPLPHdh7cP7tV
7jyj1X9JvdPD+bVudCZBWxP50f+sbwiKS2UCo9HPKLwzaEBfL+U19tupVR6dor3XmcmoJJtil9bS
SDs8O5yZVyyOlf1D5+DNp0kpKxzmxFPfeRkPh+dEd7uFcxcUV4ErtVyTgfw5Ll1tJcWrq/eQ5N7S
UG87RAEkA37TV13ysoLijGfnTDtVHAmIbck4sgEntivJdcblDKAfx71fluqkk0RWBX5/Kvc2BPmW
voVG+a91BdRMrs9AnWpDlC2dV/dT6SvMw8FuZUmPL/ZuYiCuSzJW6V2+Y32JisdmAE3AmMaOnOlY
Tn9vyPXOcJAg/yskEUvUM2V74k3NtdaSmEd4lf/Onrj9Ybv6qyPpD5+2UXmcXNw5FR4lz9FO/lJ3
FJiVYUK4XObNLmDYhFJGHTWGbam9qFr4YV/aL906W2+rFS3u3s7IxHxKAZrIcI+3ch3FJih1P199
1oAPa3e+NcRphMC0U6E3RDQi6uIJjSI3QHrY6u0sfDSv+SbeSQf4nZoIBGSW+A0gUGS8BW0hDKhb
VklpVahSYOv7O8oRk5sPbqo906foUVYLt4q52sR2a2zjuIDo4YmiMD+P+0lIQH9oT7eqMEaGzOAE
Jmj5TRyFEpjAGNfnhsg+cgt6Jb6OF6sD+PWRfRJqHRpgUxW8pSPjYdaz2fCtvk/C7m1sAbtVsJ+q
4Z934RakjVuENbnxkQktWB4p2/ka5E/Hw/c1NzJOQFFdNjFXDCPXgNVsk3k97nCJcOzb53Ntu3mZ
TwGu3u/S/mTgfc3YuBQa43cji64LYGoSXHtIrZDppsW3TsAmHuTCzjKQyhXK61m+svM26da6S4Kw
jRjfQoASGQHl60VqoU4+EA4449G8tk19FLEAfv7qH+pn+tEDFHcMLfaglIKfd4IO90Ehs2IXuyWw
LII5wuLlZJkOY3pU2sLgr98ySle04epr+Z5UIMKMGqH6RiSN5UJci6pnXAqGfx2hIkUl7x8NtGQr
CVfWqaK5V+0g4p3kjdAz8s7Ah4OfGlEFzNpjzt+739Mr7cn2qY66rNfLCCbgNBc6Ajj5Go8x7M4+
X4hpBR5GIcZrLQsgcRsKSdP9qunwmZRWwP59mBlOM07clnXNKv0jvyJSfnZCNoAQNs/6irvTBkSe
IUwmg0o8clEXadmH/2W65S1mSREPl6X14iiE2FctvTD1KCuSYwdbFSWz7OtJXiq+8/leip4wXKHV
xkd3CFRceov5lLjCAZOrx8X+Ze9CSXh0Zf87pisRY06nBORBZJbDikBSG2wYhXzBNmo8LN3AdcyK
qAQXniUdf5BunvZsGpyjDTyJ+vCTiakF1RSdFiWOhquQY/GS54VunhRqPJUJ/TLM41/QjUvinUHl
y2BAxaZVL75PHlWT8cXA6xDXxa6JcM6/pmoWLRqmwKXLCyUg2Xhu2eWaV5Gs9zmyAW58PMq+Wpxn
2PQlR4c8GRza39QRjobMWh1a6gjqK0OYVoUSbLJKwa0GPD7J1IFOxYkh7XW1ETjTC8zbp3aiTFWq
0KjuwwLkSAgALl3fLQ3PylKGd3uZBzIaLZjUZ2LMnmFeUPWoa8qF/64ECuj8DjLL163e4AyMSPoa
r2dfztL+qi97WZy+c+/TZsnmdGVTr+x/mvJuU/Sm2awWhhcGPvUY0NN3UaGdjn/+5jZANtc4QVse
co/LgjV4HH/d0VyI1cKncxeyHqP6zyK4OSt4ofApQ3THVBfmPP8D/tuBY2nnQJKmci+xKuhUCAZN
uBp+BoYwGvWs6OHBj/eBdpq6NSaJv2PPO5mLFJ9tSgbV6YBQ+eySaxd+eL/I3s4827gxRqUsnNks
KD0ZCLkomvrkYPJoCZEw00uhUC+skpvwLDikpZP6+PshCWQYNODbEwto+mxCHLM3Dv2TqSHgD9o1
rPbXaw3Y1TH+mZhBXzITuvIaV3NK3TutpELL7VS0XFTGQQWaf3wHYpeuhbPAAnkeDP1EnJF1XTbd
Abq6HnOc4nEMTNuULTdPrPMSYKBpB3Jm8L+C0YGIABaEvtGY3ePCF97C3fU/fsGYbWojWuU/iZQh
X1xtSZMd3ZZ1h9FD3zI/VgYP31oEOvLn8afEP7iSdBpZQnkxKLm4sAZYdYaPGeo3HFl3d66oZrzC
PEdvW+WmtURtxYT/xfQ94utU5LCKh0id+ciWdHZIOJ0qI5HBYyx0Ze4L/AEtppsU6NAeeNcHq/CA
vqyilLN8lGPuPJ8tbHNcauE0++DRmhdpVAG7aMxBOoExZ1YbAF9pJB2AERDtsInIFvBsURHvhl1U
YsLYBfzq+EH9DZEzGkJQxSSS76vbP0rMLCMgnhV1pWBoFokZz+B1BY3Y8dSoNFKQW6hvAzTwBedi
cNZ8NJs63+if1lGEUOasSQnE7wIc2fmcQhJBddZM8LW0WjD98qFJGCL/rZE0ybLfRdMVvJ70Irhs
9THcuGHvq8Xq7tbXJOrkqgNskJooicfhMWNCox3XEPlrEDGwED3iKsELhKacRnROfxQs077Y89Zh
kQnTTlwWVQ6E0/+ilt+5ivBHk1H1d70DB387vlEahDfy/HYc3/SKrKgdeEjjKXEH58oBs+TYdCLE
HFDozhcBDlHwjjg5JdFTCsKmipm6ONIZUSUW/UWgQlQsNzjnHnIqxSsR3OepPhq3RFPZWdEcS1pQ
l2AHTvKPHkvTedDSSFLKSVuF0o/b/k1sTIVLvfF8ccPOGhqPdgZliZYGMK+yw6QCH6AmaqlR4ibZ
+DbUrqbvoWpuDKWYz0hUlg3J0Empc9EA28oIh6kwczqVGB7wKuI1M/PHDSXLvlSt1IlHPD3hlk7T
//MdZedVEV/QM2XnzNExQU+mM5Q30Hz08pcTAqM9PjoVHj8i6uCr6a0YDu357XwcaevrKonldrEt
Lgg1dn5pkkRTQUvCGqEYqpuwvCHkzWY3/q2jelvu+vSBpQvl1j9Cgb/qyzxSS85G61kHeB3s49nX
KJj109lN1zQwHlfitAsmeFq76zTW/vwvNdWlAPFdZqk9xRGnKM1vzrww4qONJoU4RNQzdZh5LYlR
2yH5zoipcFM1VJite5zfCHEPqaC8d0Orbvdbs3BIfxlBEPQu0NjQzBqp0jqxfMVeXds3t+WalO62
gef6CzQht2yNfUTHbhiBHA8llDGXAF1+hIJASQmkksyiXJ5Z56LHtaGOrRKY8istcWRk8EsmnRnf
cVuD65I8R7IiadTQnELJEGfASjub+AKdxTTmwClMrylwn59iBZC2nTRz9mWbYACFqpkRecJb9fcN
a7eXbiQNsaQ5GuACVnueJTKSplRuZyc9tcpOV9MWBD/PCRaUBv18yTi9v8DBQwQQ8KpPXf3NOn5p
Nkho3rQcl2fnMw8tReHKMxCws2ngQUUzxkF9qBfynjENyHD9pdlI9FK3C6TeT4oziiKeNBWtTsxp
rrB+DX+2E4o5oxgObzm1f1ZpcNxVIk1ol9cL4NFl9EzaA4llKfTa0SXVShhECICWLM6SUZQLWylm
W6BXJwqtzNnA/n3ol8SNzgkvQf07yE3TxYCzumpiJXerHQrafoN5RUTSx6LtzsrRLNiwC8nq9sGp
Eydq4iNiEF9SBXIrzRaoPd7sOz+5zxc9tjyGB9THHW0XJhrHmz//zUctXYcoUt9EuSSAerLbASR6
oQ856bp6XQhhUbHAXI+pwbVxVyvTfDr5a6xhIv2fBcIZVzNceQFsN9XZnP27lXWqm3+DhOhUCKOt
aKAY35bcwV2Z/6fdtjc8o8jrg1ri00f1uliQhTDRGxM5bZ2VRPPmvbxsNdXFDcKqENxRZRkhSUfV
jeoNx3WTnInatD24oFC0RyWbXgbxoayjcjLCLPEMgd5XCHu8i3duwejXQcASVwuc6X4tRqL6eJMs
JJZU7iakjIdTUKAmfT/LtnERGrC8eVchEBz4K0lRhKq3xbsGQuNnfax0Mf6aBWcctyj0+JKPs6GV
tZ1wrUoGtgrH0jGsQc/yQNszjfJBksDKl2nY2kg9KuprdyM1GIrRO5PF3iVUmt5Q/9kJnh1io23K
WHaqVelvADrjtVhkPNNLO3yUU1xjfbmxZ4xaomtghOfz0HZfXs+2Tdto1dFwivX99Dk5qNbJZMtV
MoicOoXgy7tkKALd76yo0cwykmcom/oXhH3Uh4R3iBBM8Ux5Gd6Wqsl0KYrQ7T+H3RLRHJ6RwidE
9Byczk8kU1b8+aDKD/BH2kLJN/qM6Mm2lVPqhXvr+ydpq55iQpwq+MM05ISNpl3RoxSY0PYN/cm3
NytAjTq13vl0BqCV3JfGi3wQG6YyQgBUeWlgj+mVqQocMHgom9FUndYsLfQVu/IAcgHHqm3amYaY
iixVhprOlOW18Q4uRUX3n+7KEW2VozFbW86zHilDUTS78aeuEo3Xf5869fnWxtmbCnDf0hbr+tKg
i/3liE6NZGc1H6SJ7aeUxfMcNr2Q4hMALT/YvB7uxi8Ta/S7YS9wfAU55I3IRfe5JxoGxYRvwBAL
HyYJE3D6Dy/FPaeVzj2gRbAKx1q+m8J6QgLUvviONAw7XAfxUp/f2uhLyu3xCTGo4uibsDgykqj0
+3p8jMORIEDqq3wQPIBbUy9RLLhOA2PYMcAr5sQdF5YcaPWpy7+RIUj1zYYiCphDNCQZ6QpyfYWe
bokbFQ7qVdwECyynvma3DDxxSVllt1rqBZyAj2okFAD/uGKFEupH4jIKooXLHWgYZFNNAN9uW4QJ
vf8BvBx4lYaBkkirwYfILvQ2BknLzSUK/ZTe/JXtJYIs2LpyJ5A+MPqFYPjUqYLuD45No+uMbGDd
CSU8KhQIG4KrheNmyJdnuk6bYgme6kbBRidRRHlcLo7sYzBg1nctSpjPC182AKBFZj943JERK7PD
nqZEwEPOaNqR0e7SY8vmXK0apBkhjgNpKouynFBXyPEJsBhh1qT/DXlP4JJ3WX8QRkDLnb/C1NAL
q9jcGCKB8574bEfrCJFu5ksMpSwEw5pVhfFlE/anItLEt99Uww7viU45sS+vCAOVWCzW48pidJxp
z3F1TwQrNXrjOddRXBaOdwMoTJxDa9y5lJs/bu+jGHCGumDUOT/ilJ3yz9R5+HKE9PF2kq4+kgQa
jgkL9JGeeQuXIGFL7H4TDurreYQHkezpl5jMN55YDQpvUTTg2gbErzQ/IjrqPRi2c0muN3yXpJe5
ZfRHaXQoOWKIjmStaqUl+BjzcY3CnZ3BXSe34b8kntP4lkfBUiX9cNpFks3lNXrWvWaQz+5j67NK
a3SpoNv8iFKV4F+9oHQr/bpKFrwLFG3Vt4PTTT2eQD0cXyVPW04y1XOZ59HYhMsG1bDysv72cKXU
ErAt36OSRcOFZZSqrod4EvC4kBV9pcck05KA1MZ9jIhM6Q7ozrhf5nPHEaJHl8XPlgnb8qdcw0KM
4zmorX4K2eVAUORd52qh+cALTgKiKkDZFITNI2T7FsMUJtYDq9YRX7Ifcx2vVEgKS3dO4Qf76KSh
mVIu13wge/DZJ3bxPLRTmtUEkAZSDSgVzuAU4qXLIX6Zbl5pUthmCkvBCTySgMD0OgTSaIdI7Lrp
9HdefBjgMH92iEeWjC3wHbfBmptZddeeZZSbAz8CJt+C0ER6R0mnSSkgboaajCqWM/Ezeo0dGqM8
c39ZpBwQCAabtlhq7AvBpQsm54+NMxMe1QAKhAYV+yCVNJM/vi5vreemulK8Yubtf3ye0oTNehD0
0RL+SNpc0YLgBIyvSVFnHT4Ix2P/e6puKglC2NsyXwJEn0o0YQlgP+GzpLhEss0RCHez5HLC6J1P
NQGkLAmsx1cEXZVZ9/aCZbK/mgE8rbEDJV6C3Tm4QdNpV6cAXTIzuh+C3fFtLRdM62ubgOejSKlo
4IqacwcjDo+YVxOezQzr3Nj2QXBYhlyjWeHM9M5aoeRfHioeRXKE9NtngmeCIw2/wMqMfjqKmoeJ
Q9s9NfxHgFG2EmMVG4p1Z9YPzum7HFW6vdQawjVHQZmVfgGkj84cpb9b5wDwpt2CbmAfyph7LnzI
LzwvZOKtPoG90oWHvdnCwzq6CKBN3kGTKLc8cK3GlHwluuCLMBq0MPJoZeowMkYsV11LHL2fNDzL
BWbVwQvV8BL8JjPL9njlCVd7m1tVH5eYp+ZJFxZgXvwdSWF/BVZ4lz8DD/6Qut9QPy/RUduQri0r
1twGtA5FJcMTJyq+spQxxdASF+UEOYE67ubFyW8YJwiZX6qxe22egT9S+/95Jf4syu7soFBfOxb+
WTocuCl8gET1S3ywOkwsqK40MmTKY14CZsV7bwrOecgx7vpTHXJz8wJVe4KyRU1EIYZmTEsUh1Lq
KXCUR/1hgyhLAqpCkIbhMbTee6ZEMt0iYI7mj53IHDmiUxADBOMsjRy65vc69bJiBCvdG3UCTA/Y
1VMtWR+2dNLkSWJ3OdvuQJJuQTqcK4Iu9512rC90nG1N0dxuIkk6VKBzF6+ubkTRwWQFgtcrvmMP
m3EaMWaLy6uIs0nsJ6GMcdvMplJuhc2X7eih2f6pLFMFlxZNRptBhjxIU5FF6ZBHJRFWLvD0hGiP
Wrx2Hy26EgTAIiHM6hSJqnV095riDz8Z1YY021JCm1Vbc1QOW4ONYvE4FPVXjKEaP7kVhdwTUgi/
BcI0cH9LHW1IFJPRKI/VEtO9TmnDoMTacLEfDCsFmdoXCeFo8QVEqkiaO3Mh7fFh6yG36GJi/+rz
PX9n2b+bhiOaV7aQ6wZ1Tb7+T7933OjVIXfHZMPWKabVi5oaXLw/1Q98umqss6BbMiIZPzQfM0Qb
KOTCidT5PK50IdzockmPiLDVkBLy1cnLp4S+P+Vn3jY8oPO+NdPVhnfD9JHdk0M40ow5hecsrJ8A
BAPuUrvSt7VY48eci0kKfYRH1UFEGV50nUoPMR+sHq3sTC8xqoMuNAW+8sRPKjgANIB5kZJd/jRj
x+q7R3kvTuJorECVyMMhg8FZBZ9QkYPwXsnZg8rNb0AgTQ4/YrdDn1RbhHpwef0Oew5stS60g4MY
Bf41Jhx6QqR5t0p+CCaFC0xX8cdWz61TT6e0k+E7QU+O/ES3bFAacytSE/xMMRn44a5O6hVfKaZR
CbMjL7hbum9y3YMjF23BEmo6klyF7oFkSfqTfe93z18e3v2g6oqbiVV4Aq4Q1MAs+i4pTpgxSern
GuHgb09laT6NxOfLSyZL+xbyMsQwHy9sPPekmtUtuCVR3VK7FopIxR7uLAbodEcAqp4hiCyAhit5
RwR1TV8CyI7InVBTyt6XhvAHFN6BVBslbUzu3SiPBI7brKfizPRN7fDpxZZO49NOMZQ1SDwIqb3v
0pMd8d3CmEA4C0MFfcvboQ1rFypeZM+1E5olwGPTvDBZ6NdEJV4ScX0+anBYOXGsHUTID1rsCOLd
W2DOFRtH596h9EMfHcbdgMDWYGIJLcLhHfwcio0zL/xLgc1x4rk36bVXDDwMXa6Cy4/zNlzC0FrP
9dT6tn1W9a3dHrByihbfPJYuTMDHBpj1/QdyIQQ85uzqf0uc57APLbtFTwXRV46vEf3zhNprgtna
aoLrdin5YZgq/m4chjgXe+qEL3Lp0kKzDA8UGdTqi8eUPaNL/O0cj/YanUrYF8XvdXR4jN4qWmrl
tow6ILL8tgibYUnJIiLn6xYMnYie2kCE/eeC711/eraPbREoOW2kFKwaxYssqe/Z+8os/Rj2RM7f
5CDELfzuPi5+hMDHq+4ZN6etNHN8wzXu2kOEsCR3FwUEkTQ51IjqYj+1pWqHS0LOsqEii911KKYw
7zCHYpdPcBikVNq9IslDDX+02Z81TRmjdxYdTZyStgZoKnP+LHbJS84mD5izwVgoKBa1Ba/9FpGn
szUNv5CX8Vx2K34OJBoU4iCzRGGq2TqfdgmAOJPDKH8aXptiRhZJqYig5us8KIZHng+b3ItEKDNR
Vypyy96jf/Miur6YM2rsds7vqdAnieAY2YsShNh5Fz083dAQd5gPeIUXkovpFz2tWY+4p/W7m5uj
bIx379WScUO4/PRIo5tbcfI0xoxBz37NyLFBoDs1QowSTy/ljgy+5QBcn0VpiulmSBz2tNdivhoj
ZmXKKyAU+s23+PvZzEN62buoKQtssjnPTq0avf1kbAcxRgIUJJEGFjM8n0QQs8AP9i/xEf5BFxTD
+fqINl+NxZWlsLCKt+icX1rYSdWA6hIG7T7rcVfZ3qxk44UdXakT/g2JF0d+mcO/bHtchLipkqDQ
88AhYjO8/zq8wpWkdIrFqjAVOvQnC53NhY4RexBByTmkHDvT7t/upOc9S6x/+NJvJzybkMieAb0B
/yEusW7lAadEa1fi8cWXeiceABd1A026/OnxdUMLzp8zs+c5XmWV3+VI937kCF04mQ1L1ZxNiKSM
sKB6XjVjPQYYOB7JwuHKpSPbJKRTGFjhbLQl3ia1aypbLyOgj4BD7dBam4NBLo6y8cNzQ6JlVbOB
pzNcRHAHc1JJ0kPdE9Alf/t2bjvw0cbPViZ5IoBEU5y/SPUTerB+SAxl93947epoJqxm42VpTgSW
nte2aByTUm0fvwCAvCnsNCOyWExHofuQmYY+cnvZpYbsng78vInyVFGCYYTw9n2Da95ak4OK1FSa
B2fPVllEsozV18BvaDVinNfYGNFMYfD6CX0GemURYFRl9W8g++xHplrFWYqcxf3ycXhz6Wwb3SBz
WY6QCxUXm2pO9+wwJXweTgqkXnuWOyQJNkqyE5NFMMx7CH5MPyP+XnIbjViF/jbKWO9HimpVh9e3
as1T4tzXsHaNmy1xNLz8ap1qor06S2pNuR4D/s0XBvc+/ulDQ8QpDtFZYVKYzLiEgF1edyj0IZpV
33glP7zTn8Q13541RVC1V0j3NsUmys4iDq9bZPxU/bgeeI8/Q6N3O/PlFyBedcV2KNbErAz4IWC8
T15SldmM6Jq0vjR/a2Q/bLR44wvmMNwVGvj3l0V83/9JHJQo8u9MO1P48Iywx4aPDIJMqtYvNMuM
rJ2ez7tmft+Xp0uAKNyS1UGAPlrW1gBvRNJjeO454oQvg3qxGH0Un+MrNQXlhoiiQTZE+j0iiw+t
zeXfzvwoLeaFrYWt0s48XYoEuKcfvjmHnoWazai8S1a5/FbvcBvn5oOdJ+3lBQu0NmoqEtq0zoks
mKeBZxrgIbfeR9bxsX7iHwQEvVr7I3LGrKhLw1hPO0NkAXkfy5RYZzGwfVTUa54H2BCTgj5GIgik
6aqSQXjPew5O9gs547cqvy+AedSsUy0IjByCo3oMhyUrapqfxhDo6o0XEMTWIhMgTh1amz8ikgnA
O65K9/6m7UD2zp2V1xIKXgB2Yjmqryhnt4OCEBfz2xIjsgpFQl7Qsf/SZWnCWf52IfDjRJn/L3/L
jUdJcJ+ST2PO5f+rhyiIzy7nkWwkEXQNnrpxO5u/aHLnCMrzIg3DsfEkbKmOq84iAspDUdptmUsz
8ZObYdGSxt8DlYosntGMtBpsqAFubT5l2q3EfjnOUvUP7K+U8AbBt8htDMX3Efe8tic4wOYZd8O7
0LsCvBvuoQdzeHGPTR1+iSmgpPwg+9pCfl3/DUm3QgKiAGYk1tPhaEmYqs8ObK8ceWIn/GKsBAiz
ocoMU5yNbzJleD8kTTeubmVxQvQVBht3uVwh6S5eeV0SUq/3W6HGVCW1RF4jUsRHXYPmN+G9szGI
7aWaiKRbGR6w91q2Qr7tDjPmtnEBoLWWZ3K19eqY8UbidLn8UxhUU6hddlpDxrRYLSN2cAcApgfZ
/46qbsEOi8RW263KIlysab70iPV4Sl/UQH6mNjRq+uwJnMXb1AcWBIf7qMXTmKYTwrYw+0os1p7T
8fTTNRGifm05hIb8f4g56csMzOsdovtQ3RIVY9du/D/TrOaJti5mWZ38yGYktVb6xNNvCXRMKVty
D/t4O/WTVazRfptzk3rST9MNvbI288MuUoPVM6RpnzZ37eQHtELchGktSnpTQIeFnzidmcMKfUZj
3JqvR1Nn/7gdGG25veKJSo1utAuVHNtYnfksNXh6sKdO1lMsZj98Lt+E+mQBZHYZhzCdMS8j3RBN
yPjDBOHQO5PCotu2EYRzZot2JrkFrlZm3Tx82SG/J69Otcg0TQd44FRRdS7T4qidSvpXfdigEJ6a
mnrogaqTSQhbZs8ip70njXK8rHldXo48pJ08rFZX647ip0ySWXtfigi1tWoc5zgvVA/sQR2cGTUu
ocIlmc7GB8On96rhaGwqMH+jSfUeZfusXF2j++UIhp6dpZ7VtOvShV739GnfBXIZeTqD2sv/sGjC
4ubIOntSgJug6cN4AX4XkqRh8erkbYy7pJluLJoN66dtwi31QYOKYsdigASKlmYD7H6GXzb2VV+r
UNMqMbAO7zRDA6iOJyE3pU1ruB+zxAAjgQ/qHlW48zRilKa7JoemLdnddMYaVeOzrKNgG7DCXP61
zJKPgjOc2B6AkifXvewWjIJM8q5g2/VjVwJyoFOxq9XZCwngRw/rpPoM/t4w7KUfperYSD7WfmCD
a/QmNvYI9MUwgysKlJJakVlG9n323XBoGpZWplhCe/ty6mZyBRBc76EiNZ/DqY9AvY/nBuqV54gl
fnMPS1rUwrybA+alecreZC75f+R9M8p+mxl1Dvl4uMUAu6fv+nopgLWi700LmOJBl2evz1vsA5HO
lKOclXHHzvNhEu2u9Uw1N5R1ocqTY0WOKCIRAM0wMC7g9RA2t7T2GejdHXwEPW3IB6vZGYW68P6j
XfOVKfky6KhsNkWUkOz5zl9Ko7uXz0/Uxehps6D9rfVuG6fU/oEr8FcGFpuboBHM8Kyvojv0ej9w
CMoWllPJvloBITSRYcBgIN32Yq9HIGDIZZ32WRZeKRosxqMjgHzBjzzWSA4ItYhm5WNfd3T6vDhJ
BB1c4Mb6OKnZXvjghnocZ5oziXZhF6j2FqndbL3W/9gPB64DaMdXNt1HABIE5UqbSEDaEpRvSFgS
jD9PONl+vZWMzdNKTvs0aYdSSU0wdYfwuVsxqiXo58yyWhba8uh7dsjKq2tvjAv5QpjX38veGrRP
2LYvoao72Tc2k6fWVjcD/m7oBx6MT1jaGNbo3crBbuYxt2jCRX1Dp+N2aasWekse8L3pR2NoqArH
g+WlWO+A2/z3YBbXKTVvp5rhd5Qi5lrJFbI6qnxHRyACaVJQTPab+4Uy/MhruZN/xqfAyy46pa27
V4gsQh1awROlagLR4qlQjk+Bhtvh7+YHlET5KBsCYbx36j3ld93QzLIWWiTjdC7TaFn6ucL4UIh5
aCV6/aN2G++ww4h7eRjx8+eaN5nlbCT1E40/pHAxPbMTiR5fJ0Wf5uFqWHL5uJPmCG4OVudVLoRf
qj5s9Yioj7CHwEAcOAZfs4BrEXTo3Y9LPR7+7GxqlHXRzBdIW+LQc0I70jEAAHilBTHST8gkyB9R
gwR0PYX+xY4OXvER8oQnJ91pKfIZjRytX9ueOqndUuw7hX0krp8DH2ZCS4Bm5jj0v9mzLTccO1bB
mxabjCbK/Nmz5+2NolRo1BOUHFYGaW87YEXl7yIeyUbPu3WYXeoeFaiLz3ZCkpl0lZMr1I4GG9Ye
H/s5C90D8TkezZhPHjjb0UJgp6jKILsnKeYk8uteFopGPkCpn5lbvOv5pG6RaqaYJp2Hke8wiPYi
jbKlAycx9KVSK+R3jS9sJu2MNvnKSlSOYQBarrzUGmS25oGTFioNR4CmmGtVUlGHqBiGbj+iqVDt
WmSIUHbtH2fBAWU/PiAnbdnSeLGXoqfBmgKJ3K2H/jJ+9CAarnGsm0k3PPzPLjd2GmqRZKrtvEZ9
MP1ZVMr2fHDdtRrRL1FiZcqkHKi9afeUzav2Wub1EnOlhczUdkgtaIm7Z2O9/3wJwFht9+JkEVNo
3Ph7YbFp0VHzVjESJUFXuE3j2CKbcgbvefGtBN9a6FW7z/SJ/50W9RbsQOFhjogFEmgrJ7cQUs3v
BDgdYolAZZZtxMKN7CoTFUPF6wK6zQKpgHJRk4nmSE15t4f13JAlpMMLJlAJXoLp42tZw2DeXmn5
QFGtRK6T0pdDhn3EKCcE7L6qbiu1pKeYB8dP3yng+GqvNGdyyx6iXSQE+5UU66GZ6yYDWJLDHJfI
2pHu8km7BBDIhr4gj7j5+wLenEwm2H3siXOLZ/mlqvLFX99nWG2O23L9hdk/FZB2zHHcY7je5fi9
az2S9gFml2wCP+uYojljSgE0lLILv/N2SWXxVTu/RjkF1Mfm1sIo53JKyN+qwmFWK8JBAvJXQXNc
WXcBqq+ytubly2sVGqxVXPquT1ZdwIUs8InoJBu2swz5xkt8JceL2xmJLc4ogyQ6Nu/n9AXQdn87
XHQlQbg8fZhifUW0cssqV/eqnmYHZKr//tJgK30qTXNf6flP/cLepyRitUvEozKqLcaGgh+0diAs
eN5UVxC0fwDAyHHQxx9HEzn1+xQXyZJXQYDTkqPMkafyd1GP49OdhBXK5kLR86BwPzAEFUViOJzQ
rlnGElsHIdolVhn8ZKLkTYmHpii1Org8VW3wnTLLlFGz7o0YyRiZSECzfsEv4MK5iLoUP3bLq7hB
SzvitWwKzAcaBCaz/SU8GDuNH9aTMwaJIRVkZWCviL07ykjDzGwsnNhI6Ec9xFNkMc7Eyzg7Zmtj
zxsCD99avX7S0WvXLaTSghN2FLGIGPuWz2f1+eGJYEtj+wn/sux630+VFs9R7o5wNR9U8aLyBbh2
D7UHxol1DG0eW0YsFDMNixuhs0rq/PfGTbl8QJ3+Rz0LQRr6W4uh7RzpMjVv6UoHXThkeNQ1n2T1
ouYHm9SnS0oiYARM2P89VuSKt+KgACMoPFEdvP53WdX5XFMaDXR/jm+RyN0Gw+ASRH28GO71cLUW
VhEsdM/1STAJo9p9QISpSW2zUfO5aOs6n4ZIGq4ZYHMkJhdly2EhjMvos19J+lbfy5ldQueiC20H
sDGQVLnunQ2MfUp6TG9Z+Hy/EqZU6xoNo2yOZ1OIxhBTE9g71mCgcWWqFElzehucvmMaCfjwF0Ro
ZCDMV1kIvd3CBgZYwJL4p5PLJkLM+o3vNi+5QMM4FF5moTCYNRtBQ07oidnl0W0Cxyhf1K1gXAeb
nf8VnU9/kRukXhvtNFM9VV/76FAaDuZ3N2h33F4HGEKKQwD6CRAbcNNp/IBND4ZDZbPPtk4u8UIC
wPyYfkaI0YyFK4EklutdnZtseNn80FcO2wH+3AhA9oZUd7YHHv1DWNKlpteHJyoVamHeQdnPu8De
sVA6syYR+XureRZRdpPAytDUUbN9EgzcLj5w4k+8gHwLnt0gsuJHiPJcfNXLPa+wJSsvii/wBCxl
6LjG/k4na6nwuJusLyCKsWrntzK/URdWWaAIJdHz7/eQSjzG4qgX3uNDgFkHy6YxwSLi66Y1PU10
HrdbrpoX54q6BgUMRtfAH3+O9Dm3oa9bpcTYxKe8baAxxBg6vWbxrz2Rzoj0jA6S+TLvKbbEDhC7
lhZlh1q12UqOy+I3zFI/TRMh5blqWlHHcs1xlumvUf1m1F9wDKDuSDy4ZYPs+KmXRUg5GWcWE1ec
o50iWNVkOzIvWJnPLhwNG0zeB3cyYK1y51A93+aLcHV18Q4U/Bh/xrXTndX2uWOLVE7boRxyd9H/
m/LZEuT8epbZbfcfTNfFGyElj3BW8mIWl8uQXHObt7wiIMiqwQwlVC3AynJX+HzpHQAxwfu+uftb
Qkyq0578Jtxs7Cq2O7brWJBOy0CH4vwRiqUDBmz/4FP/H2Q1tdmnQ7cD0q800zPvPW26RYkGcreI
LGbAPF4gV4JEHWZh0bMLswxPlGoebYsCrVU0w/oZeq79SWyxrtqdcP39OxQI+/vizNuaAdqzw9vp
joLF4KkLc322xlVGEohKCVGsak1/4mT6tRGSyENaa8b4BDlVjPfnciL+ez0KD1S5rBrzd9TgDcZn
akL99VQIQiszHBbWV7VfIrwa97CWhu2UEdNzCOEmTQ0Eqmz0hVfw0aDXTFsbmLjJ9fFzosqf8wyZ
2jrQwOpUz8eSt2XW5RgKcS+R4olvqszGJQuvFi+kTUffs21AsnqqQpss1D1zse24ceZRZbbU3bS0
ubdAcGe+3/HcnJqGZ7vNckQY8aCpNV2RuBfMIoictrmrWjNHmOkcuuOaBrYOlGA0wyTCeArbDsXX
H8/IdAuQroDgONaeqCxBsCvBN0S4EwxdVqz6/ONJ9jKi0E5jMoo+9qtEBGr5pvHsp7WqRm0KQRlx
zyCmWd9BXs7jGKW3zdwG30pttCGhKOVADCt3kJrLLcCZZJvG1SvQzMQ4qUSAIHWRT3voJF7q10tP
duidQ13hGHwnGqUqnmsu6UIy2qA0HbupB/cuQYPRyn5lOGbBYPz9BkQyRoA4kL+wGN3GgVd6z4kg
vOAw87IW16bFyUfeS4SCwhb2ECuMElE907P/WS6w46W6qzuDBFHOrakjq6shiIg2Sa8HlXZ0iQjc
wsSoWOfkKVUhEwdiLLu/S/wgtcjLShlyI91dNpsTr3LSw0D8jpW5Btqd1y7kEX1S6Wt5GyDNx02Z
jxPUYt16dLGs3wmzR9YDej2azgltiSrYJWQslK/wAoi3EQgRPuo9Vh+rC4/J9g6YE6tDPRjz3IYn
tn+9C4X02mxwJ5NT0qLQEL4mij56E0CX5zDyF5hXsHsdmWi8KWV1pC8RJ9PvJTXPvkapm76lJ+Ci
fn7ieCjl5hiBoRKSTKIhSh5Fe7TKvYFwkiNa6E8ccQHf0aqkJEGHTccDlVGwEtTLTn9psTRVhrJN
FnIlvfqV4221qbX1oM0RT2tXmJazqYFcNVhp11THQC9/Tqr6rrMQilY6lf87bQrijmwivYEiOStR
s0/6QxTquGVBDtcfpI0Vz12eKAkfckY3QezmFuFiC1IYoE/gBl0fpiOo/ew83ejDz4/FLWAsFv05
tvAiBJ+o8oPrYj9yzSjL2gRT6siV7KOzyni8LyOdXsS/xADyDSJTg1lB56OhGNuUOLuZdHYvVSXD
KUE/bIIrPVjOm0qWC48kCje9IYqN8G+s/UuOodmQM6IFG7Sl9lTodlCiLNf/D0THeFfaOqTuGA6Z
+MNNjfFfzNUd5JUHqeawGtdhmoelOKWMEsMDUQrWvIHaCg+0mOWPufAx9G9ArKIEo5gHmdd1hUgs
O8UDzu3PK44hs3tffOiKT7NsWbJj8LkibxnL61rh+gHMBBemrTidthkUL1lboOb3hGwdmPO5YvQr
RUPXg/PSPoAIH4OCtzrToh+VHuTMe5r2+DaMXS0ewva+RIFu9jUTVxhZSAX/t3q901A33aXa5nLJ
WYyVugVvjmBLszVJ7+jGgomM7iXPwswdPbq09EAJKWSPHAfDMetUljfHZKLft9tE5FTuV4fHSnoq
WKHI7PG5OIFadBh3LRXr4RCZrLUsSIYicKPwhg1TSIYQNQ//YZMyxymi56hvpFJtY7ecSiS3gNKp
+qpb9FNaSRhMdOGMLOdq5VUYPLokDHMVLfYVaBSl10D74GPO5pBqM59VbLp+fmlLN4FBM4YWL3p2
0ck38m3L6/ff29SnnAODmAaGYctPA8S6KX7FNP2YcNdg0beRxM9El80vTdB7bbTFBxiDrok4P8rx
EWuQE3gDQ2vv+j4IlZ2RjNpr/BKcKY9VFIOnhFpJIHXnodnTjKwXWmdbVSdPxPSeDyqibj5CcwIP
ddSErZ8Rez/WHMXpQoSoqlfL2Mi/VljhE0TUA+vjwFDSl9W8ZMqcsOEAF0nzOppbKAjI/c8KU/8G
KlxQh/5/CnLwj6uO74yzxdnqqm0qc46l3GE8arJ+SOb5hTl1ET3dGGE2JRBH+6IoDy+S4iOjbWQ3
kJKYStGqDUed63Xqat9b9QcFHsPgqIK3EfmUg0gKGmCBcoD4LTNhgRpVNVf/yt3dUmd7EmUC7Is0
ZFTM/qgvAGp8AM+e3IZzJH/Lr9SwqYWGh/fSx4WVC98S/T4GaUhHJQ2VRRMYaUUYg3wqFImVeQWx
yNlm2QJ0//BM3Yjc8OpBa43iYJN187KqC1KeTQQodoTnHYju8S7Mct1N4fTQGkxiuzq5mieSUMEr
G2JWtmhvYKqXrlc1ToclTKJ+ff4PKnGG1TfPbu1VNj06DrnYQ6oNGePDhvp047FBIXM5y1WXOp6q
+h60NfYlWzsAHBk673tuapu2omwacxLtLxW1Y/oDanqXMttnRaDtARrhwVSTTElCsQNbv+izdG+u
RD8expcqgaFy1M7Vp7XORL8Fbk6PL04FEG5Jd4Svt3Nx0eCTiBinF98DAQfl2qt6trDOS5Nuxz3z
Xpa6Z8tqd/j6b0hvupVZ3ZTRk8EcTz10kxaGZt03w8HwZ12RsQPWbD+dPqRcp+Rptd+wlPO89mth
7Bz0454TMjcjR9oGVL3QwrMN2EJIPsyMhOfSPUDNF1I9QCaHwcAclG+GQOuETYf1nfzoW/Ny6uK3
j45tKa0VgeHN/cWCN6B70TmRPXhUqaTyMHJ5ji4Q2Z2UgTkzvaxksDKtwTXTd2cXa32/P9/Ctvwy
m1B82iMXMh01S8RJy25LmJN6GMM4u9qycRs1dVVtcDNlSEm8ANUCmX+lp7gyzJ8IMhxKWEgZVz03
BkR0zM2AczLDwbk9LwByV20yUEESeoyf5Og2/zD0yaeqfgT6b3sgAACBEFKMp6lcaLTUrzv+lBX+
iJBvILuwdDZsT+gnbxSFWvot+TM2CDEsZMtI3ho9v7EE1UTLG/Hgglc0DCuEYEHh349Apn139wEq
onUm/0ECv1bv3f9pyFqtZvXxwyX6EIA9RZKon8sZ5tk3NNjCn35VF2zBWe1oYfoXI3O/h155gCbn
3+wdT1iCjMzSSfyd6ZLHu8H5cfm15gVfNPAHUP23YenP2xEsImBS4n0DzxdLGZTZkfAb1L+k8n+J
OD85sGXK+mNNlNVt5+nkmPvXfbsE9qJBjWiOx927FwE3eL6SpNGia4+4ACs6w4Mlm+YGgIJ2HtAQ
xqh63Dt+2nON2FXr7ctTOY57iRVwdlKWtzOYqAr0FV0yIY5LL8DM9taTz+WqcvWOSQSBsolrSfxb
+xpgBTf3omjwbkO7LgjsBA0bk0VAnL7Cz5ZkK8bVaCmajCrcGKVxSLrWHb1ELJlVViS3qrFVzvAz
owPW/G3Fu+975txgAaldzmBGSqR2nnfaDm8EVTB4IF0wlMZGR+xxx0JftVC0lHq90xTy/U69KOZU
pOFVkpHJb3xSrnyNwONNNllSkQAc0nDZLO4G9PPE5Xo2kXaYcihtaNLOVC2naYvO72T8E0ggifIZ
DY4JHPJtch0FhsJM6MH9HCe+Oo6ymfi9TRPszJzLgJBa7g7Qq6khuU8TEG7NbMgnsy7swjO6KE7T
mxl1vUs/r7f3o1/NeZjHkthULv/ztCfDbLSnaDzKpAqXq6imoCSCgsdv0+ex28ns4aZR84A37419
1UaoDZzSTClkGXeeKnUU5mOmKA4b/XugxB1a7b948/1jvGN0U6eSK3S7j4m2UyQoV/3thueJt0c7
91cANazLzBgA/yK7j+KaTv9QAxgC8PE0gKl+BDPm4FmpX7UypVAKwIoHXS8mZjUk4QHjldHIjmo1
6q4uK5/fgz6vfcUhNsU+loZemYd9zrAq6TozyW4/K/rtdDpDWjuj3rOafDR87aDqrX1S5jSM0fAj
PBWpP2wMqEOisUEE50vfAP4csr6dmhwj5/23g1eAy2PuTu//j52sd/lD9+cj6rtHmZ2onw0A6g9u
m5b85dgrD9YY/E5XuhFnYKSK9Vdrz+o8DixwQ6pqa6QHoiAlPuolYfI5FE1JpUo1Wy2QUhsmY4wa
ptIZKh4XS6nx3FyIUR9/AV0EMJHP1VdWp55g2F+on9S/PwyeG5hZo+EvWKPlBzHr++H1jVDzfGty
7eAA1IOfm7xKyTvG5jwUjWqJGf0Yp4c3/JiFyZ7jC8l4W7aJmWfE+FMMtXoej7TGF/eXmsrWMsqD
Dr294qk3P7NVVAFTB0GYlWTsryaHFQTeILuxMbINMd2UOgPNgVMpJcVvfctGJ/y5/IjF9sxmorJT
ex3FVa0xMvNAH3okm8XUjt5R/3Oy66QOxriqglxeoQW+6inmmFIggsj9YlgOtOCR+spnHPRK8q27
YypZjOC/ze/n8cnLkjKEm+cAWZJ4G4Wv0cT18P/ODOaN8GJxdAOrN7vikF6WP3yvj4NZvGvdWP7+
4GJ77WEft11ftLlSfO7z5vRnM0TR1bkDxBqf/MnFL5c2eQYEfFfC3JPDQY/Yw2KSAXApZEmtXiD8
UFycuUSpUBvE0UnNcOlT6DPJ6zO9dulEhb1QL9kjNriS2zKAE3cVRRAGz/fZ3OPr6/tLHIMzU2km
zle3Cx+y2mMa0DqBurU1lR+sqMmowUH8K383CrO0hfTwtpQIszftXF1DQ4Em5zW5NSaV95CFcYQF
fj5+er9oULWfFU42mGtmbhsh4T5wq59G1Xfblvcjntr+scDAn8UA+lipfR8Js4MhHoYS4Soed2IQ
29SZ57PDxbE8vcRpO745e1SYM1Z+mITrv3pPC+C8vl9XlcWI7UAL6wOAZzCdyE7Tzl60Fp8ZsuOR
69DJDBYlOTQBriZDrcI2pRp8fAW0UhtnGXzWGMQ6nJThKACNBjaHtvC7XoxVOtQuQjSV99yM29LF
gO2RCRn24GKKtadPV4KxvuAJGqDU0NQUpgUioCfvgMwpavRbCRmP2MNmhDdtm7i7gOZtYFd+zHCV
lpCuVftj00PrKKZAGmK+ceFfY3TzHVIVVuqwGgiq6pBia5Un2Up7oStZq9CdE5O39pH707SvkOqd
n7dfjG+E8N5zKLJVONYImsrGOxdmQsrcGySlcYII4QchmoaCTo+C1K+MAWztLP1XiLBVw4Ylbb/u
JCizuIvFugGDUG92/+yYWyd244ani8WxYeg779nsLaVnFAMHoBi464zh1B25Uy/mfmmdnK7ONeUV
QRXyQqKv/A/aLG/winHOsmQCDMq/P4445wEVaVx4QJG47vDk7SXPVEo01HX724AEhH8SV+4U4Yic
MEVynWc2lUBKEm40iXfBSHX1JHLBfefPAS1kcctu2QR8p1rHR+fDHwuScry8vghBdE3Df8xKtixP
S7KDJvxIF5vboOFTRHR6PPnKB7m/YnjKjsR1sGzQKYTM9IIOY/0cErb9BAmJTYfHXJjNQMTSd+uA
LPKIpjLElqiBGqCnLq0eXXzbIcAva/R4cMRpBhsQMiOd1N3RxOR6rb0ecGKgpDqPWQRBnPwHkxyX
DlQsOz6Gjiyr5z5vZCiyUB+3Av5TPygCKv+eJE5nxlIiBMpQ70JdYsONbWisxA/HpZVphHnCm1M0
FYGbPkyaF+n52PY+yl3gHPDltOd2jH7lWPxvfqASs9fs8izeL6PpOt4arO3Z0OHJvY1dH+96LScR
inFhCwI1BiwCIQ/OUI82R2uW3ATofjTgSk3Ba7QvWVO+mCscZlPD8N3o1j9cCuACznaqdjexI29z
zZjulCLVEcSbta6FAAstjt/kS9EKy66oQEaF+792SrwVX0rLES5c4jXhERmkq3wQFY7yardZowl5
cfwZaUzIxEqwhrM73nGarnRkFCwgP+eV3cXAee2Xcmd9ySmObs0Ys1SybM+0P1CM7c+cAkwMw9dg
mbtDX+LGbbDqBXPDwH7kTya7Zt5qUwPKSYYThqb1MNFZwhnjXILZnrArwRHyJmYPvPhndL01ncDG
iZi11b7HjZ58v48BmHs0eFq4ulU4NubA3NrjLPQg2q5jHcQiC4dBsbBVdJWifCciZgBa7kVn6S5o
5qVmhxd52Kw0zSDhDF6nl1BGxOKGzrgeK1tv1fMVmUrbAlN3snSVhI7TaNzmP3ndnuP8cLbJoD3K
xAr8xrFKuWP8xursNqJSiY7lEC7pIOZQQbXZeOlB8mfToWlfUSgtQRv3V+Dv9uQ/dvzxpFDWBeYs
Zlz5mzd56Z96kB15G6pREg374mxY4jJlDZ6iQ2AFL7LEpLTSjN05elKcrutwGwfVXz7Rndjnq5DM
1hvJu/EoA63/SUKUnTlSAY2TgsBRms+nCfUXfil2go1NN0GtKSQslwEmJtkIHRveHH544pYAXBob
jND9Num6ttG8duwVPON9ZLP0BRpkuXznsFc+x+0lkDZ/ab/Ivd+uqqzzHrUMezFZGgK7dC2xMQyJ
g9zIeC3w1FNeZmZTu6qwBbTKtuFjxD9gqfNdX2osKxCTqXIL/I8oWGHor/znpsJTEVzrSOsPep+O
l3VOgnpbk71hxSaeBzSTNklQiPcERv+nK2vwW/XGzYN+K9/E1UPbrLZoZGCHsxn+dBRDEdVLOSpt
6DYoKVDcVtyW9u7SxgpPKQQbn4ZunKhBfzKIM8n33UxV8pswG8XU6p6xZJC7hFTai+hc9BpsZMRw
oL6AvUGY9NSru0jd6yeWZAMFOkVlwjZdIoxjdgzcK+qQZq3SyaDlRFhemrfoO997saBeLm2GEtmS
sUFyyiTmcXNoFFt/ROe6EVMm6eRGVnItZKOK62Ah93afkj2/GXi/i1rFe+HcV7VRyceleTPc3vWR
OgFu/+lhxrFLnPQ9T/NKuFmq41gNixlNx6vjkQFXAvPXhvg1+8ury83mqG8uAPAkDJTDRGFyPjPw
S2VnhycoEsmxtN0SDQ2SFUdlURzVX4wpZyn1ar+XIlH+CZFQG54hTrEeUaMNBvSndra/gpK/yVLr
+FwGIvXh+MOPKMKhobVfuG9i/fTi2+vZwyDZUqi4m1hzMmjjwC6fYWKI96LZ0o2zQv3IbRaWmiEi
q6FiS0Nuw1TysHroRYKjW2bcUa1zwwDcAoT9rrEpLrYknGj8D4/Z0vsj2PZN/LoBujzjXHhyf1MU
zq0zjigFCTFB0GIxuNwjg44l4mY/A9yVAFBNuyYyL6l3UtJ9hPVhLk3Q4UNU4noFPHNlhFV2klYU
pgZRL5vPoHl4pVEVsYGmPvG3+dqZUfHXKCGKizTiZD+WVeVp7JCsU2nJNksbF+1dUbJ6e5LtIvEi
VepeSVY4ZWjv5+Iem65K8WZgr5CBtAMMWLNdxgv7fMffQ8T07zSM+jjo8rIpFjhGUTOymM0qcSLb
7GRkp0D2vzTdYSt8CaeYs8tZi3QwPzlQ7X/8bHk/6lJnzC8t3q+CuQjd7+MwqdWd2tE8di4vkF7k
TlEyi2ggsvasUZhi8CHOL0WIzoHI9ybiKp+pDN0/PEDts3mFv+yBR/NsCRvldVojNWrwWsINbfLe
eRwi9x5S53vxNfZnEksYnva01RRu0E3mrUDtOwFDwWrHLXsSbZ3Zwa3bqxQNkTSFpIupg3LMlO88
Umitx8P/mG+tpTPelP2m1/nxE0EDIDgkpHi0en6EdGWNnBfhvrJWEZjyUsHRhSDd3ia0rmPUeMRN
NjNOvRuz+mfjHncvtNfHdC05aXzjH/CYi2fY0qpztOUINR8UkQ2VXtzSlI/FkQciZwG8ypEkURrj
5X/Al5QyJoNB4H1iGDPXPY1e4YqkHsIU3ZgDL/cqxKahESsHf2nmrvLAYMjdYj80qM/95cKIOQYU
r87RYlSejuuZIszOW5xoIug9JHRsuQAaoUiaDvjegbqfYxmzKJTedTDBwq21xsUZZempsX933i04
1C7i3FkTOgP47GigrlctDwIhqjNeszkeKKduMVtLHLsGTifjiqC1M/irULpM5fqrV8H6SU81XGMj
+o1DDAw0d+20P613dzKFrfLqDVJ3/dVmN44JwUy5rEwqQVnRWhaT07ZpRg2oMMLWTMqzob9sAU5n
ooGrQOmMb8+3oNDQUF0vv9q+DvgIST5agd80107em1UpoYuAdVhtP2gOXrMPR/yPmRra79ADcnVo
IEe2cmYp3z3AqECr+qht/OPNlAr0ZngYImPQW22qaMbQFcG+Lcqq/w858Zj1FIOZFrdmiv7h3kwT
iNjir5l31gVALSq0TqrIIczm2H14NwokIDgDzFfExpxsemrM4INmCzlkFqFzrkXUvUbygVkHO/70
ry67yUVFemohwUH3eZpFl4nYs8dQ4XJTzpL+txe5GJ+tUXYUxn7L4JADtN/37yDPRry4SMh9TwGw
VVbt3gM4srvi8hIeuz+rk81SUW0DaOhDIiKcXkHH9uAsD/7t/9lbvE0GXhE8LYagVLKoy7zJVGWR
B0HUvVyhfv0nW0G86gimVwkRAUm1cEUKnRvcWu/BUTcuqumAxYC8HruM1yDVnJEOCX6FnWZ8Q5Bv
2IDcKl8dOZGgg/dAM/jCff3+qB6S9NNf8dXnc8ZMqOYzXuAfbdxqXFjSD+sxjNyKmF+0W48mhXJs
WkoGADEoLVLgyLVSzRT08fP05tI0YnBAtfSC3FKJsGe2yqXyC+HcbfSNLK56LJG9nBIp3qA2LjnW
HsvoeQ6hjczMDGp6Sv+lgKv+0hDK8LlaBujixdXiSguuvIDJgYdkcvS0trg92RySr4mVdDogHutl
GhPXVjO8vFJISXlWk/z/umSP4FRBe2vgGRsL6KbuHSh+0obBjQIO1IIKaEvAdSalyOmRsW+2KRns
5zFThdLoFX2stzoxRhK5hj2hmWwVrkzImTgZAzNWzSIKW6ZNbodgjTxvVpv+q/Kl44Iwa5+AKIzJ
9kZHxELd20m+AzKQVqDRRhu2GYNOKqzKG3nZrtMZA0izg2renKs3wZLIR4GMgACem2/gN2aYUii7
wT2AdBKmJfnBj2/NP14LBGs3QABXk+OsDCpWkDd0+05gaGg81RnwaWK9SdMMfH7rmsUtyUsHBOGd
COXGrO0gyQA2tMM2KHZXHNB+6K/Y2Z8hfWHLAb3vi/hIIuWIrjd2PezRNCz7U6ZywbOvD7ac55nz
pn5uPKItdN4T0P4QSpZSWwV3TEcj0YSLwJR2kqGBuOvLX6pzdEcBtb+iniqAsZ8Blo5Hl/EmAGRI
BMwFqjURYpcojrF22kXpo6uZQOkHnkLkRAc2YBOXkonUq78gr4Y66c9zdS8NGGtcOpjSfjxmFw9b
G9+fH/HHPQeJ9Go+KtqKG3Tlv+qffTAtwskOnLlkddVXt1y8xuNE4uQSAmfXRXiDenUPrC6jS2hq
SwLcbVNLPSOI0AwTihWqcW8CMen0k5ibvbPaulm5TejFyAE62Xf0ElBaJsb0RKt3Sqm7TI2pUGtn
n0yCF6Q2Jys/pbw+4boP1CnnQ1cfO5afoai05EPaUfQJQB0Z/Bm/zlopCvN2B4kFqHYdxAClYg1A
kY9VWq67MlFSZr0o8arOl8wf7oZmfULGy5nD2MI7lNQ5w+CdAoqXbgYZ7G4sjlKXYyko0wrzdK9J
JUOlvs3peu8LEf1yYTA5hotxp2P2VCnAorlMKq/52u7z7fUGeZDH4l+tFXv/0lmvQHFnkvtAEoqs
RFhdwJT5T14i/jadZQBJkWNKCVR8z+c2Heh9Asa1FZ6ndY2iS4yCPMdKqv03kzJIDVVoNuCWTdgz
oe7COgcq+dHu8G3ZJa2EmvLYkl2kAF6BXYc69UfgRNedZeetoNoV/LTSnNolDtq9SJ0zWuNJ4kvW
bUWXmV+x50FyonfbhzzP4gY6eFRq9riZ+RDv5jPX/tXOSVi/dXqJjMFFysAaFuyhCbtEIsvGMd3K
bWsa4MJTskNnHlNwj74jIf70+M1ns4rG4c40mnKr6a9sUgbUZNXk+uRN1DdYbL5a/5iBTHW708Qj
JWrUF7puqPx7U5yptbzOVv+hIqCXTm3d/8szgjfKJkhRDWo1nJ55T5SREjZoaTYpVHNLDkRXs+FH
UAvdWnRZvhr/G8Qu+6IFU7XDoMiZyrX+8Wf55xpv1+HI3VrWwOIoFXjpgikIWHQt71n6+SsspI5O
JgDvmCutKRRBkR81bCWLOuXqzA2+6DYIMJc6S1mZZMbGmZRV3p+5lBIoS73PW2fYCLRdbv2ZZ9zV
FSCsl21SDE4o1c+BIdgxhYI2+y0cfQHNu75svxhfKYsRhMmtySt3xsW00Joi8sDzVutud5Px26Mx
0W9bfNXMVmAt+P1eK6peqkITGVSy98Hilsp/DYLGFVeX/Y/kcEAv766eD7a605nMyP5rxMhX4e+I
q+xgfhIr/IJ9YKK0yLMy5oHHYtDmELDecGbsazJa46sRP5cbpoIyKMRQwI7HebCbpAu8T3es2OkJ
fqWmeZCJMvKZrBWq9Fx+mKQfGI6c4QdCWJavpCeUywz8DUhj92cv5Q6PsvUeCf+KvCzbU3tZKaln
8k51ODZM437kKXrwxmGL6DK7fVhzc762kOe8P60LvcowhxKe8IaR2Oeh4H+/E8ZOhTKoETaGROwE
iJXSe4V+0R3DO/+DQFuzWHgi3MYUfBe320QCAolEOmvAT//arKhbGIP5XuilosDS85v5k+wGSIBu
42MoTIjjyaFgssuc5QCQpVKuNCUNBZ77VwFVRXjVy9BFyhVKTbSShvbW7XS/IqeVA/Fmwu/qjf2+
k4YS1UrC/3HorbEWL9mWALbRq/WQr4+wOM5HUdO8vzfgqXqD06izmlh1FWlSJO5Pwz5CIQ0QUPgC
Db75g6cxUfVvev0ZJ4IHj8GAK7iNVPHxr65rrL0XYVpCdECl/kwqQHxm0i9Yt37a3SlyjAHGkhse
aXXB3hwkPX9Ambx9Q3as5tWv8LtAMTVkEXHppUq6PEBkauoHO0Kafc9n6KzsUQSdrV3sQ5eYXsMD
1QtR2hLrQWe4f/xjwyysnatyiJcHeFP/Ml+Xkp+T3094J8wT5TzkhmRBU29ZSt147tXzpSI5JeS+
6mlBrAcZOkEeSPd9ZCgKD62aBnRhzgGp9LYlCrq3cq5qDZmDQBHGks3g+xy2hwj2E5iCzWak5Hqf
T8pT4iJEm0Y7c0mSyjeQMVxkSgDzomcGNpD3KZZCt9aTurgbLNt/yvu3n2o5n9f6U1Lp3g4URpoU
vmQngH/uXactZ032ws3DSkIBBvBdTmmp3je20VsYGV4cBfPo5l+RC6ydaw+NlFMEWolg7Th4365m
YZ9G1SC/NrzBIebFb4OOUqoz2/ClH4CdGNNEYkydv0oRBJlhXtCgR/zQtZ/5gqkxXEp+/uAD1Ynu
jNESb3yOXwZfjIYqHFsZIhqrka8kq0nhWhpaCo1ckP5frqNLPhIYH39Bm4koAxoxrywCGMRbyQXc
v4vlZfVhbpOD0e5gydrmTH2dYRuBM9hNZFxoaw1QpvMl7V5uMFJ/C91yXZ02Y8KsKayQPDfAt401
5V0hsVou2SHyoXIvAyjc+bS/bFuUFaxB2o91ZZK1gcB2INmTtK+T/EqXvevCxRQmLVYaw9tYIhxM
MzFstnTM02c9FUrp/kSBfosi4piwom8wJ/ojN3LBmDaxVwg2e4RwoCQ59MuYYZRUmyEdcU8gkQ6l
CZN21XAl/YqWIXt36spFT60q8v/q7pwY3WBL/aNmlLAXHPYcDFXDpdt4iom2xORwhdfeIhSRTlve
IHP/GIf84rWE6CYtBJHaOV0mhw1kQNVDGwOjLhKPPX912rUInqMw0QKm8wKFkQxNc2JGCLq8WoJ1
EkHD6RZJume4imFuMxQUnGu7d5Lx3GP3I8t5qiA4cKm7lnNAIpof7jHL9kKQ0uPSWesvPvS47IiF
UKNcSwELOjYCUpdzoQynADZ9hv8nh+kpYPMwGNbysw2vHA17rDIIJJER4Eu1GnhK78dBM36NRrmn
BOxEBTexwLpJwVeGjwRgG9Mjyts+aonXXnh+Bby2tXXq3grtTpJfaD4tVnxRiSMuhKnfZn9EW0AV
/qFZ3cGMs568iAEdO2uWXjAE4TylZ6+bVNMgJeC6EjHcnqRLBreH37funbWGPTpWE/WN2VvFFROL
YBnhRc2lHoUqUbIqYiAhLyA9IgAl2oglDLlpBOV94LcGzk4IVy3d/pSaBDCXFLdzf1JjRNnI2ClE
XVZPGABUfpgNRbCxwwnD+hwZNxTiyjTurqbJeU819d4bafDxs7YTX6mV0kmmXLYMIodUhEhWqpz7
/tajRV2fxUIAeQYNPH7Zd1v4ZRuKmnZXQChMZgbHz9vaGQwuC9kJvEzx28MJRwmcC0NavY0yVX+a
iBqW2sb+HQJO8F/bv0/7cg9hXBikPFB8HN4MQnQcWMU4yR4FnJTTwV1e03Bx5wKAembDvdkFSbor
jOooPPTtn/54/5pTwzk8+vV2yNp4xvaqkOSfGENMXce+Tr9JTz0jBk2sZr3erG/jPcEm8mDK/bNJ
0qU/YzHgdH8dTmuYa1cgCePsvTKMkL9SmvUJkRtERUteQSGztD3ASzDz235Gd7Miy6g0cYbKBudY
nzgtApiW8qY2nlo/JJVdkaEVzeP8VOopTeuDoDnYeiMzIxVDLrKh5njkg8T586kNjM4aeTw6xvYc
qfSTmRtFGHRRyD19S6ueIOPCwWHCn/ql0x9BGvtPOYUhMriFx/YQL5dCUHNtpbpKgKjMqSebFtV3
McpwNxoBq7++TKggV4TFP6p3Fq/vm4RXySg2S4fhXGbo3AmP8s/fQUUVZwItvYot0L5jEtdIiDJv
TVSPzejg9/wKgrhUHnPljfAcJny1ZFFECQCQVcMAg4EXr7lxNnq98uzcouVf/Pe2X8UBFClwwTML
hcl1GVi9a+FkO7W2RKc75ib5FU9TWtObjAdXW2qEC5ylvg8zeeXOKhdJpT82N1nrZHhGuJ8GjtuO
R8B0LP3r+3Ds0DTM7kz+Q/cn0fDl0ezPc7jRub2KCBK6TIZX2WdYsytnpAStzbbTlpMqH2SQPIZh
ixfit14z3d+WGhNDsHwOk+/9m6KnuHYogT2v0bKLJ+SV2zciyxF7XjPYdWGhqxE1Emq8x8tM57m0
M866AVqCbGed8to93nSC8GcLgxldlEw0/u0x8wDaSo84OBKUdBIrYyMdqkNL1TQBfoXn636XhPVD
+lbA9NNF2uyghZC9fEeGp/mGLB7ac4Z3pYASuCaBNWRJ16MHwzJXNSS+X3U2hqiEreVC5pqmGo+l
IgisbBBfEbkmoDdF5xr6QGAXbxK5ojTYW0Ig6xReasaszbm/V/V9EKaPE+4j/mqqy7/aXLFLv8dr
TiRbuOAvKvi13YfSDBSeiItA1NyPHL5nYmL44ZRsVRKLB2WA8/UU1hkmZ0WqdWxw08IifoYpgtZR
KOV4nB1L2p1t92BMsLkeX/wdazzl/5Hp4v1Pc65X/JpqAlpspfw8rOVYbwQi7scD9xD02bK+uc/I
10kFjm8Zq45jodmlnsJGg2PDaLISSN0HnHsSij5d0DP7FmlJo9CVgg00pp1VYGdxeSVPFolgpUtd
MUJVZSdxR56CDuN1FsVByffLylnI6cngkKXJ8HGYg5J3vreqehlN3z7VrtuCQIsTknMkweMz1Ueu
h7IClP2lAJUZ2jM3QeG3LGyxLeeDXvUtp8MoIo9rvU0hbU70/nIlhKuJVhz3AGAZfwKBM07blrkw
rZfDAwPadz1GPs9QSbnLqPkNELv/JQaWgsKlq7Y7O2USGF6xMvSbVToimB1OLRR37GiFAfDqzc4T
UuUXld3NT1WbOsaw3NZkdKR1JYC6r84Sl4ihqQn3crG2YtvN0AMPZ3w3snHfIZrG+GdCef8q8rsl
XguddS9ZHBW+BcxlCUrxTU82pH8V0EFFA+O0UkAUXUr4odUfu3GrPU7R6YvzUXMgR1M11R47IENI
tt7d3154XbxYZ9CKfyD8Xjdtk1cTvtRgZvDIi4AeK+lCjU9h7comuDqqLNUcwrbMrowHbOjojkAX
iJ8jygUhIZ7fzx9RKKXfWjuqunfFsF1zvxDlNR5CtzjrJxvlg9gG1EEc6xWK51kvh0t9j28QPWfM
nYEnw+s2vUR+i68YR2hSpIYcNvwqzdvPP4Fgibhqw2i1vxqNiPgYIIVxvsyw0YF6+bCyfZiQWzuH
xPad1dlUAnmD1gYrxBVKma+MVxTXQpgffHc7O3w5+Y9/oxXp59keuJn+pKDLIP09Oe6aUuS7ypM+
YCeFvXbJDd134Vg2+VJgwJ4OsfjfAKIkJcpdQNo06/HLaPPPQwsfS3Doxp3ExM9qveEm9Amw4BQ8
CFg9pEfQLjhE541Eb1KF50eeCq/qN74BDul/zEPWwUjkkxPh/Wi0v7Un1djgmhlcdvzvo50dYs3J
EFL2gp0qMEOxlaf142e0gAhdPVkZ7nAF/dVW9rmv/SdqeO6Q+bJxOLLTJPkwZyGOyGAQ/3/+6FqJ
rQPeOqezTOJoAhu1MgWlIUYV4+qJt4LF56fi6QVGkWpICZUXR93RB2K1DD2nD9miecAPWbCkas33
qw2RfuFDmMC6073D0Zl06J+kpl5zWaf2OByOyx8eJpoQ1XGmQLMRDh3vuIcr/tMvWYjtLQ3nm2/A
oftBPgYSU5djCdMZMk3UQB8yqzXWDiq+oq7j+G4VjdVQSssyCOgUFu3Nw/FJu+bY0mmGDfnF1MBC
3bP8LsQdpbSxg4wE0TQcuaPCMSEJlhiZFaRM3+S/wUC+JTGqhb4hozyFKxBd6wBuLXAjbaO4iGAy
4BcXbBoVRwjGgmPsOd3UnZmeWwxcbZ+g7sXPzmGrHNssD+RLzSTZAc3wZrH1wky9v0ywufDhhwnT
bhmuk2ikSD3DiDh9cffxwSkOlE8in6oM3gbFsf+d4znlTKf1iBWA0OiGKPVsVE/7yBbLoOxElsRw
k9JxOpQDawapIfwmAPM8fpsEHW8slM0AWAvMjurQ3YgAmnA/uYpVoWDNz27ROwXE8loTeSl6gKA1
yxcdtVAk6aong0d6gOQgSNaWX5hx08evqOLrRX/Zo3Bklha6wZfrzMLJY+EkYdqc9Z8UJwgDGbgH
oqHBtgkDHz+j5xKtHZx7UdBSaerx/CPsaIGBp8mVWIiMWoBNv6/EQXgkQyD0GOGitXqKoiNi7d8c
X7ftyMzIpklcVdygKTlzkl1631OPq2HHp9m0pL27H71MjTqR0N8OiAZqFbpRoLFGP5y7Y99+ijTi
E1yPqVZYNbzEWGPUHV7nMrf42CYPqtTsNLGUzZHYeWxmfy0ues4DxoY1tbPNh3LAQAmu9B5z64k/
4rgTxLmASgGD7lx4/LWzN1ApB8n7ZaF++Cgh4XmDYe2jyQcBbiLD3lcgFGPTNGYw16ISNoIu7jst
jiaJ0kk6/tbQuLBxlza4/jYcibYF4jecqy4FUSduh657mdqSw9GNW8e5DNAqUaay39svzWVujoRi
NmZH6ENe32SfuoPGgZa1hV240dxuI0UlDkslRa3Pearod/9Y3VMZUZti31B5tblhhj+sOLhFPs7y
ch/vVbjpC5bz62Z3ITVUKvU29HDUGjHvUxoosv3CYgEoWfhRtMd176HoShvK073HMGhMXcJT1hHh
HglsJVSnLxrhRpt08a7hihcc19ymwYH+QawMUqDVuzeHbzAzAzJgBhIJA/lnmYTfHZKQ7z4QIF5g
y/cdmuvVr8/eqlZ0/l+Au3OAcN96aetwUxwnDIT1mAkkI+iIcYmmHgWxRtEECkdbEscwzX7aeo0y
tR4IWvEo6XshAalWFibOjvz048Uwj+IYY2bzWAv5tptoLQF4ZKfRyiPiECzIzQR3oL3vn4b0ElON
x1UuwiOXxygrc88MFQ2FVP83M2KwSG9G86u0+Kd08TSslDziPnFx7ycyOMYYFMj1lYeFB8SEzA2q
KF9nY8Ke2iLSjNRI+JhxaxW58AgTvIFgNXsGSCsu6+MwrtHbQmK7FR7x351hYF2/jPap7yxs8Gip
hVyG4ebFO/p1/8i4fQ8U1NEkJfjJi5EHL3AeWxAu+b4PI3W+I08tAjnW4O2DEX+eVkkeBeADzm9u
A95AGPQxgv8C+cP6ErIkGmq/99jTyw3Do0FWi3fyIJ3a6Ivl0lEycc83zgC5DCigVc4P0Wxs/SEH
Mop9fX91W39JapPjPUv0zC8q4Nmi6+3/x3zfuZVI17mw96yA/UAk+27dlh6aKlzRC1xtvI/Vm/8v
kEaDAUMckfyscmaQz3O8iM48N/rPlSagn0k9JaS/NXvtHIiRpB9vzbR7o3Tm4GarKPqYjlhG79yV
MkgBVAw/WppU2w02PFNmViPZQYX4OEsMbxc+Ps670rUIu8he+ZR/drTofoeKdcQw/gUwE1EW8vPA
uYNEqEHp4mKV65basjagaVpY8fm1rvocY3SBqq0mtOMMOExhp1px7SGSi90tkXQJ1Jt2L6Oe4hjs
rZYvyYGX9lR4mku3b59Cad66ojfOxGvykV8TECQAZkCa08jR1Bq+Dfb2rwPPQTuodMFvheoiXl1a
nBTSw5Q4I2ZM+pXKCGxP94zb5dXd9ApQPDNnZY89JboMXnBFI4Ebf7eWRa8Eqw5XqvcNsE0tTTid
AsctQGvYLDsvnYBuc8CAaVvKR8TBOSlyu+3FhSJMvQRiIN0bapNkr/JVN9m2PpLyulAITTL55eWo
MXsp6oD+s40QOPma+Mfc15TetfA5tB0HFQaOHAMdLhX/Q0X7GEI6LRMMYemyJs9lt7pUVUlS6mAi
Fmm+tu3ogH/3jfwyyulaZlPFQ6HwYGxUHTCvgDgv2aR5s3RfJtupODsjrDBiKURtkIJ3+Yj8Ahbl
OGCG+RQYeayh1rCx5NKiyselyhB3jrTgl1dRBDdzNulC35M95SjCCC3jA4evmT8bOSREDdIXvhVE
M+Xm2tevgNeyKa5PKKLqgOtI/niaTMN4KwAVAimUFXnPcLfGRwey21t0/OOWqSHGhStFYDqIpuGC
BDZjaT8VttCYB1Ur716mlJURaSOzwDOVil2zT3b/m/JVyUlgXXyJ2uHL3vhPpmCcnVz7+xwiD8Mr
ACOt7c6QMe3KH4mq72pUx+LvEtarImHC5Oer8qjUFzji3Ig2SkUeryoBnDcHtO0FLg1BuvTNzHpX
tD4iilR8IXTyEC9fOmWfyDpqApZHd81pgggxxK+H7iPUgAbap0EugDmELXEM8M90naZ0r0LcoxFC
pysO33TRKM+vf0Nu1+S0ounruHxSGLMsuLNB2qMuYXMiAALNSTImX3P6jfV3aWc/8z69Ewk518ii
gREdSjh9bxbigXU+ZvLKmMhpw9wWfNcwuXFO0kiynfv7bpnRDnbxM05E64uDVDTeeuNqJHeWiH5x
kJ1cMygyC4b4w2V9GXnyWLMFcTWWqCr2tpK9AHoxg9DFZvya2y5gC6Dc5DJOk+nNdJ6K2+0+l8h+
1UhJyARhQ+V2c76lV9CMEMmayRP4NXzS/oHmSmK6JGmfrhG4khxmOoNnBEAfVRi2VN+vMTSAK8jE
jTB19dXJfEI0c1duqkgKUvf+Jqhl3SsDwwyklmCbgvEYllHHP8xQZcmO22cp/osrxo2l5Y2ak5M6
hNx0L/Xd5atdIfHpajWCqTwFTKjLZJk3FLgr0IAykHhlL3uHfdIowEOVX2dqWcvi6mDChw2STdwS
QgTRThc6J5Ju7KcS5lMNhRcXfnu0JBogmvnSQH+MLMfJldgjG9c/lTRc291MZL29GrWLLFrFyZtG
30Pqx6GQDdYufpH+083POubwVu+NsjQIBr0GYONP+Waf3bcz6k/vX8EybUWVRzLKjStNd6WsrnVq
P8dLBJJsYfbFMbOz/wkNnmsQZuOo9k953s/W5OIdcTHPYUrnWSTcI4X95eMuO7tKYEajhwmSy7DE
cLdn91WYIfi2s/Y75S/d6fJZCSCFsSu7e1EPyrnoWmositckxiqTHWO87IBQ3UNr0aI7H59z8qbU
H/N/aLduzvyAZqYXD7YEYQV3iHaU/Rhn5DIjpRkm01EThOgGEeaXhbRvpHluq5BEQ1OLfhlJNRzq
GQO1RwL7F5o95ucoghQQmkKUPbcUwBYRRGknjDqW3ADMb4wSjZT1xAiyMJiCm/zHqo8Xp1dFzVcP
oIr8xwydqONn3A6bOCyurSVUgHzphCTeYzJhP/bUZ6nd5HjzXDvTi/N4GpcbZCORG4cbdwo9lQQ+
Wb2KFg/XET1UQrr/iL5kL5/wWn5nRBuc/SKJklyde/KuJAfttBqd2y4KSLsOdn0rzoucBRJbKAYb
U3CxLQwusPnulE7RVjs2bBRAhJYQ5gcuw+tGuHE4EWofiSNhEr+9BaPeSb4HRIf/L18z4usX2BVT
sI1SuwkCisXU3L4+A1/N/UMC7/h/XE3/8Bi9HEWp/dgA0hbskp7dqa509x6ntu4s3gM6y4M5hOQ1
P6vUYuZxns9/dLv0GVgpAU7asY3+DVgyKq+h8nJEAX9mZIwoTPaKKU2Uc4cwIKEn0TEB34HytfJ1
+C6+fST1nw/44ruN9CUDA2cbZQADHYSIIck9Yp5FgH3cngTC31c7JarjUg5oNsu/7TYtzFbNIuYx
PguEjucZHgIO9PcNqXlX/DUtJBBTwyI4TKwNrGkrjBE/k4hK/LPggl+5bMYM3EQGDSyh95a3mG6O
BEGxxrKJXHGg2PugIqsfWucJGwuhFKMQ79SbP41WjzgjGh4zqYTV3ikF5+BVjUox/BOhu1lNtOg8
MG96n6e+o/3awHtV3YmfWDrHNPwO1oh0x9T6fNejSrjQpsS21APXTDwzHNfj0mkUpX0BZU1t5fau
MURhITQvV0vUYFkcCarupUxqYfaPPgRb0h4YqFS/6GPSG6XJ3l+4l8Q6vX4ZR6wy6krNDSXBTdSi
dpu/QFHSsFQQtnd2vNYt71KWQOE/koLAzoLtWntMAN78/7hLhhPhsTI4igCWopKmFLDt3V7LDpwd
xYZXBeBCdspH6qIdWZCUWB+8U6zgf1EMCM5hUYQQBS6NFA4rxbHNLQ5XxqRpYlqbdW7qK9ds+/ct
883Z05xIIOb6VsDPTU31RjAXZQkl+RCLVV52Ib/26t6wfxROjI+k476hR5B6F48KXPBccW59Hyho
65y8wFp4DEuiPDwxHrSWQ5BEsWW/OLpky1SQKRXxd9kT5Cm3Q7Zb8FwuGahGJjZnwyv0hRumGUVl
frxR4o4BDcmJftmdtScSS55yPeb1gKeYiEjlRQDDED7Etk8N8hRpEuK2+TkuNBKoZV6+4Gf3vZjV
rY/H06PEqYqFzFYrneLHqC8SPJq/kkvnk2gul+Lc9vVu0udzeumn2bhJi5f9opOPf1O0njrRrmBs
78TU96yMlFbuGC5cCSjmwvT2QjMq8nSw8kfZ3M7bwaK46ib440Cb04VHV+006vzZBeAvZyWF+62N
YRnzqs/CZ6NUVA+P34qN+rmQkr71IJRA7WTzADrZ6T4ej/4IHhIaev8n6F+DSakjGpoOdVaQzpG7
5Xm3eqxrV7O13sXrJRePjZU+ZYklmX32S9trQI+f49gsEWstNm38ILxFxmCFdp1cW6vydT845Uui
oSQkO9neG0KHfRNReAPL8yK/Kz0NHpA/hlGZHoY8WCiE0MJvqhd6vCUTfYBJemcVnlNqXwchjabb
zvCEL/fT7s3NE6vG2OQ0vDNIYkmQgsmf8z+Oo7FrSNbUuTm61ZXIQHilbIqsgdSi3lDvoGxe8+c8
o8a38ErWqKq45WppOhEBW1aek7c/8G7VDfTXP9W8NtCDGBkByRC2tt9mnvtsf/93K0PyzJDohptZ
4YGBeqvh9zKlJJ+ivdg9/2t6u5IOAUFQaJjitsLsHsoHv8Y8r8irnFglsnADftXRB+Tg/3awXvGj
0+29GSi2W1rRweyNnYaU3PjRARWM6ep+z2qRH3ar2PO0B16yTsQKze+N07rxvFhZMJxA1MROYUhs
4FPWNAZO9SEqka+NPh66fppPSh2bCxbSQv3L6rm9nTwNdh077A+TnLEPLFYeLPdgIiNCS6vj+/jx
iYTQyexoBHjZhfA8ydocusZ7cxXTxiqlO1bHRuf2tpchsEScKiKgLmYXYuPEivX3wEog7VOr0Px0
InY+rmxp862vAkDIqauYTrleQJYCDmNfTZAYaeSEsQsrjRurTg4vxEpo72Dx9UiNM6dNTo0G7nKZ
ZkOlHmwm8m24u1zVyKpOoluLaJq5BsIPPOqlUvtrgr3pNyDIgxmx+G8VUhhfkUm22YUCSY7Di7f9
rE6UvQz0n8bEa/ziyfXdVihy4B8B+mIOgQfskBXbPamid75D4I+gvJ4aMV0n/OlACc1lvqDH5kLg
1UKtcN0iLkawjPxVCOkZkQCJMaXkKfBr4w7v07Mhm+ZjjaGXY+M4+cxZ5q2YNE343iOd1doIKS4o
eEdFiKmcdFPR8JbMkfC2/jzR0SqryeH1ixxo7alVq7lWPnga5gJ/2riKGOHn7j1VFSTCVZUvFcCH
gnk7sTc0FTPbJ4I4f+OvOE3ZVJl3O/0X/+jTR+625eMxu3jkOoF+KQLdxRFs6FsD3F7LuxdNeg/Q
CJGfUKlvWKNLjoorbmb8uCxNAIJx1a7TJZlkaUfzcQ+SNZOoi7S80QhoWAR1K6RtKB06dbyPDSQx
J9TBbq0EqUGP0TX6p9vo1palOCmeJU0Ts1l72otTJGiYuBQAU04HBaxOyeDR51n4lcpUVYENP63C
s01QqUWTzKfWb51QavjmnoLqesYygHV9WTRE0InvHSWyqOV1pVahOKwBENjl/cG4lakwe6RJzUIj
SLcZHuuE7N1lN0EbiDiNnIuVdGrZdpVhkT9M1NvW51W/hBIMCS9YwITHXCqGzHWowY3T/o8RtmvL
17IQt5sj1cTywYGKXNfwIs5GMUfQOviGVugKjQkXc2bSxDmAzCVqfOS1eZFvGwOpIN6X63uFLqlE
hkQ/DAZIsYTic4QFmJLyv4plnjhiLIerfnEJyeYXWoKVtsEHyheKGGRGiIGvA7JSZX+z3dEvgPms
DqdYW//y0GTRnSNf2lnVOzqn+r4fTcWOR0L86LDs6GUOxkIn/hZ5a6ZU+6mQ8bJRFFCZhrp/RhKs
SyDvRmhvHDWGbg8ZyOFNpsaUZMngB2vDUR04elCa2NHHL/WHl5yH3sa5xbLrLrZT/hw0EwGm/BIm
LR0Xf9Yd9v5Je+7kBbY1ZP9DieB7j+BSFKqxMdmhTwLqJqi5cu6afEBnhBmjcNOd1ilWVxZk3sIZ
0/kDXQFmNeja1mjogEwUc2h2rbBTBrFKJZDkf4JW2wR7HF0CIfyrmiGoK6t+G6/hf7eX1UKrAfkS
Zq2G10vtwv5NDlhB89quZAqIdyYmRj7NxRsuMRORK+bfGRkDxQ4jly0j1T6Tu2oh6/992oFhx4ho
be3ORTuf/8zfwqnA4cdeHTTcd79dn53EzBN5OLfY2R4lT8tUVJFJn2MQSORbQAAdrFDzvxe+QwmN
YHxMXiPgpG9N0LS2tGx4fA0liBFNzZ8Fs/5h3y+zu7PtWI3t8r3S9v4kdBcRnLcFcX/0D0r24tKL
ekSjBo7Qt9UhDvLq5QbrdP2h/rkBQWYPOfiWyOpcQNkG0Lq0Eh5RHCgwruLlfgbT/+LGBAfYsAIC
Rms0e17hKRArvsepvWYItrX5jpHM3h90HJ1smz6nkDOcOI0GVyWRu97+2g5QaGlEwV2UGb42yXNs
5q4HwJ27+/XXZDT13nsUWfOyhXut15FQjc2G3ajdP971g38ITIWKaCb2j5YC1NVwldNycylu0Acy
zWAlpTxnpzj6wAIce3xlcseSBjZ7ajjk16dnvsl0vJTbXEj7zlH+ZAVHiKsml7xkGIVvEKBaOxh/
QHF2FMPAYCkBBsJFuk2BnN7f8obM4oHpTfhN2gnnm4KM9rJy19nSE9ed+SAY+zDlJY+/JLz+tvXs
QFmbPR2RCCIDu+CCqMIbHOR6aEBBF9sC5vOcs0dHttgmZOzmlB8M5/5KFekyGuhOOhkXEUbNLr8x
11ESwAofoGcVEU5UNRlYJDwc4WhZZjXJGZ6bPHz5sf+N8/gKcFB4w+msSv982MIWOO23j3MqSi1w
A9/xiR6SmzKhpMxdcdypIV6O5iVFF7c7To/NIHXEja0vI3s6VU1CocJSrWGeYQZLtFW8rFEATQeY
Ds6iZAo/Y6173fGt1PVhnx7UG72Nrhjzol4N7Nbsj8iBDxpQf1XpcL6vUaZEXhplQkugnRchYjAp
3ammhjz7v+QJg6dz+m151iRN31QwbMmOHk3tLqcmt0pio2dUzj7M+O1MXFtr2/2IIxlH5h9S9sS1
gVC/1Oabny0oO9bGf2mZYAlIiGQEw4ztvP5+jjka4AIkmXVYy4FkS+4RHFCTpJoKuuWaQuWnmM8z
1OOST/TqKyXBSmlg42exDaqGkG/22T0ouTux1KbVxwzrD71LSbbfGKlzpFg/sYTKD9M9/wHm0p0d
dttjy17DbgTak+YIWQ6wTU9oeVNSFBIRdpIJHOCBIg6wxhLF39LqLaNWj85HU99/SDt11aQM5X+0
qCH3rAk/xdRlc8HU6YrIAv0SPFn7I45QJRAYwGpfxufy6y5rq8BuQJqrPFkIN7jEQWdtW75KmOQy
u+W+XfOu6jERaJKPjJkx450NyBDkgLO67vDp52x33dxYYBxZzECsW4sRZPTMY2cnWyr7qodPk1aE
iyTSFEzXtKkGAQJ3XfF1f7GBRdSkgvNnSsEyIEUTlWX4IHK5VFojj7u6DoA2WQohvuxna6pfsnFm
w2revXAKHD6jtZ+YFwPsHe6mFsYA7OzZMliFjGnLcShDRVxbc1SRMdcOM340M2ddplUCCiTh1R5m
K+TvY/6y+RezZkcW14XWtH5JWkggCK2utnzP4JkWcZeB5y5FoE0j/XsN2p6acRBhf9nUCa9wXQ2f
e+nus3sumtOtqCfKkm75FQBGoWgPq97sBP/gJznGlBqEdB0WCOfCJ05GHBVJiykcA51Uw08lkwZa
TdytpdL5k8mnvCntltEIlEltvyugWGUr33DrOi2+Pns33OTD1Jw6MMHfVW1Eym+0KVm3qzdArsjN
cPT+EfJymkEwM8d9iYg1kyGDULeuyU/qkPfqctzfkOoNE6JLZZ8C7CmUjJvSuIyRdQRW9r7s5WQr
RRXDVtIm6e1kPblQQWhF8zj2YXeN+7/SbwtmhSZtIoffDdPFlj6+guPkBTZtdpbJR90EE+iGSPmz
M2LvZOcvgEOE7PLvkpUe+9M31KF8fx3HLmLKIDKni8oDVa1cpbdVwpSWD3H2tqMKI9qKDPOZJ6no
bUa3lSJII0+3Bshd+JJduEL7N34RouFJDlz7QhIKfHfHZBBLkgw1wTR94XyAahOqiTepFNi1pvTf
+MTuaRElEoFCT6QVm5Tv4PvV7qcyiE3OHiJB/tUUEMDYSLGtzdoBj5uvT6nMSPo+MjQPb0g1D8qP
HnYePyJCn8RPOn4OVZxJDX2lBfCYd3NWawtENh88jlYOi8rdmugQcp7OMQlgfw4i/pvu6Xi+tpwA
mUHk2QtyrLRo1s8fWKP+OeFG0mVB6RZ7Vs1giu/9e6nkXmX2BeuCicLf3s1UsYGOnhhQvjuTg5Aw
6IYGQ6Cy3OvMiNGOijf+Sb+oZ6povMAm3P9/FH38FqaErGjmoZEBUZdXzZp8MkZRNpebZtF1/f7H
slIBICpiW+K4wbvopQGYJKCGL4dtjnW/v0Iycl9+9iK7R3w82WoVoN63WJWSl0uXxmdctMWuUFUe
XORsIbGlbLr29ETQkfZ4sidaN3a0PMcJ8W6iLlXgMaZYiHKWDIxZZ+J16uX9n6KWfwFLhE8zF/x5
r8rWcWnvQStSahaS88sfeMj5IDTs1ZqvFVHBm+TVb71PFvaURnae8ISzSS0Vgh6Kbu6pUd9rsNCM
7GfTIOCfzFTjorYiR/ScwJnnrH+nvmKFNZvioA8Ji5qBnVgNhJvSvKMNr9adPmRcmq3W1tQw6ifp
TPPnBhpfoFhMw5OTW737E5DRR3PqXUsCcuBL/n6DO+lvEFpxb+55j/wJMbJmcw/BX2x5jJ65Q/xT
cNhQXIDnZeg/4X08+QQcUx9hEUwOk6D9lrxa8QPv2w4d1ic0HUJi4UZQHpkGNtDD+oC+BI2iHCLr
hSP0fipiEfNToRUN8gp3oaFpCSlWdY5kSdaJ4/GodU/oudEUzYFQY1V2qibmOfzvkHd2GiYBZsWk
tEpVnNpkBmsF0FL3mpQNEpgtDc+PlGEi0Vayh+29VNYC0CkXPzaxugIbs9wqbBGlHKsGa0KfozbM
NM2Aoz2mpVEhMduY5j0kCARvIoU4U6qYCwnxmUCpydMVY6/Q1JNjF+jB1IcJg2Ur6fQ+Kc/eu5bA
YjIerUuoqr7pFVjQrehvP4JUAM+RE4nWMFvDJEx7hpZSRKJhOdWieC2sP25MPDO3ost7XM6kEMu0
h9x2SKGZUPHSbbDaZ63I8CEtb1TbecEAgCF+oTtGDpDWzTI4dxyMhdoVel8StbC7jQ2tu+LtXWqq
pnCNrZl59NyM1cVNiohUByV3L3D1IG/nS4dv2C6X1oqJS8V5ySnkUBLS9LnIEPwH/55idMAwlPn+
/MWZYe5eZVrrNv1zY1vfp1k2WQyqizJYfOhyvmmGDs6bX3rpgt/vReVPXdGBSJEV4XjtSlEzRkVO
dGpMeZTh16TtxJnJVC1SB7Ci4A2Mt6ed1O6KaeQHfoab3RTSflqPoVYqOLFQt0JgNpo3b4r6cOdN
0qVZIM9Rf82D7oJJNJ3SQ3fIjW/1E7XGrlDY4OWNGsuXVotlsTL9w4xa8y7ZBHAkQMFkHh+/qD8Z
jxLVR/J8m3lhddbAQGhJ71Fl1yTamf8O4Gko0W3i/9BBKlFAOQ/5UzF11NriXfXs/rk9kBlCLZbS
FVVETVFWanF/NBMFn/WXG8mc74JXzwxQzEIZP9uKKGw61HnnnoZGduJeRhPmBha/9WFJ78mKKxb8
K8SFu4mneqY8nTHHZGHh51Hp68TKPM+2UKEICcfTR6sE6UfzVHz39iXc6FNSYVzx6C9z51bYY0WD
Wiuw3PQXalrIiw1VwHB6pgkdGzVNZbmqFMEMErFAaX1g9TNGzxGXvoIH1tPT2pH4hJSuxrSuUJE+
jH2ERBylCpcPZ6q8QSh5pMHPhYhY12AZ25K75pPmyHtLWcX/6k3isSDFR0C2wdzciewoMRoQOmAB
JIBwX3sEN5Z3ZorAbRAnspnYzHCv6L84kRmLyiyulQyzUlefRY7mnTd6mV+WLtIOEUG5fR1RlcUw
wUWIWDJ8HqlLAbnMRCWLPp6gojYDZ5RWV3CYmudmfGmD4C279RGXni3BpJLxB/noqwGKkp4j6+Kk
HofcvowGtD8BYeKx2UkreBKzmyEOwI+4ltdotY/CWwPP5trqGcokMqEVCFd61ZbZYXV04lTXN53Q
joZnsP8joJRGvgw0NfW/5xklmsrdnDDrMxtURivrkuay9O5ZRrQDifh9Fq8ZiakQwrEnfCyZktkj
KprmEdaBDZbv1JQD4bEAcblFkfAET3XeKj4SRPau3nonzI3OEk2a+CeXZiTnZCtXnzfzYjLs70dB
LpVQt6jVwDV6X4WF9oDXxdAYMcTtqF/3srVLt9JUTMjyH+3I209+XaLiOipf2XFKkv7DpgWR1nSS
JRd4oCmBbEk6ItKx8xLPQ0Vsg5Y79IMaZBpEREfdrnRAm9W57LCd5iMYqv4yGyub0pE3GjPwEF0+
uBizN2i3aR84Y2yqCSaKad1TWvYlb8TSzqbgtuXoQYfqy0Qys65H4z0Q05H7joaFU6b63x/VTjOw
sKidQnX6CUw19H0VBiSOjDxaYNNiGBIn6DMwfWdfH1UfATJAKngrSd2yaDOK6qYI49QAlL5bT61y
3KOCwfY30m1FIRKIlI9jS4MJFkmPq9BF8bfxRbBPwykx6z/tbHt44k4aoNCj7TBkYd8t2zPs9FSV
fbgvKY6Mph5rufe6P/WxsI/MVrXkPwrppS38LN8CqpEhAvseytkzwQ2nlleZJYqPWjqT91urB5ln
y1kH7ube1VMKzJ4JWwlTkXA8KrO7kUoPnkcPmmEA01CBcVsHrXFVV4piuj0socYlW2tsDZJml3As
qRuSTIPj3vxXPZ271lBY4Kq3QGRxYWVaNSueLJ19oWeuvA4fFMpY/Aifc196ZnMDLRhFLaWBK+Ny
lMZyG1eEWBTXIZmRFzOIx8sNNJXotsGWYglCsHMpMc9/mZXtmHKm5WQT/hbldQMBAoiwdu/CTV1N
egVaxiXryViOCbS91e54rOeCYEhNtvVbKG8rj4zGrl3fIE6YYa0vrNPFgjmgwX22d7nR0JUqd1fv
OaNFOn3f1GiDByuxF1ltJr/cY3QuVjuwQ+ZxzPeWZm3DQ0hqtLfqHb55H0sgAtQR1YhDQJJ7F09w
k6gXjtWmSA/bMJ7jOKIj3kiSC8pI2UVfU/oEXUyjw+WTp9ScPQRBAy1lBnm9NKpTr+eg4kVY10o5
B/aWfp83StD+ie8OBLUhPeD2aEpMT+I3q1Rra4SY1NIa8EzDbYucwJdiE87lvxMrPWpS1WMDw9im
9Fo/j7j5e4LVl0nDhgqENo6sRD+Q6/iPGw7vJ2zB2Sz1d1kGF+AVAJWzI4PfLMP7b/hGFUgmDDzX
5fu4ZP+b8CpuD5w6KIFz0/ZfPCTyDCxmTjvF8jcQHW7DVOwEqlhNvbM52kyYqHr2R7wo0Ma2ZHuS
Frt9G4ZSLy+dSJvp/a/9nAX2osNQ/hMW0gcwN7674ooUcwlXwrZoCP8NVrEzous71U51cTczjPQZ
pBr7xyqHrZ43048grlHX+m2nNwAPigQwu99n16TsRsEhIZpmjHJs4ZE35pVb3c1i/jgM1VgDk24+
AfKkrauRj/w6qCVYRuPbDyJbImynV7XNfsG8VjX3fqfvuDdUP/hp7nOAK80OVjSkMUd9MvDHiVfs
iuMBXLkCdrly0a1t7ZfqwfDRYA5KrnhY0Vy2QRwsexTNjPVhBMs7UiBGOV4bIKCHBwvV8juwW129
XEFa5zFlfKAW7cHAvzAd5K5+OkffU3yhIQRCx5zuqf5D3w7s4shmGk7UOcGPQgTF9ZBSgMxGpGGN
Jpt+kUDHK/6tBtSbMCP7wf5fNu/EyztIBiSkdB7q2SpC90TBlPuhlAdtJaEM9Wfb6ZNKpHx+Dl9c
AFUlt6tDWXhnbDFehM7j4SvqDRGJXe07qNHaGPXi5c3uvnce6iE3qI/RwWHu96DoJzdPy3Pg86NA
Yajfl9QGhtxKosr38qMrk1D8tBaCI4w2H3qu5LNk40nGLct45ERXXrxUswLllPpnHEY9IsDJdD34
UxbhizESA1SH/82jpm1zrXHmtC2DBR+okPohWKxIMlVCLL705vC6W0hfTTu5c0HA6MOZWDDKBrnX
zpVUQo/lpw2oekPCS60kuEo1S3k8lwiV/pjaH2ELt2imb6mqE5a81vQmiKb16r1EdLvPXdMaGEqU
juvloHkPp1QwMPjRszyr789E+Ou/BhX8yd1XFVZyWBkFuRlUk/v0Vz+2j7WvUVDFboEGfwRIWpU2
IvFot/QGyww0hPZuEORG4ywo/a0z/LdoGSIqolYskoXOBe25BMMf+nQZdzNn1QCETP6EhWIaWgTy
kx5EXepzYopIJF3BD8ZQYtLWccgZYnQnfeWpwzIZkbqKGEdTGfEq1a8fZcWM032aUHXvdg7YyHU9
8Fpd7KtjpPfllhp+sJNDP7iEJz+clnr5kvpiyGJiKEbhS7LZ2UAKf+Xu2EQz/2HfE+AYhL2T8GFX
n2GDHZGs2wfu0guQlm0Et12lGyuAJXt8s7oqboDSk9JlCHPLbiixEpy3pxX6UgWmnmd+eohM9die
kqI2LvgqlN5wHVx3TXGbwXx+nMNqtMDtRAjtiw/a9cnfiRZS4UZLAkboXuYdfshW934JuAvNNROy
c6ZD2RPfBsVyIiFwiblJlLJv0XsdZoRSS17leeHlXv4lZnxHhjfg9J1mBkFF7pUEZE1Wde3f2I89
y34erdzvvhbvXlSdmpHe2vwtRH2v7GQI+8UjeJtQnStX9BBKvshKEBZbkhrFDrxXiByTqguyi9Vk
5MSQunmBuprkz9EmNe+yf2jsVs8JsSfMyqdSdq+Eiv4orNcPhkwYEEO+Rf2UnNHrAIa5pvfCdrpB
x0sAEOIDBi3mViLHReqLkp0ge/l+oV4DW6+CFpCjgkLyH2kfOdC5jXePxR91QrDBtGTCG6+wOU3S
zQIntD39dZ6ROzQwhv2flP+B5vkqs6CCL27Nc+oxax1lacLxC8/c6Rkh43j23J5VeY4PyfUh/v5u
eb/2qRSvCCd6ReNmDitOy3CgsE69g/7gORs/LuUbqVuvjZ4UcnfnGAmv++cP7pWkJ3G3jH6HNOGM
oZ4keb0I99MHOwtbqZlaMXzkKtsbjEmmfqWvt6Wxy4BzYF/Dgb6uFw+vwCkdxhRbpqz2mbAtgwGh
YP5/jVKWFUb2HS7+p8AFRAy9GM0w/g/pj3BYMhRwWMYeVld9iPFlL3AUit5IIb5qLMB7yMBn/XVD
t+aHGGjSajn2kXPZqptAcXm5gWVSoUIoTg17KksSo0NKKQwmM7C2GvE/u0MtgG0uwcdiBkWfkRKX
Joq5XNpENfsWYehQw+pTrI5VKyhVnyJ/aBCLYjJ5srQ6HfTgNfX4NvLgIHTCnlocOTCxqK2Wr0ZY
xuHFBd5ze65YVKm9DKaaOYRpIeLMvMQ979loG0aYmGf2eqUmvKI0fSAc+Tz+vB0pc41eojjiqCbY
BVGGRXFUR/ii4NDmtXT0gpvRBobj6NO3k/IStjyWxbL88Uz7SiWncNu/ruw5is6eIN4ZNpjYVtDB
ElAArOp+LidEm36AXUqIIvncFYL7I7gM6Q7yBfHuTlquFJdpHQeV74zvryH3QEKQ8g/9tvuymH/2
FuLMuRlYzVY4AjJDkzmei0kLC+gs7QNcbXtn5CL8hopPi+KskkNYEMVoc31mptvG7AizGwklvOL+
6++SUlYGyj3kOUlZMPwIrrWumIq27gRxkWgoy1KetntvZZXA9+cJis/ovhU9PdV7Int+3JBaGw4W
iiLPjbKFAiW1v995ugzP6q/PtLh1GGx9T2XMDornGkTTSNoxeHgOtHiFYaoqHz34AIkPGwT22mae
psqh0UbtTj1yYkj5ZHta7ll+UGrg1dvEbTeIYjkDv0xRNsUTlGmGBBfYdeGJ2Cl7ClwXFg5ic5/2
GMNeD8aGUbBk/ykY5RxxIhIWifo7tBQja81neJh2AKhNv36vsP4jGXv7/nliAi89+bOuuYkpVUjU
jhaoF6BLH5HDb/NQCndYzDMBo4obd2XDgzViVHEUIafCMMp6VpJ4ST6drkuxHAdw9h+utpZ8qZeh
ty1t7YQPqkCPzyiIU5D2/Gpm+hZioPSAZxTNOUS9jHBrTz+bIRhLaRzqiWiu2CcnHvbtJrVVMTKh
k0ZzLaoKvWjWoFNyD+h4wW5gapmivpq3tZEZFHTAAp6RdiVyT7A5yD03pZTyB8WZbfMK8+ikbKyZ
KXozx1NG+zDWNkA2hQD8kqEpaEfW5rQS+t6oNjMKRCBsf+85kvJnGJX4tLoYxBK1qZi/wmUnTVrk
VlakPI2/U/4x2IGw6Rp4kt2MJc+DfR8nYHVf+i906Vjrjj1LdWgdWy7vAHiU5C84MCT4ww4D93Zq
bkJoBMUzPpnisFKO1PZdi0KkrYRInjaO2UTrNmsCsTaBLObEcMBQ0WDmXr4cSyuyxeR9n9j3z/bp
YDfDo5tlrfDa0nVdgKtigrOqIcH6bnZ4i4q6lHfAB6CQHJs7uir8C9VUwMxBZWCc7emc9sq3aSGN
q++6GyCvJfmFQvf1hChYHuWayS80AwL4w7rIqXhw6BzddwMIVPctRmhi3sCDymyxNTXbIJ0CkeiY
laKNQtymIE2sboaxWynT7Hmzm4w6ulfCwp5FQXDDMyXASdvJtBPxqZSjZy+7mnHP6DrgrbaSKfFQ
F8NfZlFNOSvs4YKE1TmWc52j1Mrc+aZV9Wp28RCcQxxhmHy1PXx9fEYUSqpu0Yt4aUetCpyeEjoP
E+BuwmvHt30tOVkat7wgV3TUAviI9XVapc3ofkCJY6OPVvV+zvRH8EyFQIWsuD3ocqNaQ8hB60qr
ttPwqGzwJsY/UWaVTa8NavprPzvCzXDKMNkpknMz+w2z9PUKVTS+YM0bj3NHU1aSMt/IRoRnbZds
QXnfl0vDI0wOT4eXMResTDVFBePsHbOTvC1utM8uiI+BtmgLRA9zSQyVjTR4a0jSflSRfKJyo1C1
peM6iylFK+uuugyoTO+BNAPE83LOiCURNaRtcgmnCFgA59YGCtWk9I4f1BcWiZBnuz+tiRfWAbfx
gDSm38ITP2cnSFfT2CX/2qEZqTHmUB/r3m4Q3lLw7IGqXdK+N2yftw948rXLBp/kfU+s+cl6FtZP
WlmZ7sfyswMcF/5ov2HxWhBx1jW8BQuTyvepBJpybClNtqL+wi4q4I7APqnM3MjA8t7KGfyX0ys3
wmch6DDgiFLDgYmsf99M5fUEj/EaUHeVn1POkL8HnAGVz6JRoCZiej+3BA6vvtIg+xBTuasxH2d1
0Ha94zuNYR1z6errxb/Ake9ZaVYeQChch0u7bHuZF1ak1dvbIYVhNUBkhLVuZsRFPFkRpV0jy0Mz
uHzXvIASoF+Q98YsaVZmKo5ZPKtKOhM5TWERi9CZExunbhGC5TYhtHKQmZNAwGuifUDmTYn5tWQS
44Zz7CFYT2Z57wdTI42vUTfKCYBxHt/dGlbzD71mLYm9/KHfEXA+WKwIjMsT6/xtlrPrFC9RtKnj
dFcdtQBDu7zerOD96NisJpp/a4/l3WKskwd3o9Z2yLejDuPD3kzQ4qxFIrpCIFP3g79+InAyBjfV
9TMGRZhcFpBweixGGJ69KAVciHmntFw1zKifp1srFjT38NSgpaooHWQ8rQ27Le/NZ4n8HMyHpHZ9
MYDK4CcjH6pHpDyoaVdONUcl3htWRqYGDaHKTYWgimZH0DKLTcA1P1suKJs5VeEckCpG3sUVU3EC
XUD9GMluolqP5XSZ6sX1jm4nawlR5cNdZi2LZempt8nPwUFLDSzxHftglnaAyoFPaPLnoqLjkdev
AnlUtHrqtu8aoPybQiviIf0N4+flLNe8IScEWKd8prynt4m4jKPtZwB8v2AhaTha1BmkWrKqBmF0
qKYfk00hZFg6JrBEpbumecNeD7+eoV5deVmfsKuX8FipRlrE2yNcl2UjyPPYqvzLLF1fg+M6Mquy
QLZyBaTRUl6c0P5+NuUPIfp/WmbFDTax0OCWSy/v7KfZhYiypZ9jF40CsKq4YlYq3anXmWsypyCD
Q+NixTLAk0PrX+Mm+oFHwvGhlrnYdPZOZ6HujBL+soh8t5ghgVUc1zEoG/u+avWwECq9+ugyLegX
GQQM556GokmzZ6ST+ddfLELHC52IbYNORnnvZASFOyFn7kjs8Fge4FFE1FkGOci60zKApRrb8Orv
+Vr5pt7ZLDG34s4Xi8mnugWa35HPuB+BPDw528/BLU9/EuaM8XUOyzhcl7VsXRPpNIp9UJHjkUMq
nWGekeqvrWXhv645uTGQ3glssRXtxjW2huMYMfP0xEHy90kzS5KormgHApR4NeV/BVCPiECw3VkN
gTMCrYRNx1umc1kFlNcayIV/07SOcjBMoJm4kHDkj1I+dzvBDI/rAjyIX3UjGiH/wBMulXUPUFmp
fIONq6AlOmw2nQ8TtHsRIe5i4pXgjx7SXTGVYHr3kEKtF4QNNqtdn9cp7c3zYmsRT95aAiwNB/7X
4hbk/9zMoxIgAOe6K0E8sBSbXMx2Bk6bt21ctbDNOdVIjqoJpl7ycEPqGrAciWNFzzBBWRikemg7
ffGUHxUbP++DOWkJ9Tx3L70EI3XmYl9cW+P3fXSGLF1v83YYXJ8krDQLlWdPnKSCJPjVUy8nB3Ul
wDw+dEh3k1NnXajf5SuPjrOY+nBOllkrIbdRWO1Pvvc4kRl40S7yqbQbzVVewOnF7WpY1Wp8LgVx
1tTW/4RPEYndZZo1oigKNL0rU8GvA0l1uMD4b74GizLgJZaaBvltfSzwKgw2uqyAepLgR+oYTOd9
npA1+tdieMCBAtCJ1EQRra/fL0/nCcC/RCjCMZ/Y4bgGUnbnl8T6osm4cA9eP0HAQi828r8BlaGC
XipvEIHee0pfqBscEV8FCyCl+Bd0RfJlqGAAmS5v4uQnGXnuHHzq6UTHJVYNg6g1n8TAqS3Crrue
YLT9P3ZcxXj2ZR/jjhHbAMIsp0Wq6uPT626HjOMFyJ3goGTPV6YfBQ9GCsn4CWMS7IDwWxOVl31t
QehCwvazomnb6Q8NtIkw/PJ9AIVSBMOW1IBHejisZ5+bQbaTwIg8ovxQ+Zl/xpHlrWj+DSyDGkVZ
5wd4kfVB/dy0ObS2YwVgwoRcTA7cCyOmYb2k+1IDMeTSotYlo+Y0UFqGuypJ3gHOhR/MQQvuN5nq
annAgLswpKN7oic9qTwQ6bv+gbxS/i0brGy2Yvn3UJr55LWxBjwFqQIsJ9G/Oc9oK1ymfyabMrOR
LNEj8pTXeLVDTpFjjhzox/IwU8zve8vFMPkEg/HgQotW3ihcW5vsaFPvQIbAnAcrNqjJSHFDbEY+
Rm5hS5y6SBJhryTSoybLg7WreIS0LptfVBGy0a1w4eG4xA6JqZLEW3ZfzC3XdCegsd/CeHMGFqfH
qY4fAuRJIUzPZxtirllPMS/pLhF6Y8q/1J4NAvhTRWQUhFiE9mZlnKYigkUhisBLRz3p+j6bN0cr
DJKZ/q49qtyRF19mMA7+/c2i3YKOs7j4GZbWTotdBRSXSOZWpXlLhOfoj1fFrl94hDORYiOvTZrV
trS0s6M0h9oj8uLl31CcQJ9jjxlOK4Ne8amFGupW5GptHI6X9qfjY2s/8mOTd+Cmz77lIghg5I+Y
PHJnQ/NRdLFE9ouZAWJb2PP7L7LUS0d/9cgfjLgh4hzHMcrhxIMW+4ocmDsp9t6kF/zfEW+y92mB
O8otY5M+Dt6Kvgd1z2WIMtdnSFg/o22c6nUIv2jRu836nwGwcI+sdo27SHFAFc2RsTE4N1VjEUO9
e4OUFQqA5FpFe6decPSHFOufoRtQdrAOGsktnFafPk9mtQpfmSSn1DVNW+cyUVu8ttgGk2SwTpjs
kAGsYxCJS+UkMTMk8sKDfz6W6a9ECD/GTv9Tg6CKQq+Zwn/3O3aSH0VrU+L3AXkKoOuwjYDqLD1i
Imxja+8Jxfl2y4Ua33EbhCS0ENQLbnq7mavCbj/vjwmYt0Fe6CaXDQw9gBFDN8avHZAK8dI7VF4K
PyNK+gojpvDHjmfXZn6RAC9EMmPeYBN2UZGzJrv6mfqArU/XfGE3gfGbjZwxaj6QsJ6eU3LexCde
usvHxNSkoH6MrlhdUwI6X/pTUZm8fQxOUh8avn3lKrZ36UsjrhHydhvXiheg+gAiEz1yCu9PMrsl
LBvT5yQbnWJlCnsfWqGcHlascnqWu11MnoO88rAnwRpaPy0KytcMJSYeXaTRjnfc9svv3hhFdEbA
Hi2n1/mc10jM4DzBm2ovzsCRQbTs1bee4pOA3hjYCqqPa802gPpV4L5G6Bx5Tcz9XuEYr+GepAbq
2qNqeDyxwUPI2CXHojwbd7/NAv0JlbiKkPhi7Q0jynS9oSf5FV2SWxGg0oTs9tBWg8iKOBCwK5+X
U9Iil8/3VbyFYKkNL3nckeXB7sqTOaeyYYAXctEjU6habFWm7NFhFtJ7y/e54urCOvIUukeUiSiG
rh4yJkeghH9ZeQj8ZQBilATAbROshXWYpHYJevYtv1gpg71EEXi2mLHnO5iS7k1fEzT70FhytVq3
s713a3/UhGeH286/Dm7kJES6K6rWuv9DWsTWpraEcrQZRJBJLscxwT6U5I5DhZIX8g9ZTujXigSd
XXIyAeu2yIFKNjBTttfvhq+ThQCaF9KD8c4gSJz+B5UmgjMnRfXEaDqi0m3QflDErgD8+p5G0i/E
j0SpTPrmBTR3OCdwbfbBY8Uc0a4o9b1EBUhuiugx8IGlNeO3uSkBbcVbsPFAcQxioQ2rvlJEzwIy
0TQcQN4TwXZM87XhSKg31niDtY1WSFd7uWVglti73JJyJ6RegkygFFuAe1fWN6pSvT2d5kIiVuf/
VlMq9DOJ2L5leU5cTs+iwOwXadB5newLilqLGSaDrACjSTdZzZ+ByEyKSaZt99y2GB2jxdjbVAEH
1SFvTHKRq6+0ccDcpDKIAhaTp3JZEbfkIgu/e3tIOZX40q7IJryoYS2MrcsP2kGK89y/RpbgX+Ok
0VuKfL5q3tajBR3n67vwiVbR6Q0Xx6KUh6ApnhIPZgLv/rxTbp2MQAf1p82meqbFbJ+PAKO9ALgn
If9ffKtBxAVcooBtfk4yGbG5xsoZ6Rwk3LkF8550UTXnQkdZE/SwPPT60LQJH2KO1SbI5g6bYfrB
zrudz5bKP0Qprhhu2B182EwEc4Sdf/hvHMd8n26n/MRBl06pp+EZIrd06DPYYR+GtxfzNLnTi61J
TwwwJi6DSyZbY3zffcyk64mIFD9cwqrwO59pl2pjs5INOWrTQyaBIAEWKlOmM6ZRurvkjr3Z79r2
wYmJT672TiN+tnSPBvRi1eAyQVAU5nTaHN9nhRAkugWxyIaYfT1yX6/djvENsw2e3Jl1nhYNuogs
RoBUqXaPZLkZlNi36kjCTZiEaQzSJnDKicS2ZQoMpaU+oZ2kMv6F+qH6YQpUzmZJoKJh6W6Ir/0L
Lawb+RLDdZ2mUP0mmPN8IC2vW3ktB7QidfzQ7CvdsXHEipQLePz0PeKwZNyx74dzxsBmgI5yRBc7
XtdYvOG5NYxUPwgPx8WvafB8qkSHSaRWm67nwNexYHzEmS1KgA4hvTu0XNmWYryTBL+7N4GIf9t5
jskuQhTN7lAcVqxGPwd+W1HJ3aqGjX7X/Wf/Lpfnx7peOl8ms9hybvHOMfsRCudN8N7G80ApOx0a
P/dfzVFfYPpYcbvUlxvRWdYWiyiRpJLUUht0zUnpXkbrWatqqfhqDnlTAxnoo+2GFXzpzbKwu0Bo
0gna82UiBzMj2Fu4zCh48zPRS3FG8spsYH1fnW0XAntW0sjn1Bc8QtmMT5V3e90rmt7BsNNianj8
ZI4YmcaPzdgCHQlZSOX/78Hu7U6ivVnx9SANuENasNqZTAqpPyOSd188WHcLwaIkdnDavMqf+Kur
3XIg6iAWzAO1dOlVthIQYZR41ZkQCfbLJMsvVNSeVpIerYJnk4OO7zYez+eE+zyXFN1UFzFt6CkG
2fE30/I756799ERenxMnw/ojc8XJoJnzZYIn+rnfkaxIy3NfPzkZaUJuq4SeIF6BUPLmbrzEcWKk
nnBBOheblQBJ4WzEzdZOJq6ZkKBjWlLiKIlzE//ihYWOlTZToKWBVngcFTjVUI7P4JsY+SmZW3ed
+hSHzw5Zwz7rmdk1I6qCiJpr9EeHSzhSKY64A9fLoS/+Yeg5I/NzRurlxqpYgLmycfBea33nnb4Z
jCvo81u++eiNmIXaSN5cx9Fhc4n+bTeAyIW0vlhVQ8YFKQlQRY9OXscoMBhbsgzag/5D6xI1aAzj
fth3O9jHnE1zzFKgAeycZKSXJOehzM+VJpX7/h5gT+UXc5MMKbhrtyKtgUu2TRQ82vLDaLyx4Pxx
CAAmfOAjgSk7OjVT+3+NoENKiIKqV4mawONscMjUHFJRXk3cqI0lz8pWO66GPRZLckwA3cnyxzXA
rYOKPkCuIUZCHJ15V4H4Z+WzmOhhv/ciu/qXZMx77UGAvVAZar47tGrwAYBO0+KOJMDPEytPBQVp
xAjwze8MOZbC9ANRM+iiuufp0wlkZ/zakHtZZp6IDrOrmoczuPizKfsW8WDEz5d4daKfg5H5Yb+Y
jITkJGisILr3+k9kLEyhlhpODNSHcUF7bIXYJKhgYwn1EtgdC3/MkL+2Hf2ub6MROE1GKXiH3WIG
NEqCylIus21BguII31FYA0HBk/oATkFPfK902JjqBnY9fr8VRcQbEIyHJNRodfD5KTutmb3J1JOe
BlEMC638kF5IHAshtpdn6N8fxjx3YJ4oViogsD47FHpIYhD9FUTkFDIcv0QGq3ILkpcfylgxP+it
s84sl05lrZJASryNZUZ0MzMrwr4jkOSu2BJ6ZTtheodYbEMMJZ0214HYOn5R88or34uQpcuMYvIO
TioLJKqzlFKpTZwWKxOzRdli2AMMhT62oPWNhSB0w3Eg3QiHNtQyDGD2PBQrG5o/3RYMByMLvhrT
QqdLwQJOZBLlWzi41f4mutetswkUPTu8XLi2Bv1qzn2vHcT1FGYedtoT3N2dy91K/TChLiC1/ZSi
DnLDH4TFNJiaeOMrFbhfZfBleiCpRj7gu42VN/koRYlaVzDta8gbljJ5HTlbwPhluCK+KxEFJRZE
Z+HvYob+MKUrU1Etqywi0WHHyM5tQeDJQku62JaW6rU2pqAfpUKMfjGnHYit2a4P6/4lU8G1qfwy
EkRsq59ZRbrR0kX34HPWaZQsPD/7f8490pmYs1Ly4zBGZD17z90G9XKfH9TmmEAC/Eolaj77FauQ
qjPOYwzpIihDAPvI9Jz1w+bsRYOTnfGNZCD/btA+vy0V8GzixsXy69RnilV4OTYTDzD/4ZjVv5VX
WdDUJB8kZwLLCEpLonUI3s1GftrpC/+r5AoBK3ovXaKlEvhaIKB5zgzc/pTaGLKGR5yHCwoAFDge
1JV1+yDMU62D+AB5IWnjC55kfpzefy5c1WEiW16peakny5e+BIc/TTr9T1N2TDgiuPhMZuJuGBeo
NO4VqJWPq1RD7+5kWTPh6sFJbzrQeFQgRpHyLuIp5VGI3ZBpBDCEQAnz6YYhsWJE07AdgnuTPEvU
3iF4p9TdS3nRPjuovm4QgmGvCnQAoYdBbLpD7dzXVitQQvtYLC+SPGePhtD7zGmMdrfIaclRxBw6
MBwbUTLde+P/JKazDGEpmjOJxq9zdbm0qI5m6VOMgrXoBv58cou0AolKjRFLuOpvIDb9kmZGM+K9
0FqJ376poPn2WlTPmM9jiaD5odDGskI2Tlu9fWoUGA7Tefke2W3wuPWeOqsIqEvGeb1u8I09R5HZ
AITRcSoYKo0yzX9tNRLFSIq+b3jbAZX4X6P7zM8U1FCAnSNQwhhY3lwGA+dap5FF2iNnNf67f6cz
gMYk8QlIG5ZrypD82+G0ZqHGbpcRhgcMnLY38Rdwg5Jc0ws1+Nxlx5aVUVVIzLr344IVdGKlU+Hy
6vhFvLjwGJqtv+OxFyLTmsMfZ180Wx3IfvzUSE2qCrDHk2VVQoPP63pEm1oe7ep3EkRF9KUIp3D4
es5c1bnVUWoO7vZP90U5CaQMJivOzBSoWTzCgvW1ct2amO4cvNDfkggTzAy4NPqW7GU1zr8K938h
RAAtI57z+IzJ4FtxnT1EV4UygW1wC9mJIqTx42MZEPNwwAa7eFo8FWODjwSr/D/DYzph0VuA6DKG
Sk3mRG62q5//e/EDeJFipoPEQr2ESsNSxncU8YHRAuTDXc4HuwkxZFSaFOam/pSo0+ve23G98E1N
CBvWwO/lt7NkUU14jj6wf5g/3nuB813KBXoBTDcQyNKF2FtZk84Ualo5+I6ihjFaTteMwTd1LN4e
2RzDfKixYNXMnZBt+2cu6kuTKd+eTiFij7mTtPCGlztD1GvUS1pBXtzo6teNgAUhUnYbvmLvDFPW
O5QHnQO3AiXTsshHpZOuPzPAm0r2ctut8LR9Hvcpwr2m9qKC5T/+vNiD6rscqQkrD9ICQ1RdzPAE
Obh8DuwIJHVgMAuFJdNq9no6ftlRg9z1W7lN1z2gRCRJRDUsGLvxjKbO/sWKHmJNxEAxwYtKw20f
aOSyQpQWw3YgS0uQ+/zLATCUhIYmr+ib4ZzJI39Pl8buPWUMQ43EsQJUO8NTUJ6aOrbBWxMAtWSt
Fu67X/kaCtKDXnu1eqzuKuXLfdW3JFe533BJWJk1+y5EMFGNyBom9aZdNWRHMZytg33UCzxLD1al
ezqJiXCuhYqnd78UHlAX2JbLiOdyiuf3RVQNl0bghUfakAk040clgw7H/6uBpHAWT5GhADxd1SkW
WliWysdA+GydEIJM1yOJ1Jp79kufZm8+BdsR/ahAers1jnk1OlQ/CeX3C8RUl3EkF46bb79iDO/f
h5QN4A2anRZNn/9aC+PuMYsrMC5JndWJ58MKzyLs6rHf6nTwNe4YZdn3dkuZRjYVIJUfZcOVOOc2
2g0VYabTBFhySWL12pL9/pKhLtwiMMQhZzoeAhOvWPQ9bd0JZea2h7YNY0boCQTHBvAuD++qshaA
OSmSgcJkP2ddCvv3/KeKjNlftwJb2obwaqSxRGswoEsoWunfjzJ8Eg1ZE8SVvsBcWWgRusPiE/zA
x0WQ0qBFYByunkATzlV+MGAK9S3mQ9PYfSyTGusRykLNsOZVSVNgVOyGr+DGy9fcHvpj/ZVf0dl1
p2xqBiRiE0CIcWiTDVdFD1qjY6qFN5TJM7BFaQ0QY5a/JgGbn/6+7PE8p8JEmFtY4JW9SyyKFXZu
TFe8Cw/Ky8DC0geRqM+ifWornaLaKAuazZkl+5XlSQwzSmLTflv9qmPnS457McCe4gVHV7elT1hO
au55yH+B4qA65oWDBe6rIppdqQdy2DkqxJLJ9T4i/EqFvhuuY0sP1z2V7CviEhvVnWD/NoEgwfds
YM51Pk77bFzyjN9X6E2AbZ8Bhbl5gG6WkYw8xzEBsegTkVbKBg6prCiyhUqXklaY2weVji7ihgpl
9LD6wp0fozVqOdhHR4vwxpi7vk7h4Ui0uez0Ohom1aon5h1kGmFRiaFdmdtKGQlYPxnAul3RF04l
4vb2IQgXpK4FlzGoXe9zgX0MxtYg6heS5xND4oHO75ge6pu4n1XQcbmnBKd82k8z7mvPsg4KVOHk
BHnC90b5vi13/rH6SrlL4ykf6Z9z4tGKNn+DPaFyEFF1kB5GublWyuSphcnnoiEiB0WPQv4Lgbl2
gRag/pIhB5Vw4GIa6biZtssg0/vS8OFch3rEpJyfNMVx1tPy38Ubz3KlUXfQZqZi2fflY/ihpJjW
MlPuxF2ZFipHRTDJnxSypXVzcr+ERhcL2733yRj/Tt9wL4XK5LiCcIrKnRG7jDNLGKDAJRJXGV69
vAVi5r9k6j/Qq0kBktrAg9BR2MkFJc0tyCBo/65IKMvrjHaxmV7za0nQrgLVJd/+lR7l4qhosTyb
OAivoenvxHHLg2k2FEEIozlhByb1YleugWo19ZOjCRpGikIYnnyP9Nw/LmFjLM0O6++glBWhCxDC
DE17l/PGWju/r6ynzy7WlLy1kgz/sc/gXcdhrNpe9ZCpS/J5oEkQfOVkjVbe/C900ZD92iEm3Aoi
o+gb+da1T/WFRtOC1YNcPb2NQmPSDplx0CWjCb9aiS6ImBWJLEvB7in8/ey31MXCDApx1i4u0vSJ
Y5mFvDCDjz4SVwS9dqmHCqDjZ0oq7Bf3Pv18HwwXtSGYUQdrtgfKVGcNb4IdUV2VkKbz7+PeOVfQ
MKlAC2+KweTuiCwVKSHJYHi+tKGpG0qRVJDh9BsPFYhu5PMZqHSrPuSWGIX0RG3+IySwAFsXAZFP
HgK0xsDIJxrEBz63HnqpM/7C5Xd8fnzCk8k8O9AM8cbW5GJa7uRBJrruIvSNZ0QP+q4ioNTST78G
xieh0txqkmnfRSzpjTj281JKkizs3tYKXIdjSH0CFRaWtwW+7J7SkE1ZvKiPSqwWrdGddNuwhSd2
faFjGjJHihA4IwpMdYP3bafIZDJlkTKIG3vXIV62QnwukbOUECND7qZZYlXKQZaB/BlTC2iNoBlm
cbsu2fLy1XeUqGzapwMRV7VzVH+HHLg5Lkxof1zsCgtjh7HaepAuIJDvzEUwA4WmNPqGuSUHcV73
K3kwxS6nujC2+fEPq6T9p1VBLXWKPEXQ52APm/1ohI9Y0PQXNHgrT+rZqkcW/wYNnzJbpf1uIBZp
ASvp6yACY786kEiLExjJyKGFACzEUDyO2ZvvQNUzquv+5ru86Q+0y0gcbaAU2fg5J195OcHWP2wB
VXMgPaiPx8pT2nHuIA6GdYbPCyJkNHrxcUDoDD2zVop8JTRaiNVhGS1RYjOCmubSVLa2/pti/hfz
9Pv6exW6rBbH0x8t07Jb+3FZDP+DA/rYcw/DSq2zGnRF2w0Rtg+NIfso3MYIRYpIEMiVx13tTDyf
g6NSAltIJVJXf86cxZ/nud7Cs5zjz1undZOCzDqBLpStQ/p/RqC/PVPU91+FcbaGBwQ1unoU2l9h
DmbWQ+7guAVLmcW9QmV1SjrxUjRX8uCZ2WsempPQpKepqPdQebWKxt8SNi6w/CiH9MWB9pbkhDSw
2hFaGhTpxIEXeZ+9REwQumtpl6QqufR44dmxmpxaBnLh2EtmGSrb/HHUAxEmnEaephdqccfOxcuR
C2edgliWCAdJ+PkYdv6Lp+77hSJXZC5b2SZY5ELYnglwA0CScxBT3cV2hYnGzaqxqOZvY3CZwszB
lPACNkwxf4oEwarAc6vDFkYbZTW32uy7GBtcdKWGsf6Qu1QqcI1xk0tvCGuxY6K9jiUhhRQtysPU
4QFJnP2LAmrZQzxKprIdlBcXNxRDJK9UAiWD6JZo168NMc1gTwrFdFMaMFSTuaY0TRWLCWk/FsLB
esmKE32l+sYuKpCAGK3XMw/Q8OcbSx33F2HQIi0hwixdia9CFijuypTF2GoGDMRanNez057z4MQ5
GPQtwUzyl14NtjPqKsNJNjVD6+bX95SxKwAbZRvQf3CChR0DtVqhpP2FscC/+9uTVLzwvTagayGO
Tw1vSnuKY/qEUYxBNW0QZP0GVIJPxogJPA+FY+NCqHa+ed4xl6Sobn5T5pNqowY7YpnOZhY8j/cy
DPfziKgI00fzk/jEmshFXhLNaDd3uNI/4o20du2kM/P55h/u/D7Dv7b0+nDRHEGg6RQBX27f++Gh
IMJuIfQ9+1tzSv/o3MkaDegU5z8yHpRP0ihq8PMEUe0wTn7AOUk69BCpdd/pTaml+J04KxvM4uGq
dK+lHC8pZfGBLVBUQZdZ0o7Q5xv277lFjd3JnZtwdjeg14TbAldvB34+MykaHfz6ccPYOQ7U3Gj6
gahern63EqYmo/MwmvF/4VDzBM1jWK5AgjhA3Y0hCLk8IboK8UcUjM9Mnf5VHQxA0xZLzT1mGiz+
RNzTNNgoyZz6CgkZ34D3yf0fsuj4QqRBACBtevkibPdz5JlyIQ8tZheliRobB7RzapIBIMk1u1p4
f3y6Foav/Mxv29L+cIcPie0bTxfJawNcpkLmb/YdZTuRvq8szF8OGfNZJn6DW2BNZbeRLcaryn4s
m+nosHGGul1WKXLyMIlBjFSBEK8dTUR1Ja7EfFlA8csURLsDlxt9jnD4UiQEK9csM7iVTzHvpfyC
UhyD0JJriOnHZv3MdsUwSdfi4bQHqZP3WQUiDdyoiQp7B888Nk56N2Q7fSuBIw/qqqX51x2iOFQn
jMSFQAoX7JcvsSXhdkNKcSYLJ3eAZz9oz5zfHielDJSNZBiHQ/X4Bzy9/cU/EaLy9wfgNxz13U+4
0eEMSU2M+9p6cH7KKoHKG6kjl3z6z/VFLhDvAvQNOYd8RufUmzrYJTXYKooOjyfK9ikPp4I1xq5g
DQZmO51pO5+qSor47U5Zku8UxqO6kqbnXoa0JywvIMRBiHmO7RgxJnw69+cCtaw08Tng6o31t8dg
OavUaE+sy6gU9y76IvB2ULJxa5+pFkoi1ORZGYDgbSOk3k+ttDE403koJ/5y3jJXt1WYfdVZAIGI
jqeIbT1Va8FeDEM7QT5ZPjbjaCa9eXykIoLOS7Z8s4beaIb3wCy2GD4Abw7yniyMj8hmMTkqsfi+
vVR+XOAN2WgxBkilgpZc7QUouMGushyzv8KHGTGRbxDYIBPF/LZSjwYsbTiYqIle8moegOpDo5eC
E/NsX8hlM2VjttbyDor+rEuC5/EZLHh7Ct7Ep7YxNIKGMtkftisSRiZ4TxS+8sS1m1O8y9hN4GP5
695+pYSZtKX80gzEeoj2SymK1aDT4x4aNA5hOP5RcXE/fHeRdz7AxNGRI+mTZFl6GAtxQUB0o5/9
F3jRmNTjEjUK+e0UmvYE600RycbWo0AZeS35+HWxLeZv0nU8O98/r8bd4FJdZNOSHSU4wcGLmtwD
sJxEXurPFEnQJDymi0Y/JzSn2wmXgzN8SVVrpQWKZgbkLICmZeA9PFu5RmTsOMH8fCYQ/umN7nCB
u9qxvaoLR4aSE19yJ1lRrMlD6RpmHeHoDraRPLtCoUyXIr+4gbjR44hAFAzGg5aAFo6/zu00emyD
RIiZRkSYUWfYxhBFImP0zDUilcywlS7j6uci9VuO4h7ep/ZF0nzqP3vN/hj0nD+lCApwwCxVREGc
18i6K2She0rHICIocHd/i+c+rTjvx/vsRge1VzDZsBO6YPfx8cFX/t3tgmD7XZq3lk0vF8vmE9s1
Ob0ddmYSyO+J5T3OIuf7R0fG4cjA+Y52ft+6SiAy+nEIMbVYGDhXUWVPCmX7vNV0olGtgP9by1RX
RoZa/uDTRCvBf6l2gBqZBTxNckZSoSh9M7EqTnGEp1uuV6seXpOmvTMhPDgvhdbP87Mf3oVt6Of4
uSRL6+LgGwih5nf48ZeO4Cg7TfoUn2PpXq+/B0fznJ7CZxtnnSwhn4nLTtbWAjAfl0Myl35QmZZr
PBA8riu+BKBWiQamA/wwnY+xg0E/5yUSwni0093TkEIAppYLUZmMCIPfmRrdCQEp1ma9FJqZTU9k
nrw2k/N2q8T6YYT95hcgf/5U1xDCRqs5q7iQZBi3eSwKyrsv2I5/jcspBZGiBtuXzx1/ukYCuZax
JVQiE42yZXAMPqjwOjSuFKZEVYjcWmPO+SKlneWsWd6/TDsJRIuaSEA7ZwUP1D2UWfbwblMlStIg
o5xAkOoicVheJAhf6CfJd6s8raadzOibF05P+2DJjVnPfKSAcgMyGSAP6suLi045GkV+I6R849xh
jdvc2gsK9jr/cIcVZksVwefE5HtEs/aV5Rt/+JULJsWN5vKBw4VMaWEvj+1QNyjhjC+nJovgletI
ltcsWUZAbFAnGv1qi3/XSHvRqTMi9lK8FLCJJEreTIBskQBLjlnKNFXJ3aQDZvOcWbqGW1/3qLc9
RSBmcvt5zwFccuoFfh9nAxdkQbXoslpGgEwTfBRftWyvM29WluJLf71LD/ummxrMOilvim3XlAHJ
C0Y8xr8aYoZW/kSGWFINWEB6iis6MLrKi2EiLKJovELnl6mTZCnWkAcb/WkSSYlefTMRuDyWWr91
gZZzTTbD+cdg1XZ5k2OBh6VDFdd72wu9ZOEbiUtf1OCvTiRK6Mmpq+0jhm2V75qA0MTPD8zgALoR
pPicVBthc/1Qrfj7ZiFyCUzJjgFyWWpEkViO2+MslOTcoHlNjSyAmnT2PGBv6h9STwZGOHcUfCFK
6BpJLp9uCJ/q67GzUjmiVVw1ke5o2OYyIv3MIdv7qnpbeLBXcJ9sezg4KLugmfVmuPTR+W/rBVEg
Ai9ZJc0HlBlfh3EYeni+iqbdNMSFF2SxWk/mdomjHPXbM5RApouBndsPjaXmkyds/fnvIOcmCsT+
CimtEwEladmNQkjf0/hBAeQQZEe/Yp1H0X6cLmJbLJLsdRrSsijE6WKvjug7mK4U7p4f4a/ajobS
gYUYiAJ7dXfOCdOaSiJfsaLssm17ztDiwsX6uPH2oaJy3+3lvq4hZbHYFrsyoY8O7Lo1SPrM9BER
c1XCha4asF+dPlBe5Meim7I2zB/i0nVSxF2IzdYwG3mxtkFoGnuO7PUyuj37iOPdUzyVC0j1LybU
0pdqlR7s/FPFaWoFV+oFXJZroe3NO5cHqimQqj+JERr3uq1mkXwPAQi/UE/HwygD3rnzJzneIQnb
RxbHhRxSfYjX1POCzirZa3yNUuXNxJY87zcH5l/w+w57NS+/j2Oa1QmgXssvLiSjA6d/gGdwMBqX
VppM01GbmekAaT5aZ8rNTh1FG0XgeLW9Jzoxc5uZo9DiPu26fOxvaJqAN42CIBVqsweqiuHvFO3k
06QWc2nK1S5/YJpTugMNWaVe640v8kBkcCugYPW42YYP3dGQ5KOj/NVUDAWruGLcaQSg05fsI5VV
i/QkEyEabtGUm8OBTukSZbo9PFzFeUrIHIiqEDH6LKZCvwQkL7HfAutSpkDAMHKIOp9F1p51eQk0
lmnhYG5otv0Z19Zj15YNvvvOHK5YHJ7KCkPAQcmbT7ITpir4C/u58vNFm1d25TeEvAHJKkxJX1Jm
pQ5FfNTsW9S+2Yz6132jSaSLjCmHpJjweadDq7HDwjY4cw7/jGp3jYS9BSiMZZigmfaOuBOi0ADf
I/N2uJb+2GVcf1ew92WbR3WX0bED1CJm8IcpCe+vq/7+GCOADzGgwgAyO626S7my7FSe7D9L7mLN
e5XyT+AFwh7C7A7WhValKQk26yi8qK1eHNT4O7Wr7hNmQrqstQPFdzloPVgGEJrhLVH28lQN3SKD
JObHJnwULm4VHsranmxSKk9Xy/VwSxfe/FBMjc+cPPz0AggJG1ojWjYl9nOGsWvyjj57x378wOMf
cZhPx63QQovtYIkAXvKzXfvncvm2b6jTG/jDtPHWbW3ENj7ZmKKL+XuuHCdSfdcO8TMwnExuD7IN
6wS+BlXymdi4Ao54cfiYGTxPIC1XOQwyHyfluaCzTRy63NGYerKCFQvFWinkbGOtNYSRfCw+dLj0
jjBG+LZI5pi0I8Unu8UARVGQHQn+63qFtGXDUPg69oMCzit7fx7XWCo0fuwbBLRK7LetacAdHcSu
iQB6vSqP6H0tGhqzhQzD0kJua91opyPfS9CYEs49Xduin4rynMHEDsmE/0mwMVaQUhdvp7qjni9/
uY+SpS2zOv8W95jDSnbslVT1HvLplK8E9y5seawcwg4mr8r31A0nZSV3E936/mKMlCvaQwDyakHY
Yp57o5w+SSMZ0/eKFs9/oeNy6BRtbc3yGe4iTe0E93kvLgGgwMVzZ/tvplHCemgu1yzrKGgsYPON
eJMu5NY3EDiX6XMfjURGCXeS8ONiCeoLKk7v2LphrN5Vf2L77dnyN57q7y4SRGGVJpVMmaKo0wzO
hDvaXHKTCDdwI1UyXfRNunYMxEodSy+FWkdMtV2mvasmUBH6q5sFE0gCVRnUbKXKz5O05DJn7vIU
aPRgNPbveAnVCjyWgYOGSml6bJNc5vuiEkq4MZ0Y4G7XAaS++682o+7cReuLUof5A1JfFpKaRqQU
zt3mM5A5NPK48EJu9iKpRa9g2rb5XqAdtHIb4jOTJd88stac+ddiuXbSaYTbFIrqvfGm52eqwuha
7M8ap/Pd7n4/T/L9O1oROqlT06DZaryQf7wRVF4TZc57eE1q1m/3WpD6SCn3tNu3HgP85DpqLTyc
6AfA3ozfwVDYNi3cjRa4vjcrEGKCtRCt+W9AgYJEgUIzqa2Q19ql9oA1G3GmbGSgDZ8cFr68OWIT
/bbusnGmOemjDurTa0xxFig3dwu/LBMENF7GE2sr2SPaaqI5kfz7CkaQCWjznw3TF50bce2vDATa
A1dJKHHYkufHwpzaoTaQrf+/Z5haz07nRE2ITinqRN8HOZ/BcmLdWRZQRtr+sRJatgDv/czGTcVq
sci+h/bd79+y60rV3o2TK3tJJKVdl2WZVyoFWc2QMPyzhPYiZvvx1soI/OuhQMWngBPwf083vSfz
Wkeih5MLOvdDIrVuFpfJORYfzNaacmX4+4nru9VWzKO90ADD6jZhvOu+SJ0+b0X1ObslfDQ93VAu
M35bq8NrFBDAekXvSDI9Xt/qrSwLvX6yF3bAccNFfBGvnTkvvrnyz3EcQ/6SW9j2rsltxthavwy2
s1NNXEPtt1wcmyErgJx7vjFts17SsfyyXfnwdD2eag0xqHAu+8PVDO9/oWh3sCrjV4Tat12X15/S
alhheEA+ZOV8OvT1C47V+SAFrHJuNSRjTxDM6iLkm33Rqtzc0rVcbDvTnJ77b26gNJOgv+W3SxAA
l5hdLb7Huc95MKcwkzKonydtevH4EL1fXRySY2jggyYA1cVSUd0RnKAtZ5LgJ97xViigwtpQLurt
CGhlnAk1VqUatNPBKYaH/eFI/KLJcym++9r4hNrxYGyN1ahpPcqQEoIWlHWVF+5GmOhN2OtWY+VS
L55iGkS05eC8/v2T2bAkhScAXEeaVU5cjSRtoP7BQhOnESpTeT95D1SP7duePQQ4JIPEeWVob4lD
fSpbUZq1FomA3ytGBTisVJWkYmaOPv24pPegFjMB8XG2MecwjVs4TvzBiWk8M7A984aYaUpzq9cI
BTU2XOrSaMjxCA96FhyTHbOy9fckdXgABHNB/c6pBzIPR9hD2uqKWlbsmVWEEXCKmHJxyuwD73A2
c1S2AS3esavf27ogmZLLFI4WCfO4pso97nNgjnVS4h86tDdMyA6O4q1DzthKwMPQCWhk19MTsN1M
AFDCdsOBB8cOMeIf0jJbdsJjX3bMDRwmqo7RNi8yPHJgm3lVqk3yJRfDOxWJ5PSasOPLfOH1b1Tq
zSlqIMye8UvDse6jAMmKLXWew67D2JDFMrD49cev+W20oFC67KGIrIyJIDnH4mFSd1cQzkMb97N2
hWpbDuhrvc6AyQrM/t9m/Rq9Jc8eJdPn5rQ8UFZtaOtopaFUd8pM0d8yHc7uk3mWBwPF0+5l9o5q
YiZkgDqay6QOkvHt8HCtwkhNQVMc+nsExzlYfxoLDw+EGEjI4FByJtQSZYeWPDRAEYmpVSaOm8yt
Wy/RUzM+fCHD6RUeBDDElW9gaqwAPbhtB4WKnE/Ma8b472rqkeEesRHExADlTUDtEx7dkVpmV8df
Jo5ZLaNsjpL8XL1Zrj21fPoWQH7P4IVU1u1LC+Xwwn7EsvnA2dTTYPFgOvbfPp1PBJPs753WBZXU
rQ6BBBZswxyeR6G7vcGkJ2R2bAZU/jOF1JBfo0i2QLPAZM096GM9f4xR1X0fQmiEibIbAozQ8CRm
SopNu1hw8zHQgvLCoauKzXK9JYEZaqpR1KyzgbSo2AL1QxPrJ3A1mG0EolHEY+iervLWwcEzvXY7
Pajl4AH9L3gTrZEVMayvZhe3xPimlNb6KGNPBaE7Plt5el+naTOZU6f7MG53Et6nxBROPh61cucu
6iAe495/DLZh3K1Rp0sb183ubnNZIBXXfDbWD6KqNoQCdcJP5iryGqaO8BBll3oJ1idw8+4blo1q
LA71VWn+9dCDUxWHuaxNJsclljKaTb5cF3isLnzrmpdau0UDj1HfPxUgMh7VdnagDx7er8utQeL4
4tO+Az1RzSUYquRdRWLcpFLQZAcoF973jzlz/8cVAcd8vb8nMCBGLGECrre8JQwrqMlsVYJiV9Dq
DBlsT9bjigysOvPooJaJlRpTkF4mEUTCkc3+xCBjG8D5c571hDH/wpGpb9riYq5fRPjXEFinD0Tz
T3SPtN4abRHWQ6OvbsJPVZZD/HE8+h5BVmNoGcxZgM3Q16wWNJH7GY3TvRLFcfot8oW5ICmZANNr
BwO+TiACxuXCfO0+kCQykY7vTFACVRwjvW/G7VksOwBtQvEyqGTMQHh7adbUiFCBCQak6kZJ6OfT
jj2M3/9jY28VzIFIOEZ5kcnbyEDe9yZ0k5pNBqQdCD89ivgarX1BLgvoOYCJkTgvBh9ujs5ujqvW
kUZJNPBYrozdjZBFyAX/tdITCWxEey54kC6XTntIiJbavnzTsh+NDeFx+yoNj/foq+PngBrtht+R
DPerISYXqTxdV9sn9MawrZTGnEi+6XMHnR4ASx+wZiizLS/MG/usWa6ieD1ePIS0fgeGxn2isZCi
CjXFlBsS0OZtKC6bD+9wdVy086+WhvRkVG4J5rIA1EXOzOa1VhuwF66bTBo5PAkd+DtSjLGhzU9A
Ja+09U9hhCfk1/lytsIRIK3xB1LcLpbdn0hegfLgV5gz7/iniI/oq8+qDhax/D302pxds2T029in
U3dLdg7RWa65oARFPqrbotehake8O0DQR447/japkiFSMG4Q2Akk4qBb4+kr27FmRffP7SYsAwQN
qo2dAFkYAZqfhCBeZbQ4KxdeHK6k7GWFce7iaPaALC2ka7PfhH94RQL/IAK6bKx32AaZL+SwEZhm
/JgG7B4AsTT655t1HSNvaQlwdrWB5DHR4Wr/N05be1nTsXg/WoZ7opjrF3XiHwJZmHQtT8+c40q9
F7K1b+Adwqhwh4zGqsIV1lo1ZBlA3l0NMRwt0SNtOwwiLULlI6yd+7Tm0KiJ0SJ62Y63YoLjlBSK
EOI9AON+xK+qlsfh9g7HzqQnehHat/0FRORSwL038c6m+6+xKPCqfNgjM7vhgANkH87vEjKlLChj
ALeCI7BJZQofOr1PWeERI3+hy+YnTR+iUvr6J/HURmKxw2H5FpvU/ThvTnlEpinT9gSJ1wZ0O8Aa
cdn+RTLpcAih/LDyZcsx29LkB297EcDaUukpZmSQfNK+s0cQZWs62AREYa3FBnFs+MkXN5tGHRLl
nq7cVFZWD/uJ3FIxaNJDXzt70vydEsa40c2KhF0TN5NoJZOMQUVjmRDEW9gJH9DG5iDG6wMKR+zp
UzSwukk/jlfbf/W+Y/zDIIKpI8CUZnXCr4qU44rwgjHYTEIDnY6gKyHlcY6pOS1ap5XXaf/vBSIG
H64i3+IrSPjbNUVMCjdyZqRcwhXBzgHg9gqzwkXfTSuOuGbSU2aljzwmaFJ03+dYxH1jDCJcAy3x
aRut1U/yZvv+t5x0oWYR2hBYrQ6sH2vxT6dlfAeT3et/jbGFW8tGOMf8Jy9jzyHx9dShL4Ue0I+P
HAEiAtdHwLEgNRAzeH+r04xrChDML38zz9IYLZBnh3ThILrDf0svEgiVW7nvcxGaXHaBhNpXgzl8
GF9ElbCGHgi9iuLBB5DkPmVIVLpS8kcaEOkmVrL67tksTGYVg4q0ovkXrsOuJSH173W1QRPkZ5dn
FVRFxJ/Rao5GSAhrujEiK/rmehYQFuHjht3hf68wkqkdgya9EZXDDxzoKoleXlWLwjIGEUGQ0LdK
iCtP7zCgB5oNgthITR00f0nEpFMgMrmFhrmYqOH3pcIXYq7YrPJCkyVWOyFvgs9ATbLYmW2/grcT
iBQDtvnQAlubC7DkJR7IGcOO8GCsGwSDZR1blZuJBZd7Z3clwLKNqJ48O7Wk6zqVJRmTa3AMuom9
zJL/YMeg71pIRnYQKumz+8OPCrYOsG1tY6CJM7tpwKfAVW0lBbbPs8Rz+XIuRdI4sIePs/7mzbzT
2s/FmnYHyNmUhQ3csKP9A40YpHjDN3RQqfJE2Xtrb4NNBRKVwCENMEVlUTl3o2JD78WwdXi8LKzW
tdJKdoVLZ2/NU2xb7VqpDTeztZzgTmXvKfDll/3xXDa5+NtIX7ixKXuCig6zvO5cq4U85OdmBCYJ
3UFWt7TY3V4MZvWdEuffLK+qCOCz9dAAucSbzq9X7NIrCayyuRLoGCc2ySaGobPgNcf+Rqh+jTxO
S1zn0Kw+2kKScLpJndl0aaTNoo6sEmo2luFLeYCqjd7vs+LNXcOPDxGHA46c9LRVy0qVgcMZPdSP
luCUXHlIU9HSLW5jlhneDKj8P/nP0lztPaW6XzM90nahFJSO+9P5wF6wYUlDkecjM2k9pIzM1uJm
IvTxjNp/R0bo7wXvfsVL0LqKJbOA1zlFCm4jfpzFDn0OnkU0JjA+lJfKvcv0JlGh29phvaNyWz20
SVt5ZcsCvUK6FfYok3zPvkk83QBR+fPvNg/zRe84PDEl5phNuDnVbaqZKrs7MTIPE04aJeQEn3rt
3XuxTDVKhKOTERa3XT9OaVPzuSOhhyD5SgCadXZVXlSueMpsd7ID78KI6abKvaF/afprGAkcA74U
65ekMX9p3/02Xov3cHbR5/2QmMVtxJ/VoJ01WLOYD+n56X86/2ziJihljqNEdyHUf6TkGNm5AqN+
5d1rA3CCC4556iWvmZKwpHlOF9lG5u2eRZE1CfXyMcZACRX6vwXMTJ3Uyjw1te+eNpOYzgxWmfzs
DPzzWyuXa7IIVtYNyLfBZm6Kgkc/xbl9wcvbTFMk9w5kJXOfGCz46CokDGixdX0SRRgRWfzBMoeP
ijuLmQZCPSv2mizgKqB4j99Zqb9C/kWmBwgTuH2vUDh/Hm5HP+B/yrkGvPWweY9zuFIWVYEV3tcA
QyEZdiiVHgwnvf4F5RExQ0ZQZCW4p6k5eXp7wAKg2hbKW190OJ1P8Yby1yA+HAZ4UPoXJ+IP8eGW
CZfqimCoQ68aEinnMIbDtqrE3oPJS3b3yR4kgaDg0sEIF20e8EITUTNN0gK2BO6ly/szzkFvUWC6
SdNCihUSxfN42MLVdgyofVOZwL/sPAhVQexnJPnDNtEE8K3gSBiXvoRVt8K9rA/yFAGue74oDNg3
DdT0gKNTPK5wN98q2YvGTZsHPxDrdz0Gr1WLB7mA/wBqqBLwlo3mYOPz1P4nFC/Kxwj7C1EbxJTv
YjMunoQGveq4NV3w0pfQoMPS1MFhhcSiBzkYiANSyHUlFutRSeGN7y1pg26tcIAkwTFcnhfzxYdh
duKUnX/B3tcY3TNBbciKmUkWrfl2U0ESEZ2kl3UM7uxo+JwGyhvKtRL9JP+DunviXabtvjrQuwFW
EIyw8hREO5qmUcgJJ6aYlhDKydb26i5bIR9iCix178xiQWPregRQLbx3pS6Qq5L7yDP+vGYD9Wb/
ZPVp88JyAaHOtWtuWHdwVrlrUgm0CUdtmY3ONcNVkZyZctt8mEV/BhPpSwOucgfKfBSjdCJ798zU
SvTVHBoWKvXlmYjvrCgmn4DIFSPXX8zgG5fwyxfAfCYYLM2W9hQHRFp+aVdGhwT9WhyKgyFu2h53
diouZwOhPIm7ri+OFPy6ik9bBc80gY5lysIA91NYlh9oIxS1LAEfGjlUeUDBfVRYDVMXjBkAcEmR
86AubLYrLfKV4UsAHfgrel4OkkGiTF6+P/syoFNQub14OmTSxehXo4K5KBQQUn78zyGZqZAY7ahg
JoJy3ha85hK2RRanfLroY/JXqB/5+k9P3IpeDFkEgQFTcz8IDIeYFiowUO/ixMPDvmVb7X6tic9Y
g3ry+2dJMujVGdMAuzhl3VS+1hUQ0O72/0RXWNEGcceSLVkGoMdyFMOCgtCF46iDndTfW4MYmJ+t
059nz6C7mpUz8RWl3HYrmnPeNh8niCW/TYolEYAAn/33dZWEuoXhNVmjgA2qZ2cYqu9xyhDTwcw3
6ENVoTPeemDMxSnJng6eGvmkiI8zfyjQmwyccuLPRVOl6qQPKoOrMnKWHgtSGKzO0zqShLX72wMl
X4tmWE6U7WLaWWxTJvdLVbIWiJhDZHaHpGW6YlSAyzEuJkH5RJVQEWjVonJyVwbQ24ibWZ20IdmK
0HPtua4+4mdHM5Qo1/ybSoakdF09NNvZlckwsIRxkjqRLoFCyUgox+QsoyzxZx2R63YrF5Pq93HU
FX9ebiGMF7ghFNQ5t20aOS+bwVsjCRlDTx3cUyhuOHlIOcWoEr2ODGr+InVNtMm9QpSORZzRrz5l
uK7n8LGoBgPvl3PragAzbS5D3bCDo2SE/nOAKEtCd1zkiA/B8o9TgzQD/N/8B4FR+51YkC1Z6Nmv
9sobvH/GQFsJqxIpJ6jUFGR9RjhS6DKKfNY9VaLn78mzDtHUx/DIY+KH01HX3t6nOMCVvMxPck+m
MslCog6GCc1B+xj01klh3S9CpnxRcQcLQCbBJ//bwXFndXCr897NaJcQ1HhlSe3KutaheSMrEEwv
hIZR0jDf/4ktTd3b1yAnSh113x+KFjgYnixoMAyVlwTia2bZx4zAXDr9p+jUziwfSsK5A6VLRCEf
ns06T5WALJQ36PIT0cWJ4e2KDlxqyX1cZjtlz9qMghs7UIxvQ7ZAt4CpcTlBgFCGbiVuUo873wOd
+g/X7yd0wOy0A0uA1eFcSBM+TMhtLou4lbTIlj5r/71HloXS08IutHHpjdETxcBS2psPFTAcQdUO
3vHp8QGVjvh4RR7R9q0urquLEfknokhbaG/0kq0YiCMuvWYkw4BgMUYP8BzbOmRLbgOGoqiDH8JG
s/sHPWpX6igoNIAFDWKR1kNKLWgN+iY/Dd3Gq8VRBGEKRQbYavfRz1nXmkkM/3ZREGUGHL8e5YA7
QThWAWhlsBjCs+EApVWO+8KvTcOt/W3kkUaOEK+ChkD1b3RaGo5px56QAT2p7MNaX02XczapBCJR
qongvWZ8dtxFzCYilmtYX6pjjMw6tiVwTcBsVrDDMz2etAMtDgQ4HZB9Y0TmrgSdFCkdVY161heE
hIiuXhNy06MogOvBha8YTvOC/kl7v6qABiAhZdvCDTL2PESAGeZM8zRGKkTGnyjZSljsig+0q33t
BGwCo9H7tEEQNkE1qzz14ObF6r166sVZ9U+nQ+kfXrS8y7jUVUJNqfB0YNNHMNB2yb6qN4f9D+j9
HICIXxd7gtHCETIh0JSM9QewZkewd53hjOz4snI80kHUzsGyMl0+HjV8WfJ1GJ4JQb+cyYu8AJ+1
XmQ4XQLfWTVvFob23njK51bB60fGuZLDJ2uspZaiuv2QHwxbxMIVHKt6SqJhjfKTZVkk9yowZFoX
fvjjDVzzPefUlestGF9wQR/zAjfF2q7Jew0S0/BmJQ6UDITPxZTdnosVFUM9nhw5aNAj2JUY0AcV
FICBiTy+pv6eWbq/1BuYCsS2tF/tQpaU1iWuGJcPumbdaYDlT0b/rmwz2xpCMRrvnoJgDOJCbgVA
YC3Y9vud+dbAKi2NhzK67litOk9079x7LX3MVta3mkVzBT+04OHA0LmhEyjlV4EQ32QTtiTaj/3/
Ls+q8hRcMKhrn+Vcy4vv8bs8itXOvwGv7GlE+6f3aZUrRDyR/pHXm8HbxekA6OH/tQe85kEB/92R
dTCEOPipW5HFIYoxITUMt14xGEnSUcPwSKduUC9RwE+/3WtBczgR7uClRcB3ZW15AsCAS6D1DLrO
N3iIHeE0BCVtEqpfl/Yu+8B4gZXeiWOIsCAeSFeszPKkgnJGePYsrdchFl6l8p6Z6tIte9wqRW+a
Nx4BRIHQCKQI14P8VlFGY2EZudIAAld2G88lIyI9bRWS/+t53aTTJpFV38KJxHrZRWg1Yf6P+EVp
bPGOfvaghOICyTgk0TZyRCO5B12FlKJAYOBMNWBBHtmrQGWYuWHgTT5T1NVFs77iTOPihevtUYjB
xrYuXDz9VT8iJs5UCZOEY+O1URiKOK71eL+FKvCYP3+Hck5kWugjOIs7saXAf1SatfZmw5Z8zc0B
qm290pevEXyF4ISTaY21dzDWbUvlMytmgcMNIUASVFLZlXKohAvOTdO+UgTopR/nJOqx/T3LZlFj
Sh1R5mYOOri/ZQq2GqJY2pfQc8dsMqh2e9j5MV1HsUw4cgo1BqbZtHjpNbcgr14g/tS4syg+59BX
Z3TIk772qEF/x3OUES+LLml7cC93j//1HRFNMdBCiY3EtIMtbr7hi+68CqvwJqbmxwjroyXiCvw3
QQJhfUbrEMK76nnDwbWPG1beFoAFvH1rLPg2EEP0yzvf+SUrFoRSvPONtTMs4KQSs/icLv7KJn97
OL9TEU7wZVdU/DXWcYcz5pEEHm/cxlO2aRpN3Cn/t5lS667HtBV4y/tDkMlzyeQfOXd8eLpTYgpk
8M9Gn4IIU6nvEuPmSSNBlVKmrOrdAohmtFSxhXi70mRe4B+XNcsEokR/lCO9WCOxB405iIYCNwim
Q44pM4Bxm2B9ag7ZRhXuS/yrQHkLPmwNkcwCOhDxZljbRTNbxsKiphfPkC33mPR7RFn9ytzWnMZo
CArf8NLPZbf2GFXt6d/dRVtK6C4sCKGkKJVm8PtgESJ0N9RW5ASJ+50z3nEXOcK5+8RvblVNUcoo
1GhZUFa6DevidqPY8gx6vqPH9KRrHAt6FtfxzmrsjYbVC0PrOG2epxtFyxIV4+oEgiw8BhRNZEZJ
JLyaPtSQUuYzjMb9V+G5UbRFf5kyiGkR8l/6Gj5BC4ya6K+HobfVDDAvIWBDUPFlqKNOKDytXxoW
xjGWu/oVWDqqtg/Q+WITubVc1iDSL/Wewqzf2P3wKaaB3WSCMHVcp8RAAtSsXAv6w+VuLGJ7XfQw
53mRAvlKrWNoF+GGuYhIG9Ix0C6L7LOa+iemH0ElN7lDv3vf8yqYjyG8bjd8wMrDx0y5S3XR3+d/
Gnbo9M/hpOfG8rsO1Sar2fLkyOW/2QaNMzVe05yzPWUnqEwjk5SK8ZlXfNK4T8ZIOs0c8TVPZ7/2
qp+JzoaUVlT+78nHL4d4W9RZ+98QX2q351INLH0XMm3iY8D/7FmfpA937+s79IzdHCDnVsi6UW3P
hXl4bnh9omEtmNQDQiBF+ECoHyE9BzOk+bFWyuh49oyM2+BocLKDIJM9r+MNBoRJEYpaO5lYDDgr
vjNrUBgrlTiZMaE81OFf3Hz6z+TYKWFU+k0c05JcKY5cs/zKCzbg5ykSDwtVWR23mjH+UaPYj1m8
SqqTNK1Re8hPAXCuxJTiD1472ZD//8IL84AxwwOjVucO19E/5V70yl3Iy6d7uNkcCkGQgVOhppjn
4GxYxoXIJ/w/MF/Gw3osrZ/QhNY0AWsW7PsETG0miTnxI2K+yiqgbPRAkNws8YKtmCMfYHYRwiWA
3twKwQWGq9n9lYrdVL/Put0oAOIOIeI+RplGhOTdiDE0D78Wwodf6CPtd/78352DLH8H4g4T9TKg
K/GR4aNWFjRQf3DK5pbqqLgUjhUT05cY+D8JGrGtpi/pPzl5RyHU8IM1PWnWV6Xw3vCsgDsLVJF9
eqBnI4bY5ZFALG9NLFNGY+8qcm4qp8No4FGzxl/DKAVlYPNMImfy//ELC+w5sGYsSXbHn1Ielg6C
5YJituQtp4q37TxK+eBmE5ZeTGW3YQ1tixHhO2vTmrOeHfLzV6qCD2CfrtMghL6RoibkRqpfY8Ei
rE7u0sb6kg8K7JKYROLewgGdqfzPGACTVMfQ9+sCf+h8MYWojQ+us+Jr9XIau+qm+0lXTVVtwNK1
Sdi0yP8m2Y/z26EIPaEtoRbceL0ekb6dRvCjajVyLnbek0o8Fv10gO/O4jkP67C0CEUpcQldcqh9
83g3d6o9hivWd305qQ3ln/3W1ott9RkkqSYuaciA9yV80RhsSGBeTEr1mg4z01KBWbZL/KUSgwE5
VeIZN3YMBxNq395b+wES+GyEviH0/cG/UgS7/b8GvyTogeWIHZw8BlaO4kanZHWjY1MMlpykZGyJ
2aKQFERkeg8oq8sL/KAU09rGVizNVm+qB+opnowYMEjBceQeMmt3mO9mXrK/an3ix9nrOHU3uED8
DGyQqQag7yraQwxTa9DkDqZm7izBwMwqta1V3CA2X5g8uqU/bOHTmyZ8cDCQpbF90bTHblGjeEAf
g636UFmYE+LRRCbeFkTPgijKEkEfqwoP+lKaVf+3QNSSN+y5WVIlB22kap85HP4I8KrSDbW47NLc
h3n1kiHGhgVjAvguvSpW3rMiZKJNYEQOOfcLsgsFlfVNXTlxr1d5sWdwwM3jsJ9fR6eALHdmK2oU
hVdgroUY18Sir/C+Al8SerZLzK/m+/lK9+MYtPQ43y17+zywIVcvUwLtS1dkPlXt+8QCH1eq48GI
vgNfaLzmny7+ZxfIlgOdnMJ4MErEsBBku41UjwxC81bfvR2BubldlQukRrHrH6JyYNp8PkgHgqEL
Mq42vkG8w0060LlThgiM/rd4ATXyJeg5uqtT/Hry/UJ2eohHjn7KP8isPwLKcCMm3PcmKNOR/CyF
hrQVMls3XTnVm1CkAclo7/QL5hrkLNmqHC9bAOWXiSmzlJj+T2k/5hPwiszssSG29xCZ8QAmOJHn
6Bm4mMeecHS3a2LPDYK6fN6ugu21iVkWgRCTeK0Jp+/RCYdT53cVm/bNboGh8+SdwQ+5bNtto9/d
6t5EODw/pwvy9PX0/mwMakaWSinNHnQprlrs2mZnE+6kH3E8nha3sF34Pt84HSekflWEw0fA7+Cp
ZxG0Q6Ivp8U5ARNrSykVIqYtXWvMtSTTWKHudmEYJljuAo2Ql24NfGM8N9sJhL/bUS3wt0HBpCvI
XeX9zXQWaRUSWwfmRiSLyYpbtoN1R76er7Fpfi8f1x8q9Jq6YWiAhrpWSlfy/qn3ayjxPm8cELKW
wkl9ZUBaBRChzbUOKocFaYT8LibJ3lEXHqxwODBA0KG5kG7OQsq2baf6Awmyll6lfZwTMztRZKea
l8HgFdrXGbtoWmsogdOLFd9OgnkBaQs+QYwYKjSlQXPVxkUKeXKn+5TiahbJrJuj6eDde5q2eazx
PanlVWJPy7kOhLSAjoONR6PjqgK8JXaNX2Y+vnZbSw6ZI2jT8aO5hY9UXF0pOmAbLXosCjKgqffH
vIMaFPMmK8PmmApBPFwXLQ9JMs35H/cyM7ilEyIzRfD+/JIkfwM3+lOd3ss5asOFtKZnvX8qM1XL
4iD42cnvZ+Z4dqTbYQXQwEY8qJcF1gLvA41ixrZ8Q9kLi79nWKaNxXR8uEcHsVSVI26YtL1MY5eg
Fcn3kL2GAMo77gmP88gyhAumrseoZ5QS47tHBBUggOG67Z1z0lDC3b5HV1fecxOeeecnISAv2AoX
lzx48bLHxZMUdgkpGWHxmTZ4O1PmqIvVt04r+Q3pFZkw/eJXOv5oj/AVs4YmC6IhHcdVrzBfi7kc
iaBdBfWfbxjWf9xbhRGM0Kk1flarZfurTQBPIZkdZkX+g9/41O6JrmGE+V7vWX8Bz2+D3c4XeIYO
JTJBHtrmorPWsDGFIX4fkfzMu8Ipfx1sRwVJAdOb2fqOoI2QndqoA8BJt8309m7TyQsZq0FmiF9L
jRuOU5RjPb0aIJ0ATelMc3d2Yxshp+Z+uHRf4lG2y2zmmCQNt5LJmwrz2tE8Cb0RWKFSIb6GJh3N
7DqRJUKt/5CXYdxovjekNEA0YWngSM3pglRYspuhBLAPBaLOLLuc/3dBigsieQV6yEYzob6mCQXW
vhKnYJQzrhwWC/LyH97SbQi8tQHa6prouRbpnaXXhskRh1NebGiUmHQ/ev9pAkZsORnXXxHJFd/Z
rz2lpBx3cG0H/vRSjmhqSElTlZNq4R2mjjAXCWv+mDntd3YKjtlCmpxa/Rq+Y1NLK3DxkJLhuMkH
ZWpcgw55W5hpOQ9a2DbpIyZcJ3NQZFxOcYvZKNaPhZ62rx07qnuxJCT3YyFTggwsWcIZ0J+K6EOz
6QWmJ63f/xJr9Qew/lQN2HBgIgKHsyCcQdcc0Kn/OEkBfvKeq+jBT21VonQV6XdJZ5bpP0G3eh17
kmwi1j95wwS0jTg/sGAyY2MOGZZ9AZj6LpjphXoLPhm9P7zxTgdu6gMsEJLP4nMzywRfMexrToxA
LnNUjpjs/vBNR+6fJGqf6HbZLx9ou1YB+GZoyKg8BpKez1TeEkR/VjIofMtiGrpFxy8IZL+vKk/s
G/tTvhYleJb6PN4Qu3B/cQGhH5YxTGbqaoQr9ewgqJGdOru/S0MMsZKS1HajcBkz/98iSdAfuCuK
wWPSAK/u3HUnlbSZyq2pLkPqw+eiGjm8e9aGUO0ml3AdQxzkv+vQ2skTg8rTm3TVUvxEPgF+DWWL
Q7LeQzMuBN4qHB/wGqxy4AadpTnV+Jnz6E6sqLy4MvyEN62Am3w5RW33pQLeoKZJ5+CZlguGdAit
YLoFFMtW1rxFjyAED2h7/Du36GTfzPdi5KV4gl3Wk1OCi8Qkai7ql6FnaX5RrmCMCm/o/tNxRxYO
J/1OJBiJQZe9yCh1/hEHNn97ner3gamUV5jEQlexSeskTCo5BuW4wug/ChYthSVUBmFTS1t7i8hQ
j2qBYdYRxwmRT4pxaMepMY8KLUM1zZeQRUy7V5v0h1TW6j0SsZQGzgFMPSM4GWKtyXbvzqhKzXLa
SXPEJ5iy36cho4/VYljK5rSYfjiYbuzOaOPvgZYtlW9vWfRvnmDII1dpZ2zjInEUBVyEjsv46iec
MCxokuWdlPgPzuaKPJlPXO6a7yOUatdJs61mRd/Tu20NGDNc0mS3Wt+oo1wVUOqW/Lhh7ooydi35
unZSO5YMefqSPQFfff9Ne9xuhYpq3MiXJOwF/F9UQHfxg2HETUrq+ffyx6RFwN24TtksdpoGo2ek
/UIBv3ybpgISCiefuaAHb5JZVBg+aCPb1Gh3kfb/7iTWv/m1SOdV9Fp5Yp7K/+3HCVIGN+7z3vP4
EzK+EF7oXTQ+wUtkDZ4/zRDlV/uGBidC/W86nnZmFk+uiaqpEnxSiLzD+e2zfn33SLuTBe8CRGM7
kJpiNO6jtL+DwqYfJHMrZKcancugfEIDxZjFZdFjpe0jUaUzieGANQZqhTfrKboU8IfHEIzb+bgm
wy+NcF/h/oeb4TahX2+m85S/zGzJzS7T7b6sXKtSlPHJNJV0RDLw0bHs27p0M/kI7wcE9CVkArLB
4dUvD2sWhnd+P4tKG91P6ixr4bQUYSfy1mjW/RG8I4zjeS/Z2ZKucisRYpXc17dCHb3DbLjitHQg
oQoPN62nxQ/jQYfj4J8WgF5pbQ91WqL9/Ml+AGYPD23CnXhvAgSqxSEH/dLuEdtnHM9YhxpClIkn
agks3BPegv7/mBa7cy52qGVzza4i3paOqCwD5eut4YncI+rTzAitmGBJg1EQf9JrGvtEfOowGPfr
RFxOm1eivxTJQOgMZRKxqwQW0yX5TbhqP+fDgUL9KO63yBVFi+BzW7n1C78gGtPui3DLt93CoQ3m
tvb5EBhdJj1ZBgRS0CpEclmhUYAIJys4+mvtci6Fdcl9pz+Tm6P6Jj93TXlWvhw8b25yAGS46+ib
RWLDCBAbLU9GWe6m9JqKzZ/ZjtOhS8BR5bCGWPDwXkYlZYp05+aEUmhhntZfvj4Fh/q6SMXzYHQ7
tJhaXH98pKxxJkNg7fEU1rl4Ic6pwB/ykxwJsyB3q5Kdz4w6xNXnoDupdn5dUUJ3KGcYlwQAG4kJ
bt5U1HiBOfznASUjSB25JHmiDExwf4QGfxkq8v/4tnCdg9Dlmtk3InvWV3Rzwlrl9Q2ZtTjQ2/sD
Pm6PrWOJqUBeby1/MLpZWmiOO7KHiUDh6sOh5K4qh9JxWdHZE5+LFUe9CsitnRI4riEX1bipMnaD
QKTH8TxBAuNFPjPiXDga0yNj7ML8QqtSdb3CdrEd6oF6f6xZAABOBH+PEFqFGiTm23gXj48oHius
rYVbjWkqJqvnDacgvoYEN+kRZNORpmXdggpCmKnik6vCR+zCPE2l+hW263qaNFDcH4CeeOFAO6BO
DfwvJ6lM0iBxY9YQsnXLcvMfHRCn12HEW/fwsskJQX8m/QEkqV/PV1uxFctNpd/dEO4zBonxXbcB
2ykDZhQffH2QVzI81hy8+cyNZOJxEkFhOFFH8+vTYtm6QL5Qh9TN4gbJuqcP+/d+A4D33oZuGy9W
1RyXVlJyY/C6LIAUS8dFwDy6jG0Nt+HIXGMcb/30M/nKwZ81/i31BJsgRzc4eyKimzt5RwH9blbH
aGFUfHyJhwR5wBzvWYvvXuv641D9/ZoFKS3//e3wahTBvSD95C9O+hp0FS7G9x1sCz2pPk2uEKPC
1x509rpxcWaHs4Lu88v5exJ/RxDUL1MsrGzhgQSGXNeMcoXt/hxd1Po3W8u9n1EQoo7auLVMCPro
52CAoO2v/ryjuCQM4iYLQPE1z92TJop6WWWxxfMRnAfgG9BZNxObkENeKXCl3D3BrN7tGAHTLdaT
XIJj44/WRQivI8KAtL9dnGOnyc82Y1JefczCxa4T7mVQZsw6QsAz7Ul+6QDOhl0yw4iivfP6F1Y/
wlRmgMYWKlq1ZyfAsreK1BHWDLioki2YC/q/Cux6QkVl050uzx84cU5GKNb/AKqcfSnFjeZm0ozI
8PqwDLemmU2RtHBI5oq7U5WKd/OV8HQHfNz6huYStOF1UJIsx9bbML1w1ccp/HlpLSAmKZlpqzvq
Tqmg9BUCyJHk6n7SVxmwt3thALVxfWhh2ovzna4+8e/S6vI9IGY6Ms0d/VMmymepn8686UUaymLv
cKfLCBFZz0uMXtIlidDXeir2UD2uJbGl9itYwaoFzCeLXRpkhYABvkufgbJETXggQFLby25sBzJP
iSxlejA1FNB3s62CfU0M1JoB4mrOzGlZ9udNei2OQjGsSoeDnjSMZY4WQIdgZ5JOIs2BAovlstza
5oVLNt1LeeBvETha8izdcR01WWumnQ1eE/GkqgxtWC7+RCn42y4QKQ+DJfisMblgaxD77IxlYotB
c05dpXOdg5TBzbthAh3GsQQ2C17S5oo+FJ50xDeuvDGMuE+NdRumRJ0kTVQErW2Qxqi5h/d+ltxU
jbIIgmmHCknfXnwA3O9IBfZpfREvCZn4CgfsTclhsiHPcW4aDJdGa6kykm/NHmmOmq+z/WVD9rND
zKyW80IUfI3/HNnBjR4kH7g/WpoExRaQZPEj/n7JCLuBnIwMwAaDBb35NkUPes3/ljoLcbctx6F2
7DWzq0O4PaqE8aHkZi4j+JVy6BWONm57DSbKmY679aci76hDObHq2ws7FkQxVtq+tVRTAl2PGgi0
koyigmp0eA2Wqb/IN6oqRdJNXT7gj7HvXPeN/XIzBJwiR4A0uYfUf/57Nbmw+tqwl0lJaf5Cz1BM
BmMsG2s3axJ+KYjSJZojZBW9KvmtWrlbOYzVHUCUPQOc4v2PNUrElhXlZ78Sz8/efPduIpXjyvAF
wpvY8odmmDUqW9Vxmp0yDBppHr9s1uaK5M+TNapigm9cl8O6l0MtX/wppC35uQd/6H3OnyemWSG+
IKGOuZXP8HTAxRsyELBUqjqYd6mYB8mswlDNjWxIE/BFpGezES1YUxavf2xVsrPzVa60qG+sE80z
SRc0907loesgQPyKP44pvccU0lp8lWY0m+uuqcr8uIb4Tjagbo4n52Ax3gHUMhIUULwi2zwLGCsP
sQdV3w+yxs1izom71SWvhVhreGTBmbqyl0icHFXg6Xo563zPl3gfKJkaxMRnWN38lR5A9ukb+5FE
bNqKK/8rqzlgnYrpswnbJRaONsNssCGBbpkUnfZPjtrg9goB8dlVoD8jw1EARSZv76x5Ho0mQDSk
/CNj3xRX2PUw1pMeagzXd75kBPYaE9bJMQsmGnsdgWNPqQb6g7yI/6+US25uggH5qJwrP5LpR9i8
EV4uszqDqDAA3+SFyDW4LFO+p0bCFpmRbhfK6uGPhhNp9vq97DjZQWoNrQt2nlnRPoo1AvNJsR48
3DCp2tgj6aS75w1flPAXbz2vkUxJwMXhj4HR9BnLcdLDBElt7W91MAhTwdzUtybKZAxV1xKHXaCN
w6HckSsB3Tq6vfhEs83LdKL9vWBUW6D0+9ETTRry5shrlnvj1R2xnqqnU0hUBvhWbKx3Wf391vco
6zVLwrtRigLscdk7aZ0rvseMxVgH+RwjwtaUV9GYcbtwgJ2/bsFHRSB0Qd6jZ/GptP3lAS/fCZEk
54SrX5i1StdsqdkgyD9uGtXK/0KmTIH+U5pfCYddUTzKlmF/bHiR3620CZMQnhBRfA6m4WLGghc1
CzqKXftzr0BEtpLNkIVjrkrPT9nEqSo5vhGpEB3UGnTMQlWugMdEccvjyQ703g2RsiMNGMfy/4W7
0y/iAOOMSkHcfbcJOH+iUqQncaSWW96Um3rRWLzaiNWkrDB/9jD/WnW8wJcQe1Nmx1RVbXbQ65ul
ymD4+d9vhimz2W96J4WZlYNKbBjiWcIJxe0uIostVJug9vaNXGmFnwMFQFEXYFQeSgr0NdbmLNnM
zVKOuMEb41lTMUCCluXSmIR2T7J2kcUIwP4f3UT6BgVZsLIgQvVBOeafWsx8TVztw5zJBSj70Gsl
ARAY04hFmy+i6VB3SaeXSBlEeYrsl/W6zrxeHF3DNrUok7l4PvYOWq0pe7bnxrLLB7/StDQmzDQf
zfCmY8gHDmyRso446NH7kJjvZgAi+3mJG66/GiywQHiTQYZc9lxQlC4YEmyyx5PRuTggtDoe8xiC
fuJbuM8k0rncyFUsCPdP8O9e8+VQxH+NUWWwQYRJJXZ8M/nWhmdhyQnxz+zkmNZbhjaGO6p2+S04
bsPI/adxhQEjraqerynN6XX8uZcXODpeHc/8GM3u8dBWwUN6BmX6i/c/z0wyMIZD1qZKdsVwZIWO
gZ4MO2z/QOyfgBf5GoQEi/zXm0SQtpdG6ZoJ8CiR0EIKKxXqY3ptV5P6suNz3V0n4qFH39fQQCWA
jKK3AfQKDDuCV2bgJI5VZKerIIwtn4OXOWD+WxvJEa2ADg83d5z2ytLcmsZR43V2phwr5Law/6tU
F4YVRgGU8mKnjNln0R/kl0gZqpdwUR8ceKJlXv7t81+3D7LAR598DHwzcsiz78jgOM0/yw4b78lU
ZBNC7pOphXeFP6wg3q40Iixi+6opxPnWw2VYQZsORsncif1YPAfhNN63BDwWmf/WIUMu+k0ImSXE
l5zd7YP+xeixiNvilDmKFsIX7zvLD+66JPQTvYmPABYtQ/b0uXJMC5WIYPeVkEAzJB4x3Xc+WCWo
xHRRmZ3KhBLngpHFDazl8S4MsafD/U4D0x8h/ca1o536W7r/0G4BhtaUSDsCTzQk+eHHMZPluhu6
mllbgqkQ/tF/sqDfZvCIH+8yBtaL+PmvbnMqmYwfTDa2A7yHsQq6DTdInkbYqXMw4wsoJYgPhTcS
W11Zni5+cciG+T7X7jLAzpFo/0YHGjnnrblGcck7MD/ddiWv21bE2eptzjHKzCqfXBBVso06S1Zc
JeCiNBpw43UCYhnq25NbxAKwcToFXb/qLTovOZkQVAnMWprkztScINp/aJXJuDwAGWPFl1KstK7G
/XCih0qMQVsLS1dkNpLb47D0JmP8XRrqotjlXhFtMi8GF2yaLfB9YKi+ym1K3Cuj3O9Zo5THXRON
8ukQl7ty7lSWsDXG4GJEMc65eG7xDAdkaY7OmbU4+QyIhXtNnmSz//3s2IGj+xm5upRsbVaJSPxQ
q8gjouhzQLOttFMrzwnXFcTHQNIy24g9hR3UKin1gM8lYfBoCC3mngAoEqX8mJFizvJeoPlC8t/Y
hwiI6C5zysclKuCZ4eMWvtMNl3vGlAYTNOSkDAKHAMBia9L6MFoizGUzVaAtrGNuYGh8796wMUoL
9NzrE7yEeK29cDaqiiTLlC/4AEx2rzfHvsJr4ddLlyF8byf8H0XcNsSaBIpVBx/cFYjpBCfDYUEI
/uUlx7T0c2FAw/VZk//rLcX4lWxnFQhMh+PxwYcgU3aWVX5ze6V85DXlmaw0zK63naP1iuJ3COGJ
mysA1EVV7gVslnmK9h7yhNbSmzOCphzOpdgMaljmOijkYU6juW8P+MKARGItldgvAuL9AZApero+
qQoRUY9Gqc8h2co+VxpSYPc+CJDkx6QlaaPZBw3SGvsEoKNj3fRYz+cWCX8VzU6MtmLSPKMwjGLP
77K3mmyWeTX0Y54vcAN6btoMLCeKaUaDSjJMBhcgyR4PcWrHUD1F9PKJcFmcdOj+9GEbrNWyUDNE
k/Kisx39Xjy8315DBhNut2nfqLGuQV1Efcg7GP9gVnrsbcT65HriXbV5Yn9d6fqhhmb3ZiHJ056s
iPtcp1gGNxYHw01EQtydnoMqGvfdQAe3q9/6f53c2IR7xa1jVo3XXhZfZyqgI/0O1cEpeO+TjdYM
nHZ8CR/W2d9egPJ5PXQFSGDF4M1Tdp3NH7y/C6WkIjJtmGKgJ2yYc7nSGyeXV6GXtIW9kP3bqkza
RAXk7vlxSAW5VZhfoYgZ9j29MBZW/7dLpXFTq1hu7lgDWas2xKvtBNSi9mb+CzH9iGAPpN0iwc8g
84AzHN1vUh8wNqG0mNHYSfwmIyugAHy3MPQI1jCQFUDQWTb310+RVobmewNQf558RCqTv9FetOGY
mhJSDq7ECD2QaIjh6puPAtyJsg2KgU3asCDMf+hSJRq2+JSgqazBgqeIkhgfNEafDtgypmPwVQ5Z
rNnrQDZVGUr1AXirwuJ/cn3bMN1ms7XJyrZuKHU8k0mDeNkitsRHVjmb+rMtfvg975bafi9d5Zb4
NfvQoIxEnFvFfqpQeMDvwmiiqiWAvd3/zYOddM+Wt7s1lqrmTvV69E0aYcWTTlWAUmUIRAYOxElE
ihXA5rN2F11GSsKJneGtZNJYVYGIvvAyTF9QK9jn/oQGAcQ1e04EPIOxkClu3nEAc5ysDJ0uoxk0
4utXEAAk+xDMt4L/zx9N0vYIcGSKMLVL6CSw8Ay4mfN7Tz3gD5hs9B8lX1DrMSIgQC6H+6LLKZQZ
YoR+CunlbPKCQ5s/TCL1U5uDrzEuA2+7KEHKc6HMXy56g1hcbx8q0S/zonfVYPsh0KadprvcLjlA
imCx03uawvYRRCf1dcrS64ofezop7tH3FdlWElluPuu8fnH+881jkryoR6UumvV+HGZzqEkb+g/h
IzZb1NrmtSrfgKohyI/HEr2MjtqtL/5bYFvJxClHNJJ61CLx5VCEUp7eigecErSeDyqNbXHbgWQX
ROomg+irz7njb1HnvjVSzs/04UuZZbVHPqT3+VWjtj1+ghxZACsN7sGzg0k1AUNPw9s7OxcbXg9P
VSYVvYUx7g7eEZmF8Og4I115GWu8XSg5saUzt83f4ugl+14Lgdcw1bJjkBBNpyrcEV3WWovyyY7Y
AjUjNvINx+6cL8vBVRDICHFfpOExL0Xx1lZ+NVnQloOHXWsD0fUFyU7+6cW/5sFcvcbg/lubLd1M
Fb7mZyHDNFMc1DvS52g+Z1c94Xpg7iMHCGzMYC2KYQknb4mNhWJmncrTzGqxYAle/fEo+ySMF7Fp
EJpv7NmWVs9dsG1tSQEQHh2/G+SxFORY5cuCiOfmucz+QVTipGkhX2AVUDgetXkUT8SHgWGLPlSM
ir57axJUct9LGCUG1uWZAGN4vnczdZHMbJ5PGDQnrP9vrVJBoFptxv6P3AhnjT1eeW/bMnl258kq
vrOn/QZBfdOSOHA0+vMhqtzVnmtHC3hlTnCAgie50lDmacDdF63jz63OJu5pyjP3h3UZtI/szbXv
Zu141NOq+dztMdC2OivaVTabFmLt//0doltmGWzh+ePt4MRqZ2w3SY5FhnLUHBUdyI4JHhwutbUv
sWVpHBAG3j/NKvEmXFH4lNuS+VhRktCzGNTU1WTr8yUQ9AlX8zSrLJSUqj3vl8qvf6HTwDgEqP+s
qmJMfxP99dZ6LnnB9cAdlV0F9sT+D1tQH67PaceTGOsH/eyQ8v8584LSZiOo+IgX0P4CP9Fv2uhC
KRSOh3qduXoBgFhLkj7tq3IU9Kq3+I+o4NucmpVam0LYvePjGkX035oX6lb/gWJN0rtWdnzNYi+T
K8eTDYsOvbQPCLyDUed32bUwzCQegFLxsy6jUfU+ZWJ4kN2oMLLzkbSsnT9WGwTCg9OIyPFlvuxy
EWSsJL9QFL8rsECb9BdPZP27EUtRaS+KsFkskpLCGyvr65/tb4kN5ti1fxICB2f2eDqiKkUFzKFM
5OQLmeNpL4DET6jAnMtDFNVlZj0W8yAw/rye9f+EAI9e6oziaHCvTv4a0enveVrGR6jSeVvEXj3R
5t2zx/U5L6WEszQTTmimTexC+z0WGwloh2EvQOARPDqLrLDpYIqgKi3GuyKCf2I/Cw11K4kLRRxv
F+9IVVGjhTEvl2TG0PE6qbaxHK8qF8RbkHcQ7xsWRc9aZoyGza3jNWnUPakG3TNLSdJ/lMFlMWRE
34Ni/jIyrNlLVpXzjW3r3+puehO0OHBsCSiMyqkx12Jky5POwJqIgOORrpAXd3TFxwAiAq12VUZE
KPlzUXcXBdpFbsKHN8YUGH5bsWPRgnCO4lhw6cjRLQh5V8f0RMhHTehebntJgECYCdT/hkONaQEZ
0p9/rG7mR+SSxGd0PY7LVFPaI2dIiiGBBi/4Wl+zGW6meS7c5dtWT2wY1it+OnaguNFjYKJ/LyG9
o2Vpq1PzDC4nXQQdR5v3R90HPPrN7eyGRDsyXPyQmARG0w78QpwEmY3Us0PH2T1d+ixmlaSZaVNy
4thR19zI1CWSg6HpunNIMH8ZwDrg14rmuB3PMbIUTzTCZ1Gt81c5zei2MRD5axbxIiq+KkvI26Ay
5pVPrEfKffagv/Jfy7otCBHBrFccerut36/CATGrG6Ht9xMtpPXBXyoq6I3cmnjYJZVeKiepK0LJ
n03gVKgguTNcmKy8GRQqFLRp+eha5hZBOVCUfx4GlrlXlPXK8QzXwUREijERDY4JDRV9H1JGTA9F
hgQin6M5UrL1t7ykHfsJCOce5Va4eVOt5Z4uOI3riKjIebvUfhAIHqnHT42B11jq+H3jZDkoW5Yv
yMYqYBO7URuM/RYq+m5eyF0xp4IZxTLzDlXCMpp4F3GOktKyHZyDu4uidvx97Rk9qFoKizq6Dmhn
Qa+KT73emElzVXnsoL/LifxGKd0KKY27/aZd8rQ+i6M820HhBix0rBOhqun6RV4aWZb9x7u9MUxY
h4kZj2LfKowb5BVtGmaOT2DphPjPzhLifwN0KVs5vq2ZMRH76j+e/s7fVAqQcxUDhAFYajK0DyGX
Cj7VqvC7xiFHgS2OFkqn07LJpO+3cYchE8ft2RqdIHPZeWw0ixhJEJt7+LcPerw8ZovwzsWSQwTe
TNSEFrFCIpJWlgzZNQYC0I8OrtlBexFWF07TuSJiZI+4SinBxeF3JEnbiLJjtbSm4BYfY2WBdvSm
GfACJI7aXZcgbIQqLQYM9EAtk7uZEHXMa5T+ncpbdmDmdwb/BOrUzl/kU468XBqgFgI5l54U0cHy
85m4Ke03RJNbHCE75Ixq/a+nQPOQkJApjQYfxPZ5q8PbD0bJCkl/ZOnLDmCN+X2g7uzPc9NWZj5M
1SKQ4TwGE5UnG6HxzFrU3oiui6sD7a767AwBBYQ9M0xF5oMrlXfXrm4BDiP+cKcEaEBNEKkiMhOJ
ywLEF2jhgashV7slJWUTHZBrhWu4uCDwUKK+4bswGNh1NuMLCPamHSJgrc0K+wx5+Gqj/OQbCd7D
zxiotPgTaRRFLbcYmu/qdLwzT4TCae9J8NOKZOpySWyKIgYs/MbtUrQuUSiKE9oS3gCMOjHiKpCD
CpwzwQ/Gq8Zk+dO6dfz5H4jvPYKAsYdijOfrp+iQbJbsF2wTcUt60ZvWkK0CiHoL38MgPOgmuJ04
Ixi8J+yPVJG7uEBpQOCYD7E6kOtOGtcPs8OtHHjCJH+ooC06vAkITt4xn14xkSc0bjH18C8zw0bx
PLqdTul7Pwq46E8bi158GDLzCH3kuMIF72REMyq6aH8DVo4XcwscrJLtKCMNL5XB8jAU2jXvCBOB
eGskD1ji1ZWKDwIsu/s77WPZpgQGadddrZkG3TWtDJrKsNdnFnCfcnZ4Y5kypKwoSm1ycSnKUeVL
ciQwBgr4lvSKKULj0Mohj9BalMfEou9PSJqlMQd1oUjy59PabcluEZH1mv7seawIyETYs7sOj6l5
2r09xfkuPvv17BTCwZTFSB/HUEpnbO1nE/zfXsoIDlBWdzir4yf+oQv1ub5jc3MO9vHq1753T/uf
owYw8VCPTgXlaKbkjx2WFPQD9s265pyApeBDYAPRd4NQu9DONE/kVJ7Wlek/kfcuEDLnJchV468k
k6yS98OUwrpIUmSZi4ohYYaJgj2u9jH3fTh9GXbBHJNHjjeXSuZTPdnNf3uK852Wl1uoRK5vPt/N
kQwh/nl3nQKJyJtkZ0DqWIAhfChXFrPkO6KVBFIumq3rpiaw102k3YRNeLEQz6nKW7Qp0YicvVU7
ANar3l0KpH+IgCw8w7jmsngeXHpvdRk0psGpo7GE+i8cJjNq3PWHoMD4O4++b33CF38Mrj5U3/ab
jqmp5ZrKJSxR5+mQLElrYjOqjPhcpX8aCznymX+UVwBghFwhcDlSjeLdENR7Ac9do/RlzdG9VOZC
YpP02Kognjvi2AmZsjOdWhmvgTIChyFk1O/6ENXR5nlWI1T8fm24xlbhREKpwT3Ng4TSSlDL1Hzy
icMa0bSKiMP+2Qa8N1JsJfYfwOYQgYTLxxxsbYmPRvW3X8/XLgqCp1KgIUZIv706ZXdBPLDSUwzd
sy9R4DZaQhUn7f5FkUh0t1xlDz6l7M+vK9eycWP6jI2NEOhF0/nNPkFO3dDJHb7GOc+hgqCiqw9g
wIzpEyluVWLU35I9EEPCG/Oi3dIprOoBzz8ilObGeXKOl+bTQ6HwHxlAA4hd3LPP52dJU8xNRazV
tUeHrgOelxNsRgFOhG1RCdQvwcqdHiptCglM0xB2xmIaGhA4EOIvXZrJdao32r0vX/hibOUpIwpO
mxYFwz45ct2781Y3dpH15ngSj6MB8mqdYuIjqX7rzJ7sTPgZDwBjVCFg2DuEsKze/0CAMQkUEV+s
o6ZSFfBBY8yC4j4AfsqnBl8RNPelaGkv1x4OPbUCnI/EhCVOAx1phD5GRW1yzRMjrvhjVx0p0tXB
8x9lT0ORv9krYbVPIW1bWNGJVa6aoD0ocWVo344cZee8eeCAoQAsxfeV6KUFWZAb50wnUjkdEh90
InsHjgQ4M5gaw0LfbcW7Utpk8N/R0WKVqZOA/xAnDRgRQ8yDAHjv2dmilOVlWltH8H/5V9/HLVbE
mWDd3syym9ztMf4SNLe5hA9QezjC9J1Q1d3tC+tkjfpPmUj/sT/KYwa7Ulx2Ovv4X7KVIz7O1MKs
Fznxwjp9DOh+AFcIrMP7iTBtTqAoMR/H6Tnhd2k9xMkvyyvSea9FuLro6gplmp7MqGFnyZTqF73U
srI2YsvL+XOT6Lcf2I56FNjjMCTKfJCnXb6sjnZiZK6wegFe7qYOcB+VRw4jhxzBMb9WuDXd85JZ
5pdO2KBtH1Z2+7zLy3xw9Kdf6Et2MnQzI551Rr518nMniY1BB3Y3HVqbrPJ9qsgaOm4jpdHUGfi1
pit+OuzVFhgLZ+LMcr2RWPar99atwBh00MDKnnrrrL4gjcSinnahKd1hPT82GLUlssq2/7ZOJFTq
UMXulMuDsEoLX/CCSbahiHZMNLQcXtwBrXlZ0ZNH6Ql1PKSdLkfUr0OCAzECHwBOia07ssreh4F8
6ouSDA0dFiiQynZnK5ghNemutrsY2bnN2Jk+LD1S/9V4m4M/10m+CPK/7ua73zxgfrJkhgmULI9w
M32OY2+/hSKI4MI5s/ywCUgSN3SbkDuw/ezkOGOP7afreAP1X+HI0JxBOslp5DvumjLV+Hsnq4j0
ZHZirqk+uLppLp9DTCujNMH+IZCrXRSDrDKuTIp5ykWLz7luVHHfISgEOkxvAHFNrn3qo+HSPcBw
cchQJ9rrUm/AtOxREDbf0Jc8Imc71wLr8M2uoJpoE2vGlg/6fKsX6xHpqtuGRi1DpcURUbHJQh+a
/cYSXJJoWxa9XOFOcNmkjd//kQ+nGHYxt55g+D7Dqsb4SqCJ9ahJP2MPVrmYGGGIHmjnxTU6MxPE
bZflog06I375KRp3SyaSFq+1kBRHOjHxg4KPPVtEX+UipdW0i6P7TXS4AldR/QS9yU2gfQAFjE7R
yi0sQX7PlNWFKGWNZoQSe2/gFeW88xAkmxJF820ggJD5r53WZ5wMArFU8b/u215lpZxW2hxp6MWF
V4639TsrNUV7lrX/3leuLZWKYE8j0n2OXtqRBHxDhCtIWIuaNVP+lONtvAAg3A/bkwMGBqZlei5x
i6Q/Wn0T0IRwx4m2CQkI/Mk6tI9xMB0Lysyicn6ZCbifnIswErCnrKTHKV9qvL6IIa++3mgRrphz
UP/KaOsmRdOFwjRiYITTO2QbmS7YQBTMs4RCAivRdngzareS0cSf3ScGNy+5xlmUVwrhq3eIl8ry
PL+8W5C2HZ8ePKVEznzg2DAPs9PYSy6ukai/jlYtQGDVsheGACyEaARdYSsb39R6qcBcpyKoooLS
3+jYwS/ePPNucPLKDvtD2lyWXUwbDcdC2GHAl9uqarIzpteLpk6rBfaMELg7SMWygfyLBH0T844f
ZkaMMVozlW28iq+ocaLzYOZNymdeqgWyg0hL27IB43nPYg8PohuRVZf3Uc1XzrA9J5LCJS8nISQp
P9NG5oK5bClCJi+B7Z/d++shz+/Jjw2Cw0J3ur5YJk7PlYBjxmcwvo6oYosZGJyazNyFTMFI4W8H
h/qmtkM5BvUYgUCSO2H3yADH+Ikw2/a1h/UI6zJnhTjMWHSlLXwVCzkqjhJjGdmxvbzLe6PMEpSs
/lseYMh9DIssreLEVn+avwq8ZB0mBKEadTjv9sI/pUbb0bMlwhjwA045yXmRHqFONzpCKlTv89/w
RW/nTzFpnkEZHM58Ruo7KA8dfBSvUtAh/FYyj+NCXrw441cVmrHRnwcy9JnWxC7KCe9vjm3KZ5yb
NA3sF3pqVkApv0dYJJD+55rZxgita5F6xvw/b7kZX9OmJ/hEOFlI+vx7Bqwtvb7UdwbPhs+iLnN+
I6EOGk0ALLbq13HGev4f9aKkLTCWpf5HwPLOTA4Ml0Pq7sUUUkn6x2bxd/y3phsjj3W4a+XzTEX/
uQ6fzPxH1ksMC67N9R6RzX5oOZq3+z/9/bzwtXel9eqYOyNfMC7HqsRpNKpIlOhqq54p5xIlCcGG
iHdFU7jOsv5sIMdgpkDo0F/TGjFatafPOyabolIdYZTknLut2I7lmtqqu0jwpbjISN39cVdpX21V
EPjr/HfYPXrG1uqyWRR/mXEZHBDm6o1tZWq6w1+2eTtGLjGtDBEnJpJrOpi/flow2FwJ2zXeQ/8o
C2kq+7weCOB0EBf9GStzY3YYHirT0iLhIgjQjnQ5NVCv6O3tc6K2gQcs91Q4izjEL+KSdH04/fX/
L//WAOcIGoLbdgaXLF3vWU/XA2bSQUSbNZ+G79dhvdGtA/sT8+zvWE2IfGDx6biNxzvH9ygo0Xsd
Sc8XliM9oOVXxSp7+msVCJ/NOSOwHaGzs5bnvEvwENUIWqAM5HIRFCmav/oOsD5iGlV4Y6crwsQW
uD0pjmjjoX0S400yFadUieMKZzfF841Kig74lrmCBNFqYoqMajipw2IxtZk/Se1TBDao525pvp2I
CFPxpNODY3prXaSrkYWxNJ8QZeeSEhZQ3z62LgjJkaa5qwuHNzjU4ZgRUKAAsxqU6Us5RPOZfn6o
TnxQ17kfh3Poy/cpn8N7WexvibsS8opaMI0wCaMkOyKRV3Ulz8/qTwSKyZ/swQDMxsPrgEtpwB/V
Kz/LUoI9z3Twn4CjjtVRKtZwdyXcJgZeYIUEbMF4uBSnuOPVXybJjL7A1OnbVbHE13kHIVjb6KKS
OVhd259fPnHBcv+pwJUAqq4Qeb9fjYPeXmenvZZzPrIMAYhNbLcWo6B+t2u0ZL3SB/IFDc0/cFUi
x6dj26W6+DYuressIwtyKI/4B2jcXP52ypgBosoxLwWWaBaqbESjYDjl6Kp47TAX8WasE561DAF0
CxpOU0zSRYEqGK7oJvVWMNVhVfLAVKqWvdkScLbITm94J3xXXeI+932xCVWQeyCa1+REPEESgQ+y
xN03FffGpgnQZntBOB6mHJ+CYpJYkmuGPnct5SmlWxxwh2MCGauHbxmoAf2uX70xyaLpufaGUQty
i5DVI4mDWMcM3O0VYG5wc7K953XdCI1AwujI1IZGm9a/YYYj+SFMy4HvYSPUJPMsLE2jsvnlDRuR
TKE9yV3VJXNCNKGdyDrI5Hi2tfirnF3i/9ncwSo5cFn/qJA0aFdgaziRb83kil5L8/ZnFONnRVp9
wiIDl5N+R2qN8V+PUEbz9kl6sC2N2A04XnmNsrd6UcW85ajAD2sHwH2En/P5svOb/cXb39sVj41E
UOjguyItOfRTwI08Gpn97jteyud1ckajQEkNSKeAV6BkOFNA77G/ICMvKhuFRwHlj/K3a7p9pyqR
imFmrqVISE/cIUJ8l15f/p7OmtyWV/RwqW/iltbrwCrzvuqzx3/H2D+CEAd/WFhzopErzC0SFVir
RboxQpYGUxGc8Ry02lkzI/B+v/SfNkV1OCKxbkm+iuQkMrer6ZAqVKyAAj9tRRghT8DWAmBt6APS
D5aG4TTc4D9V5WsmJVk60ex2M8dM76jtG2/2Biz49xNiuyhcO+bysud26iPIkbY8Y3heYTEES+sW
QxmZyse9lBgEkfTMPn+kdXAgez/sig8q0OcxRSBXFzLrBnYclT1i5KRV3mJnH9SbUYpANU4XMX+h
BU4yKmPcE0C219uMfXkSQTTcydLSm6EgLM82ruQoeoTTlPsg8KS8hBK2hpuVF3O62bKujJ20efjw
Cio0IhdNFAFyJkO8QRskcex5RG6bGfHQgzumVCiOUWtshBR88rtwLNnF/70eq/be1U59eZmWB5S2
B91mEHxTSEy42EalosALs4VFZ0sUUqAigXBMzGTYfPsCL8csOz8EaGknwU58lU4ndxdDiNXBlmN7
FCdNd5M3lD9jkHBwRwXGGw2c9iWcQTepln16hXPXQJ+lwCOQgzhxssvuWw60b8QPSoR54fsIE6O8
wNB6nZE2VClxLj77muq5q8FBfDhNctjG7MkCrSh15qjDSxwUba22PpUsf8ONIz6pS7j9yzlid/jO
T0dJ2cpq8X8FaVaH0pZRwV+ZjVDMmjUyDQEDKse024roZYwSGBNGeGB2/YpPK0itSBBREqeqmBj6
XzEnh38Zd5Jm2S4NrbohhVhFH7dlMr7sKvdjkkH3EV5MqX2IGM1f6dSoeLBJbcV/hQFutqWiFDgE
Q5GwunMsUl7ViotDV9Ec1iqiflFBqw/u4yS56lFZWSHSpb1ke1V/IGIO9atQVrwxf+/oBS/ykdzr
DwkfNMdebGgrrjHYnfZ7DBwraJ5JqPZ0LNUviNbA4nPJuWFDm5xKQXDtry6bEVUgCgUwx2CoZBYm
k47xlyG6tU9qRh+VDOzaw8J6Oy/236pefxT7JX/pCVgrlZG8Xs99PIduCAcxEfbyP5PYj0dxnbH3
OPNJ6Y9BZ4wCgNRMpfoMOyO515f8sCkTifWbpA36EWG7uIRdvaHvXl1g64hhe6PJR5BHI6jaKst+
zesavleuMaLFcQoLn2gxTyTIwJEWHxlVaNEMt7UjdoyH96DxiDSCfiVvGMr3Nj//ZBHAFGVyPPNt
j9cpsnp0WBeZq/R2xY20fAB2oHypQ99cElKxwjG3Quj0z6VjBXdBDxl5Ku4jLHX8yjOoe0IpEe1v
rw7SwL2R1F2+5v8bUpeYWu6tSFPmjoCFgFOxm9UtmRbAGXqzLhLu29Nqt+7Beg7dyaserQm3vKu3
A+v7kruOdvLu0S3o6UECANc4CNIfoQv6nPNNF6BXcN9TseLWBoDXZlpi2horGRPseUpZwrGJE3p5
pC6AkOQoeeCfiORU+gCvuWF/oOy+Pmfi7cp7Qff/kRKGsEFHWV0Y1mPni7xR18hWg/0h6Kh7y/sP
2+hk5Qm1J+7y493niBueN6lAL2/JoySutBGBr/5RsjXA+nIcl1NJmz1QlcRLzcnEBwQLMRusecsq
VrKzciLFrEyzC1KyKvz/G+2rXVdfK9nSV+7gZWLENEbyhQUkob1SgTqlcn9SP0INZjTmz6Sq6zTO
oV7s5Dr0Kfo5VQ4HZ1La5gx/nYKmgeGepYG66DldVsuZuDDlMcQnmJkUL7VNWIZwefZug6nGNsx3
AGydnYPRHvNPxswLzH8U0tVVLiOi8iR1P/p93G6KZRX5IndSmXujgPfm5h5q08SzWvRPWjR+iqZ+
Wz9n9cG4m5wCIKFBnO9jMV00NmiHBIyn0NN2zPF3dnhK9pfafTMih0s0Jc110DPGGmqp0qBan2aQ
ZPXs4b6hQ5WES76k4y0AnirTGT5KW1VeoO4VQuGM5FI+Cr2jzxnQO0IVu2fRgak5S3ozlJeIEsj5
A+VDJTRkbGUgM5i2aJkJb7RBtF/kx8cWWkI49DKjNHSzXwTcEzu9L4Ro1mRmBC2ppAadfFMA93fI
WweaSQF3+ViJtQg4i11Cd6kiYbleFJzxmOv2BCucvYZPsXBHrxwamBL/eIH9KFvxTLARh3sW7kl+
4yS0m7c27timj8v80w4AAi9hie5phzddEut1uFokZSOeF80lmiSxhzurRCc7k/dl/eljAHMk42Mf
TPxFF0Eak/q64HvRPAjH6F+AiL0uQrrJjXRUNBIJxweuhaO9Cpu3Ew0Rc0OHtHJCoJg/TW9UDgzk
6RtiMJMPD41ioqvIoc5CPJI2a336fH9fbnU/Vvq/3HCzNKp3Ds9mOmIBclhIGVSDpduAsnA5fyyc
sTWqwCJdwYLxFJDt6ZtqztsEaqVy+gOB8FzN9yK1/V08aG4fty9RkuL1O+/t7lSN+aqOzrcHT0L4
zUgDjsxa6uuWc3zgKaaQk2OCcEO3Q5Y8RzEWtz0SgNyWi6So2PnxXlib4RkEpTJajRaih0TVpj0F
YPN1AS5grEI/Gy9p7Fjn1zBjHJOobkOpFo7kJBj9hcEJRpVL2daYi8ph6i8NLiTZ9su4WpPAD65A
3yYw7OPqyIHkt9gJ8H1SiNGTIkNyfK4DR3pFhXOTiw3Bbnm4Eu/NO19fF1RF0PMs6b2Sj+kxPHAR
Mg0pComRCSohxot/u0ffIg/B2LxG2wC63DY8rFVZhlgJ/l1DnQIDE1lnGsR8M8SVKo5WAErA2i1D
OkaqdQxgeFMH/nPi4mEtyh2OArf0TaCZF/LglkZCvgiOdMhm1ovaLUwNlQamrZrAbzZwWpEDuPzd
oi30VOFseQSl9ErWTTgh38gTJiVK9vRkhnW+10q9O8P+Y+cZkWH6dsslpj7NsldlqW4tg1RciRoo
BR2d8P7w4gXjLAl9UgySMZA3PXoPY4hevvX1SsCv6KczqfET7LA6BUJ+7JMwFXRmCBJhWuB2plUU
H0STHMcp5HnHMAjTlfTramb+/khORwarrTg4a8RY26mdoCkZhkDyLBqLNb+Ev9Nv2MzoCyWlK2Ub
X3twzNSishPcg67MtvAnU2UUXKJ78w5IriWCXrlndhK78xZ31VWlugYjP6Y9va51eHxklYUVadiW
Rn0OF6rtmIWn4I2VCrL0h+yKkmoAs7g8bHcVBawcReupPhN0jI94E1BrZoX/slOWz4Qa31g3rFuB
JFp03w55TuyLPhp6WzLqF2l56V8BOf6ricgyVBCQnCkOhmOiQucmEBzhawkk+K/aRTwvGYxtTAaT
z4r31k57bxCsXzqJwXwkFnsOW9Pj1yzy8wlVHaxRBisIGEIkmtbFSyMOSjs2VsKDJzLZyjHIqsXJ
devszLBKzq90/yKjHFEjvqXQRmnZFAJKrNWTvswqQF6Pll24+oCJ+qd9wMU6EnnheN9uLy/dFWCv
M5RFji+DD8vbMgL/INeAij08eCtZG+pAorgaHnc4yg06Ci0R0P5EYYrovrtqIxg+8js2ZXRtoQti
PyIBeGwlXP05GaMaObjxx3IjCPUEqmu1FI9Xbudn0LraIEbQzDHk2hegJZnV7chcAjWvlAnqJAnw
VNDZuIOAZEjQbokHgRMWGMiI0ziKav7/e4RLbUIG5FUbAO0AAupkjt39D8bFd0YtqSA2RiCfRB6X
qh/acSjKojMMCCVrBh8XeNvgJkyIpLSV3E5DWUUz2p93HQ26pWi1A9WWV+DkdPHVX2U+c2o0sb8A
b/n2KFcdlUKjE1o98gLK9XpXxLXzSGJWg2BuIS01deBekxDrnmHWKt8gLme/HLVxe8FMqjkSyxT4
Kyc9B/UIZJ1AQxYzsykg6VBeDzR8X+IjZ8ae1WY2awfxY7NFOI3Znfjj/JdFSn11FQ08PEcjGAmO
1z009naPD1KXpW+5hnSRWO+/DJjhiKIQlnHrqN+qLQzyAtqh72jtAul7g6JMMPVMgxv0xhcfXh/E
HoQr73sXdXZzaGJu5xp1ONTbvf+CRSR5I+PjriYDoGYE5etTFXgQbjE4f2AzIIGdy7rFhvBfsAEu
+fqGYFgDPf2DACC5On+XV2fISSzm8kUN4vUXnn3scX76RLf8AhjLSMcYOSIQvx0tE2y7AbE2Y61A
JTMGOyRQGdfSMVOXWQfAhsEJ/k6+tVUy03vIGrCNqWknkET7HUoWQs1g8s1bWlxk/NKvag104a4o
isZ8ZHwkqc4RHgHCpzrkF7Cae2a3wb4Zw8jNG6DS68F6MrI8i3KgxAixh+HEGMGMsa3rp9nbh8Lq
rpPoNLbVdjbtOHnqBcHz9BfTOep1kW5rk21GNr0oB0z5Ueb1cj6xl1yCia5gU3rFdHhoLUV5kONJ
zrX4qk/rjyuH43NSGA3jeDWkY5IcaowX2ZY7TilUvfE5xCxom6THKf5ldvf0ZALxlwuX+Rt6VFaZ
ap/fBclJ0Cu9gLVOaTbaihWuEqcarOfiyGsY7xw84DuAyOgwYzWjmdthq6CMUt0PDfhROvQf/On2
/q17iQungEc3LZebSd5ApP+860nOJ3h9HnRkl8XCEHfbYOdq/Nd0SE0e7CxGLDGD9yivkIcsSQxE
+x4KukWw+tfS6cLY8qhKzpXEXj1PI/AFFZtIRuJMmZgOZ6AbxEaCb85rhYd+5Ix1OCKLHsnSElSH
W1MG+B40cC5A3oSmL0ka+fb6iO3COJIsYOckRk9DxVpT8gPDdxDT8+nsYjpBPTYxu4O+FqGiWznb
JQ/qr2fLshLh+NxVbTwqXGgksR0dUkys5b26l0TDgB7iNcpSOHp+59ge6etRgE+qs+9300h/Hly0
DNHEDqxzERRVf+jh4aebk1pcws4N4bKWRuyMwmlKtjFxFkt9rUohMt7N2HM9TxHKPllAgkocCUk8
1aetRqk5dkW63aZO0QObS7DBMl+GEqbRTGV1r8vugpDLIppGAdbRUbDazdS108Hy1qNjQ/yUDjT5
gdHkouxQB4F0yfhn0UPOGYC/k9oKdCnnxQ7gpOqHod6ZXooXPmqyloX90AmpeW5kuIEsvcTOzWft
WINdrzqs4qZghs4iQ16qpsLCRC1PaCaonSHOy8kPf/ZQ+9Xf2cNnrJCcCOJZgPsR+SlP+FrVFq1b
3YHErUtfKWOKciCjYdCPbaN4c9SUAcRfRgQVcyjRjbEBapDcEmncnJFW/8OxGDsKzZNmPclTCH6L
hKwSoPrviE+ZGOuxzeHIfrcZZea/c0XbXqeHMjtviYaZLEcvEQsZzXbkCM8wYUy8sxNrkgSf10ag
fYMb8+Xm9v7wozhuNHY3MbbzUirZlXcBzM8bPzCnDSKp7D/hQgcBv8TP3kfJB1+89KnyjhiW3x/E
ZrJ34o/evj+gCLGRUnTaoPNZnac6tF3dYS4X7exrohhLnxNQbOxRbQMRjJTvsg3jSLbpgOIqRdgN
sxEXAmbCWF6Kkx7WcWNZeLRUqacuv2HDvxbEP5K3W1CbcxFfzFivPmx2GDAv5NxHBRY6jJojlR5R
ZJkNTGu2SNGR9t/pmCx/pEq9bMZpUhHqzTt84SaS5WNMSBi1sgu9rO4Vod1vDThd0HDzUFxyL7JL
yT/ePiHMzEN7B6TxpN7FSfGwfMwTWWEm/X4EzBqV8UMdK+MTVkrxs/er4u9pxtYJv0T/wYj3WsMy
Z0vPNQAGJErJ6SG/zy2DfOgQ1S7fTQa3rp5R8bH7eIQqd8cBIw9SPUw231a5t8m/aVWm7TowZLzo
lxw89KwTgGfmVVlAadWRClrGqT/nQ5VmaLXQIk+Ul5Gcug6lyFK/ywWGCwOBQVm0iz+4AupjoQI5
8+TpSjZn66q70qBXfel57ZAONRH7g2chPQgYdIC22BSv4pBjBh5YOBQa9G+SRVtw9JLicn+oc36C
McJ+VhKHqsm13WRdKgIkfBi8wlNIFQObvdrHNAjxAIPGKgUor+DnChJkZCbElywglvx4fXxupzer
FOeUMS7G+HrXsroySjF+RuG4cIFnQ3mm44iYqXA2IVK9fBshzI5cGnUt2SE8NUh/brNmfpJWjPEM
suRgv07sDJtxYmNLD5BYIN+Qy9lqW+iBIAeTIPK3Qc/qaBU02bxNdQtGp2j2GyvSCPA4zYVi5df7
G+wbXVdVmOyg1ep8Fl2Vh9/uTzWO21CC+fULM+GOBqxHNRD7NFduGwtOVCW2e/WXLbVKbMx/7qFH
d9b/lIcYTYDc5aVCY/5mpAsdMh7Q/zDUKFyIqyDevj/bnqs0DPtpG6cc1wvwxcwQdYTJh/u9BiDR
+iLShI1pVX6dcmklLfZlIbcBrbw2qOQYx20NOO0epWZppIlvy9MYfVHXX6Jj0RSmceotIM5p6+VY
c2ADYgfPsM6uA7etzc5eqGcBAmvlHopAYKpDnkPmQXsDE4rxVy2MizvezfY/hYPJlTe0TS4acqXc
wgYEPY4FAzXBAFmlrRAU8tERDV3mFwpYKkHckyoC54N0tooYnUeHYWz5ohA7rZUhyqKGe7Tz4did
uUReDfbHEby1P7Yfs8/Hxv8VIjAQmU3PU8IYcgC4p/XnM8aTMCghCFD5CYs0jbyMsv22rwtXns2Z
EDsFr8TC+1FHUM95CtindX3pxUmvfJSKs0lBiua6RCufYd/BvU1mMPHNxYTSme1nYrjwsXLF/D3y
VqduURSIxqoAciSuCRBdmRoi5cCdFciJqtarSDMeYevb4KGgATotIxEofGJUM1XdiePq64f913jH
wzVFW0nkAZaXInK416jL7P/lMKi2NCGrc/vtwfSZvPtVndy/yy5XQq2qM+4VcevoEY1oz+LFI2Am
xrIlVeLV47vLucAre0wJqGtpPswKpI4JJ6c5F5gwtrtCFkeZm+rpM+1CuuJKtXv3dK+ydQPS3J6g
q/N/Fw0VqBW+fg0wLrbwaBoGzZ1SVG5UvqyGa6VVan5MJ3i7DEGifcfsJHwCPrS59Q7CSxa5oSHy
ujPPIKAml36wwC5gV+AblxwUqE+reVD9r0UCVXepwoYA8Csp+pZ5nbmm/I2Z4cGvCX/DYFbvnj6z
Ro2Ua7VE8yalK5BfdLkwsmoVP0zAQRCVnBnavRwjZ2kis217zfpk1XIe/MJl2vfYBgT7LrxfJlf2
VW+yvCmbOZYh3HwsN2Rj0owRuR5HADhd/IoaNKBZY/P0U7OGXmqdksh0nzCjnK0knMO8aUjhp84A
W2PTvOPc+C/IXo39okxQe1t+iCGxhCOle+gXTsFu2jIN4b8+GaE904y0PBd3E/Mp1sJ9rwMFOhV4
A2sPe0bBVXhSg4/uGpqza+RakOLdgj6NkXQL3sOYvSNXhHeaNcCAAc/A2kGqyLPlISRU/6AQFQ/c
cM7vYFEwX0Djor6uA8gIVtzcNJfsCbDIMDF5Rbtf8ruCkKL74Xm9qHdsoQyTNplXpOHx0trAcUPR
UBvLEM+QdQvlBX+M+UA7X73r+iVsXRZ9WB2go5xDzsoY8iQwInJREvdREyj8KnH+0tvrSFAoi29S
1JcU3OB7u/4K77qukRZDnvsnOIVcGUKGuFQKY79gL8NMx7/rK10J/KjYyBiIU68I59ocywa6vPEG
tEIQD1Pb6jcXSWbFQKadTjZ/DSueP0mJRfV1WNSD47qBSCZ7ehDVSgPg2HxV5SljEuZp7yoidt4W
d8qG6oFhddbALgEl07qlPXP6B1/+wKS7DA0an0Sm+KLXcHkHnfQAVzXosEuj3i56q103O0klgdJ7
vNmWoo5gJUGwjfWTKWKxlAef3cfElQEoKYPJ2coqQBngJb/tVTpLSqMPMW1YozLpElDL5KWE1yD7
pA+puPCT/G5cdlI04pPgXMDmQjrn/jaFT/4y7HXDyhYBj62pqNazeNzeeVK/KN4+D6ULI47RgV0c
I1/M/h4i6+CnbbZHeYG36M/vCwEQBoDodn1q6ju61DV7ZFqYN0oZazG/E8BjL9qMpR7nMVojHnJi
MUqgMlDv0V0WEo9Bk4nRWdIfsvbY3dC/JEibk8JXyfcV2DnalPDuJRRw9+eYTv4hmpUSkwA6OIsg
bB5YiAgxx2Y4j734rHs+SvzBIBkNtOVkFW6d0xGqQOUi5a3zajnlVy/O67fKG//Fu3tnxP5oN44p
Mp0KQdtEpOMLWUw2HVFv/OEFCX/fmGVfhS4C0lLqmR7A2qim+vZHMGKEWEIpE4D8JbQeYbU+hU+m
BlRk0w3myBGEcyAWaDYelQgXOsw7lIc4Zbh0gU0mazyy2ACFSuB8BdlBiktKcLmL7/oPqlTj3wtW
ZdqrH68gecQ85F1yEjJGhlpdwm44HsERHCCbm/3JwOu1ooeEBNeI3QDlKNySnLGmjz4YSMyupAQT
wJUBmBGBMmAbfkUgMc/9C1tKubixZLFpwvOiefBekY4JUAuk5Qo5pdqoNR9ovJ8lqjpgwS2Fs20J
TeFZgHolhw7h4ZXWeMLcQq5ecLrYDSAy8zvtGZFTLcWQuGawsXWHLdnxt72TEzIuOqdH5uLaVfXU
1anp/Zil9j/KRSUxPkTOCg8vUlLGMB7iSlfWJQ9zGCuWl5CVgBmiYifZCilOtn8TGk4UIsF4iUS+
QDTMpA9gpb1c9ZlXiH8t7Ny5M+E+bGuC+MPf4PN3Oq+X+R/twsiuU9wKlgS7Wgwueau2UnqRNg1n
wcRXgIpOvNFf/V/jKeWVG+RrLaLdfQ/GYvnO+K0TE+LJp5Fo7ZArxUtd12KYhSInKMD61KiA20MY
PmdHKWV4FRgCuy6uGc/6+UMNOz3Tl+simJQCxtB8gbDJD23HVdXiO9sLMNIqLHkUFA2sCjKRgd6C
e6BuNqRfJeOHyIYxTDa3T274Kt4JK+zr8bsFZjXNFoX4aicHTcBMhD2PX9ayfKKE5WMObh/bA6LB
GnU3Ga66ZHFZmdWJISuZNJ5eAaRsxkx+LLWJNuQxtZ9Lg+hInOEWE7wvabMrYn9PMtrM2X4RuPCd
chCbxCuPWreRi/WWExzevLdiEBX7ij6ikWSDh8aYqJcPAQDAbdYdCPaJ5Kc4Bja+o+ajb/svwxTE
VZIqE8uK6OeGxfWXlcBorBSDjeQsQ1NRAcOssfRCbGhgN7c5E1oxd5vaLdVxdz+fN5cLKD9SdfMy
AYdLP7976cUXu7PPim2JKafVgLuJnK0DZRdsD8Nou1sQa+fheyQEbHs7RmtPvkOLMMDYGzmuwkkh
zP0uCVuo/11fXIjmJDC0DZEDxHZ96CoVsg2qYJP+wzgQexxqenOexDqE0xjapIp+zBlHmGOC/5A0
T+snXNVllf/e9Zz6fRjIkwiv4+4qHvW3WqDjwwUHx0gNLTTGDauHrH26WQcQ7a5wQcBvJafm2njC
aW6o1wzhLZ5olBDiM56TW94LXoHc541i97pOPshUy6NEAVl055EKRj12s3JPXf0GNhGPTPIJcOll
d6uLr1AVPo+IHbBgfqhhQlodmy8dbvuzdLX/NLUWhInltNRyIAB6MZYe6kItMLxtqZ6KqcuPx1Ga
5noBJXxbw0qQkalB8wKvK+w0m38/P63fN5E3AgYZ4LKokZ7PxAGHp8mohM4Bm9kScV27nVbfN2gU
2jvdcjpxF6etnGu77HcmwkSgN3BXjjrt6qhbx6SJ7c4XKy4SPkhXFaZwzDwYYpCLSkopPoN8NrPn
SIE0Z+BMMUyq/iOwOr0ezSjDzoJj88fkWSvtS+1UrhlZA/C+KuHD4LyABCiFUDvIV1hiHcyGY2Yw
yNKx2cl8PN6dvJa+0qFEnqTxcy9OLmhHdZWAmoWjlywxMHKaJOhITZyCBWXqAQT0fP0Pp9LheCql
Y+Nsae+2mLhPKcbf7lX9xvMupb/7r6y3C225iF2dF1Nbak6eutvUzULhBJpecvqU/SAMirRX2LRf
ocsrmAHHGxspIdsKf6u4FRQUW874A5esvP9rRcHtqq2JIlaGUAOE8VxjgdvzNB6SmxhOv7XmA0X1
hvJrP+Iq8Z/FG44bXbLFMjnibYLjtCYwSZ3cJcLy9Cb/PRAB8R7jfVK5dP4wo8pty8ijLnM3bpcL
I/0AgG/lGLfoIZH0YOKClM4+Ru+Kp9TwB7uJKXwyd2bBzxaVHiN5yPoPq825J8zbFV1T1JQ7lmFa
qLOSmtNQImPE3IeaRu5DXcWv8F2kYzgHvjGLPlVgwobTz+ZXYZKxo6LBWmANe3yooA4KvdxSJgzv
APJGlxqBW6ITC6sDAZpqQpAwWRuTsJ5i64aPDVvnif2MJTo3sv0cffwwN13MhsiOJ06h6jDvexwr
RgmAf3Z5yjdFqdwXyXktKPagi0I4fJ3lwHlkkX5W+LuHKmvKD0STOSDcd/JJlD4BCE1WQx92gLLj
bA4DNzzM963jDCHyF0JyeQXZc7z4Mi54WAHzj3772AlED5uio/Y6H/7LW4tnQjESVrrBTHkxYG69
xfQMalWk7WgEoZrohB4hFUCoXAX40FU7M0uGhtEIxomknMbMkSSfUHLVXyPRxqJHpGc0TJ7hwoje
2xp5SPuHxTCcyl7bPDQNCTvzpv9q5KOsiF/W9zLgXCWqcWh0YDxJVTBjNCNS4fG7kMaKdFURJu0E
+tAFi7gtYo+CfvSccbJ7vif/CWxfErpfnbyvYP+SjFspLb/WeJwAU/Yk197rb96MCr7ikIM6mu4P
8B5erreaNaRQrO0dT56tXRosp435Ov4g/UuZUrF9jFQsWxmTdzVnQi6VROM7GQaMsrs17wgzWtvg
H3yxJd0osLzyw9afNPNnkYZ4J7vnVPSj+hHhTiwVaWVbvW6zR08H/4yjYQW4Z+AcS5pZzsgNO/Um
XlseBnlMPk2alA+Nf+KhM5RF/UP+BwWoY7weQOG5i9aF1a0JxnTNju6/RF0WMukE00ryctFab6Wq
r+CN9xEuEB+Z2c3zKSHS/DUIRWx1KW+caK89mfuVAlGQ3TTWYAfyIKSu8PgDNZrXZzR5GI2k5Mu7
xg3dpxvbXMP8BiF0fE4+sPv8n071ZmJWLMEtlGT4zMIbFWXGBSOX5t13LVkHXZBeOPsk1UgasSFH
YENH6XLuVsM5tRyIkC7tirNxUr0MkrdRYdZlU8t0gu19djSc0mYzc4DdDi2GxoAztqaegWk3p9+G
pMhp5Dgwyq48LoqNYhwCHQNFKq7P0EyFv7NOzCD8V/ZOHLLwmQTNmVhqrkKDmMEGy9f+xw7Ojeu3
C3mfGkPjDj/xBA4Jbm6FA8IYxtTJ+ITCxoZyWQCgcNJ7Ys/tb7aB7IjV/S3hFQ7CzvUPGv2olmzL
C9dRTNz1OI6qg4DEaQ/0oaGgwPCHDgvsFhLrmkLzfrutSOYEURJvllJd9TO4Rf32r3XoblScWocL
wYyljF2C6tTRhBXDFzPF2kg1ihn2X1Z3ytjq4/ez1gQYy3tR/ZCmOBJT5ERS6jToBzKpRaQ0YVWx
UkdiSfUBdT5RRnE5JS4fMw3ohbrUvs2Bvq+NSnnX0Ry+y9PNYfQrcEhfFOCzaxhD3XEOGGJdR+WP
NZktA7j03ApXqJ7o2Y3qJdUOQal3iyUYTuVgjZy11RJkFFDimJgcDYYeSdU2ThwpOBxzjb7PZsTu
tSylxROMMF0kXmx2lu9/lhuyJBY+072bVP0ARpp4+0MKnkcqgT3AxwGAVkJ93pwRyIBQXk+IzAZB
W9xxVYubfWvFHsENFWirauip0plj0p1Fawh+yQs193AzJPld7v1OcDffHoBkDHrg2xTha7MfIHQQ
f7eN+jKFYc8IbyLh8g7k1cF8vV2gYUMrDcpPVuETnJtjACWY7eUCj8bIB51+SC3P338Xp9Jjw0z7
GgGHBExPwDBjufFDfxcno+ZXujYkfY1R1sznXP07sBlbgon5By6zosn354Pv3IYEAk6S3rdwGJ+n
cblcMe0vVO6JgYUgbRwP3ueNw4OKlHaCRrkpAo4S84dZGUGZRgZfPBlkVseFn/6apVuHRDPRtgk/
clalGA0yW/1OsKPzhpasrZEJPqo5r3ebhsGynci+8F3YtbwuTyHpMcTGtaERyPGTWulDUOvtVqv4
0+jKpprdUyn1mpbfwBp4AiL6i+hs0sRvaBAkAmSWlcFIXDcg4PQJx8T086DMdnoOv1daOJXPkMDL
P/jUYR47+5j7qThVjPN7CyGgo+o/NkUqG2VrMCBz+DW+w02PH7ZjG/UlIjeV+HAylc85C3QIb3yO
rNDRQKxDczPE/ova8ZViHzeR+XVq85WOAHAVeN8+FTpC4QD1pNFvzdJoeTO9biqRm7DPZf2dQenM
tSm+6jwmS4DTRrxs2OxxznO4bBdXMvYqDbjoJ7G9igT6r0RytuLNC/1K+Oiz/rbicshretXnHSuE
VMAv50PFsdmC/DtwY+cdsPDfKwp93F1fresqUiwC8dztnHRfY637cwVXdq2k6imckmRoON7oOpJZ
uW4F8nlAYjvYy2O5srYY5V0p6wOnSrDOFN508/jeLLy4yXnXBDXcbciDk/aVE/hNXpIl0Z6rl2Wh
7HwPDVlzcqdq6EoBXIO+wU5BgfJd0NjquNBMnIeyYEcAXV6Go//xjWYZYsDGMB7MA0L2SQxouO+f
IgmZ3pFqtNrdBDCNAfKcPLbVsa8dWV1yWSmt+UArJ2XzEtVcy72YFzSLdbXcexet0awEbIY9JfVw
2yq1qpCrpFXc8WzuPWVUorHrf6GARUR71AS/0bZjg6A+F0IdEDldMnbLDNPyYrNFRCdElFq14UKx
rrvUQitTJWND8KWQVF3y/mBiTqhEf2i45rnKjPSvtjq8xGRDUR4caODh3+EviZMqEeErZj8+0T7S
Ox86QONrsO9t775CCGzKRtaSAi6obmej+hxwHXbn81esIqws4Bh/42wlgsKwAUrG0VEo/5ZLCBsp
mZ5c45IoVVZ5WuYiW3TNv6h/QGSm6m1CaamTf6sZn8PWiNBbR3VCF15rVvAql/4QnE55ghKmQvob
bmxI+uDO/CwsodR0AclBFkhUdJu5YL4ShJYgmrWWQFjM1sGyD7FRKLxpjAmqutgtOXPc+z4PRvdH
9GBgRmGK2oBiwuUGm0UpHSx/njEK3IGDRM2AFfOI8ZoNTmi3HaEc6vrirYbS2kAtGJw8kzNMS7Pl
EEzE46+IhdF++BZS/DZAh3my/QPaBUYyPV1JJZlfQHRnsy8FKvQmMuglhob5xsrs+tZrs/961bq2
bW9EPtm+uURpQPYjQai4aINznrALLCUAkToaAe5ZmFD8mpdFxPgaoT7uu6QH4aZwzu7Ud59yKs5H
14K6byiNuiLdwAk1gf8jaqp+uXHWNmLBt64V0ozvoeqIRKOOx6yWDjllE77slM+dlej1LFDrEicu
cu/y4a331GqDL5rWUqBrrG5d+ysxup+M3hG6LQ0FpUDil6FGMtd5l5vf3gnMySYQ7sF9iPLQCH0b
nTb8cwPzb3spfweWMghpNs9mqsLeTSzD0LlOZQjnj3CTMuLA0H3uPLjpH8c+CNznvh6AdWmvaKmD
82n3NUkKNklRviI3znyiw5gB/k4ia0iCsJvaWlLRBUeD2xyPHPt4iTLvS+150IpbuoqpqjWacA6/
xzBc6crHekwcJcryo9Jc2TuQWqLUwScTvXf6UZuUSLwgleAHo4Y23tIoOOzFwniRaEEcbjk6Thqu
WZwBwOAm3LOUosNftndOPgGkTpnHnL987B5ybq1nC+5ul5HLMq6BFRUMTqk/JnEyJgF30Gf5Kn4s
sjjgRZU+E1JgEi6bdNOXqeNITVz3LkU012DCMpEf9G/LVq6uTzTcRjdyj4gIoSyeQ5y27T5HXoGg
tTZn+vrELmY0Tp4yWulPHxTO7Kij/ifK/tB68OILyHlrT/oJp4aQUBml6kw3+u7JA3QUXss4TVmW
KHlEHE60p5wV7YqhdzNzk4xjr/p2EyknwkgHRycitwbcfZqUcMRXBHsBr34kRWhk3vChPK3ADETF
6G0pr2mJSqruMe07z6tLKywGwiIQVUVfxZcMj+Qiaz8/IiuS0xz/Qscl0vxY4OodMaOLL32lTO5X
kh/pPMqTbw+SLecdSSVqwu7VixAGB4+kqtQMc0hQ+n4Ho6IQeS0l5nRAZzOLrooh6WNFnvevwdMi
c3uweMZtaS8J4wXLCdbaH9BaViGMzkUfaHIrefO1awDCNRY3SuK7Ns9w11bTTIXHA8+Ng5Y7czbq
OSjqq/2i+JVJ2+wRdyEJS8bqsJ6SkQj8h6kFd040/RiM1Zal1o2fAMgzNq0wpmw4hj9PzlWc3hTk
Jgk+aqqKU/7VewGR01GPu03ElqKSS/KdUsejwtP/rcrdbTjcP+oT0HRFFIiKooGpn9Ozk14cud+k
uaFHDQaVoOspmbBN9BXA2j52wfyWZ0rZg3vZmT6EcWGer0/pO2X06EsaKm3P0WoS21X6RDXp70zZ
+zNIJrjza4+5+Gr6XQQ4qNbPohftoQSBx/E6t5SQrPp4nGhgW1MYamlwfLFiFt/cGpK9x93Qkuz9
UOUHfKFWfnIXzhCaUAFZZS4lsXen+q5OFxPcnMy400Uygt1FpVVQ3oJiK4V9dMpsXVNt3wKqiPRQ
TDUBcOw+esJMLbUtRYoXFljgVTtfPpSqnJNa/5oPvq+nN8+5SK/hnjAEaunYENrxTSLXR1XdbiTs
b6VY+Vnzo5RFrNI6qPGZasMr1ipbhxNLi3KJKodTjQyBvqNv3BXTBSmtTFT0/D3Qk7GljX6Gp969
igPzUx1uUCOrLs84in8HAW1TMfwKrtaocZ9EKSEZASWEDDkGLW6kPSLlk4aWaZtPaoonhIrs9ee/
YB0xg5aHUaopwDCGpsXu8iGzAdFDLjVwsQwFJSQsyi2SgCJL5qfZ69RnVWbWT/ZJfL90iLQUZKSE
oDCrTdba/SiMQWQm0dELLGN43pAmm/ie72E8ZFW7JeKJ7gtD2A3QrIcB3pX3SD4kGwA12mrr0aGK
9Kq7W/qkcxQC/XAbIUanhh5v3XHGT7FVM2JWA9M0o6eWCB4xtUVXg32PumPHdIuM1d8bKOiAFpVr
E+mTEijB46xFYqQJ3s3yTfY9sNDxJEUfnVS1x9fA9b0ZekQUEuLhYvnYT0gefk9UkEGIqZfMZL9Q
0qte0XIiuRg/xBwrkD9RlCzTih11iqL0tSsa0VU2teQxCTl9Oulk/1o4PhJA3wlDEaV8Go3uVizm
Di4LhWlXuuR6XcYZ2PAE5on3Q27T17DW0Q2vYD40W0kP/FhD9B0dtkZPQS46tXJLcqJoQ/VwV+iF
34HSCZmRZlQFwFbnQTGC/WLU8bGokJAMxFPIePdqvoI1N1fvO6nLC96Ttpa86x7ek7BoofS6VtIQ
9SQhYFaIj8ci0+fWpxgYq6BLTaSDtyf33BUzL8fu+VGVXafFDzWg0kAkKWruyQk/9ITIAWVDJtbq
o6+Z/vhCQPzSPZt45G3F7Mdzi84D+by1VIBEHwuKxay1VAJeMjHFbWEpbpxQT9e2iVeM3P/Gq2l8
scCSQ49sPYIUFcLAP5miyvwzpVsarLdP01LD2LD9hE61q+LZi/hOr+lAhgRpaM3B0n0K+RGtwSMM
HMJXJnUuf3mWLPhTN0Xonifm9YN8BLOkjP2qlShrtl1JDc616I4Ukf+fDKdwCfEPGvWYtY6TVqrS
e33PVrvOasPUkS8foG4MwvK7DRXTiBSqKeJoPoW71M9g0qVCQ2iHyzDT3TdbxsDklf7QdnFaIxrh
v0cqUNaIdv5cs/nJrwbN3TSZs4TBzKSZo7eTndXT3qd7IJzJ1Vesg+8Camp0YYuGZyZSQKjDZk2D
C+0/Qz9aCTZc27mn4WzfRwLhk8+bFzkUr5E+I4yVycUUqa+UZWeerqyfMIeTJUlCBFd6tHf899Nf
jIKYn0EWRoILXe3SE5VCywch9PK51jjwDOmn2qRBwkcW5CrLHKcjzIAO5KswMuazLA9GmvgJSgaK
kBsLbWzZ5Yz5/Vm8+MIGVDHrUuqBZN+/G/xBStgEf40ynbg5j9a6yZGd+mTKGhaHNgvpDgfp9Oef
0QUFrdYrbmeEKc+zBNMVa6c+FHfe+gS5C8ZpQ+IaA1QuuTGlNPPFc6SUpN3bm/8fGem67LWW1eHP
QGeKqXuz02D4BH+4FlaGWoTNg9xPiwZybJI2CuBcfz4tbz+Vf8+NQzkq1caBhC+734L2gIHa4gN8
AzV96PfKFckNr8j1EIJPPBEUV35bcZumBFSVX10s3GaZwruNgiNxdetg1gdwJn2waND3zyq0Mmuo
zaDoYIQYZq1Ab4cQAJrMrDRXe0czFSJBE+jYYXxj4BXqe18reZDpj+AeiYv8nthX42VERo1A8NmO
9wD2PIvNW8aaTeJ0Kr2X6/Xi1L1gtCtlN2BPotTX9WxQtcnPz5iKxuuA2m7oxF6UYMfpuUa/7NhG
gzRk7qLV23QblfIYV2aPwoDC5cD0TeyKsieyZbj/13T9k9KDCzAVSM8xRaGO8n6cYrLb0OEVrNIQ
ceElVwLNfSMwVOmI/vLSNrRi5ypyvp4ul/KfMvWr1YqW68KK2W+Jfua7ucw1W944wIcY6A+Xiu/N
Nofpvy4OjhfwzgjTJXwl7bE8Jc5sXH6uE4VMa5PCdAjkdm90sUha3+uijuGHgDTd4wtM2YKBM/FS
7FfLKo+J6xoQFnGYpaOj44YSoV/lfUJNzA7K5bXU5akr6ZKvkk7kz6EfVnYRkbIR1h1q9gzuFA9U
mreiq7Us4nHc5vhF1OGCo+Oz8qC+BqOTqD50gC9G0KBJnRl2ZQi1zOOGv3Iyv3TLBxQYOfJhrpFf
JFBcyZ/r/qws8cQGf0HA5bw0TzR/UU9s8vnerPftQX0C8YSSxTzoIUhBD/oLvZdjGoV7N4bWjBWC
0hco8JUQzGKxMNhRmc4aPpxTtI9nz8W3F6ISzlQaekwWckKmVah7pnd+VVJ737H41ck3rjMYx824
M/6Ei1foFAjWJkKtDvj4Ojez/ixVmazgxASxnYRovjkLzsA7DKfjLWY8wrnl7ppUQU6GSQZGELU5
7XxZluWhgUWnZg6VlZZGwvHja7gYNu3YqVxaysb8uori+zRSUrY1JFDx+HwsjZpwsuvw8ppEMRrZ
HViIgCTn/m40Ham+1K1PEkZjLs4dm3a5OpJjbeYVHu1FQHSkCoiPPqXxtDxR3JMbrfZg59deYHx1
wywB6Hb1oNHQb7/wQjgzyta7V7goyzbsCwTsHBHvzOy5FcKHPx21mBbMbOz49Fs1m/yOXreTcCCM
47pI/KpkTXr57q6UFCQqNrl0+DpF8vSt7cny9R/tZNGygeZ4WA719pCa3zGD20F9czFJzGNXywJl
fBF8WXqmYX3acHYDGyxxDu4l+NfbankA5xhpj3cyrSFexr/hHKhGanAqE2DVelHCaideWxDceRjj
Vo0IvH5drRE/PdVHf8toGZnWIflUC3WlruQEc4aY8Em9Jrp4td73XxOtIZqOBAZuZRbH8fwxAmv9
g9FHB7alpiV9rK6tAaiYhYzQdoKxDBjo9nEdrO7phet5Ud583XztzyTBfuchFR7xgBQhX8IPdsSF
AYIqaiJOr4r/AkpeoKScwKp3V7m9qekGosa7AtaXkM2ka/sXEz1THY5epMKasKjVnS8pEqzOt0Nf
ap9w8vWC80TE0Ezl7cv9u8wOLdzb5de+lDjuTE2LEyl4u6qMHHFDEJIXWguXyGW6h2ON1e70ez3/
mxGyabmHLDMnmBkdVVuzJ4FrqZ1xUtgpN8o3JfeZserGq/hDm6+rfS4Zr3qupOgQ+GAZ5Vbm2mto
KMoklEncHiXGi88kSaPn/pkKlVnXDGVrcSMmVTu92T6qAwS19jjCoZBSXsC1xy9TGaF7Z1HErIH9
aUK0fgrJWdyaUXywhVB5Z/wbPLO6dN5qeY1MR77+agvNztNBCVveoXOlMnNwmm+jfKi6ht+nOurb
VBytvNgt1NUAXhqhlmFF/WizufPaTwEP+Op3ErXbp6JbkTwyGrv8EHLvCgCFkVJoOJ5up+DMepMv
n4GttBJm+ET7pWJu8PDPDDmwoCVoIXiu3DK2BV/NYNbPfE24BgJdZDTJ/pQlqmOgf8m/ax+nPSqd
erdiShWiHym2UfoJAnhl1b43sNuXSiEDFpoxDHqWGI7f/vZn+VDc80T2hPh0XPtIOU1DClv6wC7c
Y2Lm3rWvMkQo2Hg0V4ClwPK+FCz3mWP5C4vRNqHpDVjqGSb2ED8reEGAANbkBBUPBW6qADZNs/XR
Hjrs6y2RRh5X1A8eYthR2C7SoZGzmKY5wMgtACFEkgphCzPGvKbcqbGTZ+xK33AGmMb2xbF4spuH
SfzUeGaN+GFc6WBCOW6a7zP3goAS1ESughI+hz0FTgNrC9UayaJnKGfUENeMELJWqYlfYE2p3XfM
Zorh5g8OIw8Ebl+QMuAeklWi9MJGXrtgHnvm+2Mh+cI3YvFFDX0XIMh1ZxHktDvyxwojTZYNQZOT
ah0rsQukWxUF60kZNPVI0pFqEf5r9bWEYvofaZqpOpPBdFH0O+DlegJV3OoKNJY9uLpjY3lsxSSH
KoV0eR6mAvnVdeNDuRhZsNq2ga+5wcw8UPnCdEwELEC/wJDC5L6V3vAwQEMrPfkS5LbGDp1lVEYM
y5cJy/M4t7axBzyBGHL/44+O0nr4hFI53MpOAPX+sD4d7EVrf7kEXpDW2GtwIWG8c0fFmY+Gx/aQ
nTHYb6emaBuLSCTgqn/XyOzY1bzXRm454WpxG5ThMxxQQFbHXyfsVo7GuXxU/fcCYwT4U+Dlm3iM
oSEMYrrFOfQLdqXJkd5rcQ3B0Ip4LlD5FwF+W7008P6yrei8kJhFd2t3Bz0WWBXNie4MobpzcTpB
4zBWhQ2xO3qgNnCpHBBAslZbEG6Tj0rep52sFNTQx5czGwwxpfXV51HShDI8pIjGNZ0qqQ+B2g7Y
CGcMqcM17qZ02pMGfSrxG+AqR1mamks81/dKP4lU9GwdGjfLLEkFyii3Ufu6pQunuguePI7vnpNG
Fkc60jhnCoNsRjZzT+EEwGHHM95ISWaajvty4MBlO8aSKIndyHI+k3X35xC/DYmhDS3laVXvzJsF
Ay/whU3uY7qgY6rXFbGlA/hNk1I5W76j5m4C4pmxs0O/QoLmcU9OxK5jbGSjfkcc5nJY/TqwhGau
2E2zTOU0sxOy6ikk8YEPhCBQMtujuKW7qe/14zA4h6ad0zPV9F4UZnnx94J1WFI9cPmE5pGBqnS/
XHAwE0T31ihCib7c39nqFrJQiJt7UGHF8GmIXjCFZ1TJve727SIdl4rKbChj9RtXfiPHt7gfgmAf
eTajSSnLmRVTfgn+U4aFX6oFDzAcv4DCpaDyQuLe+rdYBSOrDC+geI15jWRJi1lku7X6uE0TEGAH
0DXV8z1HpYD4ImcE+2suqnSR/dA1c46EmbxXVFi3cUFDO3m0WkPYTQfUBc+CyaYMgMEzAKdOUkms
Q9JvM9Ck5liE/lFEFj1ZHDa6ZpPvIk4d/IxpO8/taduq2Kg3L9qhsS9NgAQbmfuDYIICPyluIxf3
3vfzND9BxGHtHJRPlgYkJeSto8aTXRQfV9JBv/dl/I6qrM7BBdCsL1L3yp9Naeb1frbvIX91B9jp
y2WU+Hut3e8mixgwl7E2oZtAoxK+CeooI45BBWGYlSBnoyVp/lPVPpkLD4Pm3SyJfSLrpbYClyxc
72WsvjFYqF6m0DPdLR95c1DsEbx9SCAsXbOBBjy4+T9P5nGf+MrAEWwAVm9x2o/eiheTXWQHHSMZ
cknztPIW5sfGYEuANs5+WJAPUaeiOQZakPOosQzi0zXSs9/oePhs4QTAkMRRvmXBiklB9IrZT13S
5ZgMJqo7UFyDJ9Q5kTfpq0/H/Iq2R+HFpjkX2PfuTg9+O9MWasm0fjOXdS/M6sWNkQF1BgZwJG2a
JtJd19cBkg7UxFJVL3hzNjIrdloVCbg8nztaCRybGQBcU2wPLR4S5820ivHIIE4DxepdfJ/k5Ybb
hj+/Rhg+4eZGjTEfMbP8pbHzbMoCEYDoNE1ZvHJRSFTnnpXovZUOEthuyOQrRR6DhfTOQ2bqcYaM
9X7MRuOgJUceY3Cn1sBN/OK+sm0IYm0oCj32mTZL9xHB5DSiF8ZPPR9zP4jQzDR9YKf7RPR5cLGg
CbM0i4e5T/LIFxJ6JlPJYNtqY12dss2J5PJRRpd7rq/aS3AIRhZWtEPY8zyQtmYDFJJ4S1SXoqjm
GREctbZaFduwpNB+/lxV9oz0mmQN2zlQtJqkLDYEIYyYG7mX+shAfQokEVG5zhWYLoR6w0jFi8wG
zKtR2+u7gx7yaMyHQPdpGZq5fnMniRezjBwSnUSvGG9YvM7lkIR1ccETZUqxzK8dXsiOYpwYxSrU
mxxyyo7BtYniZ/T0qK2KgOutHYha76C58fbKsnALlP38ttDmG6qymFLGcmWrPl/aw2f4Tt8cZRm3
dj81kcsHEVo1QDXpokw1WWqzSr96fJ1ANzme5PfxS945SuTNrGg/TVnVVXcecbSlD5bBYw3SJBwQ
p8dM6r3+zPbsz0LVW4qvN9wt6kYr8KG3OsZTJTjZTMk7+Mgy6BRblADoMsXcj/l6ut2877RFjS5c
yRxXWjGTjdeumDQoEYNb+yREbwshgBi8t0Up5A/Sm6cy/l9pAsIXyUvWfZgCa6nr+KZ2M5j0xswE
3AVnHFET9HWnvzzEhgLVq0VSVHKudDBVtFs5nC3oFSFM84mQ9/+kqQNl5CmkQxNw1m353kiXE6pB
qkHI9Sw78FJQs6npx3nKjpfTVfe2MNl3DKEdLLvRBs9njuFcZ4bBdTUwjlygYFbGLmOZKpsCLpCW
5zf6Q3hm2v7+/fFIIsRbgp7+f9n4H5C5g9U0zwU9FDxMqouiRlnG5BO3OYJwAIWRGwWen1wEu6IC
uFCIOjuToIzDLqSaHD7md2kC/l5vewFJaKCQ46YXLTrEFHzykUaU/sCb4Ntd5K3Eu9QW9NXfYdkA
5SMR42hhmHbF7gkTCGC/SJmRyBDj0d8rRxZI0gWAx6GqHYKbQ0guJM/melpgd7XyAz6jGzQFLkjE
+tq7sIlXeh5fNJN1lP8qqzh2SzCG90WJAE8kDK9WpjGx0WXy9tYpa5q/Cnz7zKRRoUx+FR1cKRUs
xJhivmbQNDYcc/Cn19g011kBVh9IHlLAHGYuVfa+JOLwtB0HITfTt+eUycMUSYxAPEDRqLQ+IrWF
DK2+IX9GuqPmfiYOPd2R5I2wuj0/54AY/7O58vhsEXGUC076qOBdaIxrboVdyK8SZTLo7SN/+fBZ
j8JuJdS8mSIj6al9B5xDHQrRqlx/pJKf0v3nZyEHCjFixYy+GqeuFMTa3X4B5DoXyLXkeVZMyC27
YbmiujNnqdT7t1+mxu+JiR3f5Nw/psVifxWa/NFCqwifSbjq0qmW4c1bhN51/2toiCKT2tqgiwdv
SYvUUwxoCbVn/3rbNk5AWoHzVZcwfAXMBnRxwga22UWosgsFmCsnIvOH8b1BHcC/LmT/nq5DbJC7
tqdKDNJekxJiXCHXV/AvcZrARqFXBeq42ZR4g2pMdLorpfKERgJ2Et77qmW0BYc8jz1XXTD+hW0e
QHmhYRyo08pbJQO8Vf9lRPTtcI7B7SWZ1n+RPKYcjnjvIJnqZOQ8lRY1GJV4p+jFv+6EM6CZ/iOE
L91psAz7WQUEGXzYMx6gK7j5T8Ny2uMcEiT1Ck+aQJyO1N/G6hLq6B0jM9zR3njj61B4YL82bwv6
JiBH7BajpEMQfFsE1isU7GDmrzhlTuC+k4rb+/UGxNcRLck88HHVxhbjV1npK6MBtadz2kP13TRj
LhHVqBr7igpztvqnwVSpKxY/wn67A7FoNLimoVAODw94sOuyKNgPI5iWm9FlXzmWy25A69vi9xvF
nvHq/kaFdrukzpeEhBg5rv+N0zI92bUb+b1aAzgGqGaP061J1ulCnG7Hn/cR+nCX2Q6rrs85eHHT
4DvN87FK4XFCqDvTEQQz/5qM2RM1nQU5anWCZ5CjM0StUW5dZyrU22zJcOlwW4WdYppWmYHRYVlT
PlA6T7XhvHiNdxoAt5Hi1NBjFMwh52Mtcg1Ah9L79/WXHPLmW4CjZuA3Mg8gjdaYdtad7DbSkPXD
4e03KpuqPnisExPIOQEWO1tdLgwoHimNqE91EgOMm2KYsKJbORzU4eALfZM92aZIyQE2rPrR+1Pp
sCMWwzNqubSHCmi/w6EYvul3PXzPyFLHzTFrNTwfkusCAj5x52oGSQ9vn86a2t0vLF94sIIru74m
8IhLHJOQIbeaY6kclyps3QJJ/qY5O2Bfs4SlR+EK204H1Agu0aY12KiqEuciAENoV+PC2yWTo5yF
i60hfWvFIWUk09LhX1e9bqYLxuNNJqxSkUfsb3A15A7kKS6Z1UannxHdEb+3Z6H8MK5768MuI53W
7m8ZZy4WvaBt1lfh/5f4HEIMwX0EGaoiajNr6RN8dF6NbWere/kI/mthjYqBilyqSzIYHzEKX8YF
bVRB9zAfwznbeklkcMgULqPnjtEvjnVWofK3EvXLNWJLyFTmJU3PRGL310vEuQq7AYRmjVuxGW43
QcCDQnJIwhvf5m5iAF/qRivvw1S9t670QZVQpanhtocpJEidxCh5ZF68CwGUZmPkMYOXw/0zsgos
QekX5XImKcJgLWWKjB8AuuDe2txQqeEqaKzCwf21oYyUvvSr0xRXgpLDEd0suErhz9gLYae+b94A
Apgo8enit8N9pFkisDulLCXBAFhw6sY/k1+MI3h1hCYpGrNWFa6vja2fUXroVz5NJL6nNHy69cJD
XOPRbjK6YVx79iwI+F73UZaWhn3qFx1jxoTMUVn8xEmt4NWv8Lbh/nY/0RFCD6E7otGXhnXDNkFF
yYqC+lcO9QHBwtX7i7OUMBCfVOyylQhppJlreW0i6KHBcm7ZBrT7OOltrRlFu2CCNu9KnhI91uN1
gIoXOWae4EcUp5OoyBK7SqzlE68oPNW/UUa6pjqOZKZ3taEKmM6EVu/GAjrsGopU6IIS/HEwIDYo
fA/9DhxvlWf5d7ZGByyfC0oRun0qlAuEDNvovQqRl9OVEcpyvwWWKROoTKvd1wrFJGBIKkbLg4Fw
Y/BAMF0LzlzK2fhW8M+yq6FhllFKHvYajiwjRoiwyG9mRBNLvsFlsMy+1ANuCNm1ZquWmDxrXNDq
HvOfoGRIOzQDDcXs1kllvziXtEQ4MqBKZIPaA8+oo7OL+ORYTpbJO7r16eFN/G0EKyL3mb32U9AR
DkpR6WCidsqRJZpBxPqk6NfgWbj8+sT2MYrSVEnXCFAxezNBD4ZoWKrKgl77ovV4xOWRud3kQuyS
xjzV7pVStaPV8A1+sCLqTOdC+fdpldPcR4fUuAL2unJHPZUaPL6MGsrer1hLFD33VTtFYihKizMX
CSpsdI/SKjW8PaKaSXuU9D6MrcjTAbdfxWlcQJfDXF2jlo1Zfm66bJGJ61eZGdwZiG3i+hIMMbjN
4RSjGqkxMGm2oGbmfdYD7DjqnKVs6qjiBwU3dw9nL1KhwHixQfcXYa4GBzIIkLLQ5xPTAhCWrjnU
nIibCjDX96ws10YA/wApimnxRt2xiLR3S41C/Ehz/RnimEQCeFSqV6VaqoN8um8KexCuky5nz4v/
p+sAGJUApTaU0fz0EHYjZ7r31oaY0KwYWCuB4+gXpNHYUUBR+HZmL+pt3H9Vqggq3f7xUYN0RgoW
1aQP5aZHucww92v9+vw45Ja9ugwkPpJXm0lYvmxgWyGMuOaVlKkCu397IVWBmGx9eKgDJ5d1s5cK
h/9fptcAJK2oDzfudorUS1f+wVxyFAXKYeWGiP9TkIESWHApmATNtdN4ZPIvBLzz8b8Wi5asM6Wp
bzql7tGl0MyNak7YHQ95b4MSL3Ntm7ajhn1LJGIvzTPJ9D3VcETKdTDhxIXb9e+r4zP5YJOpgAS2
R2cJAbF4FGP47vdSn6tE+usj3igDkf/cmbqx86+bHNuEHSWOmI6cQbBNxc1ZpMcqjLYOTd1sHzJE
vEl90andwv6FhmK2l13Sy8P4LXsuNYHW7b7Taz1VfXc1k1JZnRcKgipe6t2M5v0hTPD4v6Vr0YiB
ICAQSMNVWNvjuz5vSeMxdIDPQSDtSWURvWRt32xY2zXjOjjx+CC69qXFhtgdPsu6Nj8zqC0uiuWB
Ns2VZl0WHwEjOheUMQAiNqCJXOVgIuH4IXUeBrhNTVKXijWYBCbaZGq7zLPxLA9A71HeeNKA52K1
nyE31/wOIsYzl4GxfaKnl/sv42IadhsBvQ5JYFqLzVXB/H6r0N2C98ZHr17jKFGh5TLUr/lH6QFT
4TluNk2ToFz8KBuirl7ueZutPaXdVG/AXOJUX8hGdbBj06WnWsjJWLQAkl0e7p4O5KXM4XUURYNb
rv9p5mZ4DMySGUJMSEIn62jqIEC6upCSpfItVyc+mMM3ktva4vpS86bB0Ut76WMuHgK7BpomrpFC
MuX1X60BMRM8fdRNAGMzD6+GAF1W9fidpNFxwCkqXZKEQAYC895lGLAzR4xWB0lzOZLFELhaVuuz
ug+8YWAm/L1jNOqzbXk8jL0SmpiEDKueifHsYcVFVmIU5RNpVMhE8octuN21zLJTxE/zKiRRbJVu
IglpeUJYYUzk9eLO5csx4ud4sxBoSVS4vdA4K89lH+SBgOiCSiIYmyVMsiacz5i4R4UC4P2Q1S8w
8Vx+QDKsnfD3joO8f+dKW+4aO4lJpqhnnMx9IFY9v4+BgAKlvTFPT3YWPLPNgLgLJiu6aOUrLCDR
2uAAI7Ad7Nhd+zDQXtQIe3E89UpxCWRQVDPOyp4trLqXDcdAJffo4YJYHZQ2wgXieb02v66SuISr
p3NUVT9Q3wcOwPlD+lB3kDFERRmTInQncmaGs7NIwHmaChgBUx2HDP79JYLf8oWK8I1ZcYauanks
ptCCoTaNXXDqCogDRBoKph8v5g+zcAZ8N8f1RtiUc+YxMKxxZV9LywE4CpUoMFUelHz7r+scUvZV
deIil8O5KoVgylcD9nvDtVo3UijOG7uzSu7ooPDiR4ouvJjg+3v1VLoyIK/KwWpU5YhhWrIPj+c8
9oogt2kk0K+I5+JohKDXGrC3HgSsFJoANhNSRevBjWhyAQzeDhA+cb+ZW5MV2m3vPR2kGahw6zTY
d9AQieTSiHuQzEyMar709dEajv0QZvNwy5rBy7Gwe58bp1WQeP78QyjxOOLSTXlimQ5oUZxVvyR+
IpFtG1RkSg/eX/sFbndwXpsIeI35HWnsfAjMpm+bmDfECHEpaDCT8hK3PTB57GgNFbyrHj7/rzEH
zMBmR02FUc+M0j8jIOS/aqwWp7AgC4MjCX58kXkz7ZYLHwwaRzAgGuR4Ec2hADzw9K3LB85KBMDA
AlhCp8bJ8+5J++DoccgNb8R/jZY1kIjomzLtg9oKucMwgQR767B8aSefnuw94jA8kDzJSiGE8LmQ
Wx8pguDhQtBH0OZ8OJD0mEmdPcGbUt733t3qOdgEJKw+cyn8WYpl0PDV1FvpRXv8PUDXGfrHzyxl
/lzBR5QOMmK2vgALUIesfZ2qGB03/XH/Q9EPx3auTXA1RWkYJVFNlTYxIcco5tLKjSwxjaioY8sR
+0uMWOu3dgX3wbR2Yd0Lq3cX3cLY0s3sbap6dp/JjDeLaIqMbOLzcUnYvaAmvBnEjslImlRQkE0L
SlTbpErZliZROUly15Tbxht+Axa+sKqEjpZAJyTyrBmD/pNCL+AK0lownnFYbihUPp8wbR6Xsd9u
CzXYg7CfaN9WrB8CBY53OU7thIRMwfOVNiyqGmtkj2t5y68Mvt64K6TwcO94fY5ipzjObS6Y9z0B
pqlBpXYCWV0ijKK5f/WXZD/9T47yblpN0IQSqBu7+eCq5FuuIK52+PEpugPBrqtZwgVQmdRK/Ql1
GTqr+SgpDmUafxk1pPuL5FGltOwfZrX570TgxubBoh2PtLyDcs+B8XLzQxQScEQH47G8JT4JTPiE
fJc6rYGXRZgtdlkFxAm/r5jkxfNBq/newUoG95DhsUzEj6+2Hcf7ray17EyAGbOIe35xIieQ8MLt
NUVKPsUZiibc3bVqdwE1zeGso/QSsRoms3yjVq6EN0cdm/xFAOzEZrsJW/2it7qHBH9SnJtojxDF
C6s306cox3MeYPV9Aixu6RnJFOn3LD99cpDRLetAcgzmicl1NS2ifZVdSjDhwKS+W4T7veygg45O
GwdNGG6CG/STW1nt6mBZkJxNnKTwnliEJgYmiWGiRuQZNVZzhsktl3lnbZNW5X31HCo9zkOq3Pqk
k2Af9hZo24MmTRttpus+mGTVqMZ/Xhl8CzNBSS8Xien93BEMQZKWDOPfBsInQFGJyszsn1+clEde
L1Bmd2c2BbHz7K+mn1M1lW2O87A45Q1P9Hn9qb30GqBiXIIfP1G6aP+7ylVpl89r80hx20bmau/T
hsQ96lIw8VT9pR0Q6K0Gg2+TF9nFRIvdk36vroWC65sFldDbTfeZc+/V3xVqAKEnh3HajjuFQXTs
LmdeI0FoZzJj2Rfq7gVFlL7EneSodeJTTCcHgpxBaCjZMvm1npHvKkgFj4Iie40Irv/YbVOMqwGy
28obwajMztSVFJHwLseeJMpjfF/SxtIoG5nG/vEsGj2xIzsj8WVkTZKE8L6Yl7FrL0kHt+wmIK+M
huny8FLcI4DeJdLJ5HqAxbjYmpOlZgAF2NKcANBUn8WFE+ka0AngGu5kHcScPfqWltGs0P/138cd
5UQIzI86k+yizI1iP5H1BN3ecOmxQ3wwOrLKorgpEq1RgYMIDx8N6lCI3ZAnuDw4RcSPoF3zTgwW
9EHzbF68c6E8CRwnOT1HIOWmDo7+g+0JDkiyVGHEUE8fgmib6MH88Su057YQrqdJIhN3f0Mjp7nC
ODeppjNUEcKlIjpPUEyvzGtlCadBpR49ca2n0oPkZ4M4yVlCg8MXiP6hPySzOuwN/RX5eAa22lLC
bPtKY3/AVGtpomesGYi92D7+KQDaXyUqNz39KER672SZ1p3VhVVQ4dGy1TAMOc2D2Jcxrb/R5NLp
LrXP7SjEqxU9ximLycfOIvk7jAqKw8aR6GMHlsxI7RjD0pPKpArKyHB2jpT37PiLiY/kY3nErITy
ild/v1b1PrXrZ29ApQIJxqhPTbN6oZzlUBt/r/u2mjV3LQ0V/aZsiA78dXcJ//wU8D6awXqBzFwZ
gb3J7G2gArWEIMNx5xWG4dbD0yy211kHQPC5DwqInJt2YNXzfu+GkyMbih7Hpics2yrSHdXpL83T
ncHNOINBFgaQlLSgoZfrPTVk1ZICUzFnb669hD4zMFoG5F+M9FvCpyOi1MbJvUehvMepyF9i33j4
a/2eItcK257JFXh4ChYvcpr1qizkOM6Gn6z0zf+6FABytEAQYAqtvdEV0iAwxuJRhmTrxINMgJXR
4qhL9ajDKhlmhIshgROfDgZDTHyjKhKp5tfSl0ehW/Fh1+92VPBYtTywg009RG60b1wLb2GNYsd7
hqo6nZhpmtaYTrgPetkX3HQVoeHb7iD+p35fizKKgIGmPwmT6rznKTxUjtqGCdAXC/irYCQsCWt+
J1TR/qGYdwe0AzI64ULAQQ907UrRljaoIuP5f5keVMSBtl0GbN8/jAEUmb+oWM8RWjYpuCL8A36k
a+xUzJ8t7PADPsFWN5UWrzoZM0wijms95VXIWyxucKuTRyvJSPIfF0MVA+4Avgdn8vGCDO70wNCN
FCjQXr9DNzuPapt+nlW3u0gffZsgXbEFIIS1WhDn6PATg9cVOiQTAaMVp6801qoVVy9TJiDebSp9
Ch3mPr2H7M44pk9aT/XCG4/xY2LEWmZ8B16eL9T+17iP87sktTRr2x2etlHcgS7ofPDeZs1CUqAx
u0RQAGxiSmbFl63s9YpB7Yc1PTzf/8vzl1Kc6prCgcdeBS7SWnwzDXDOqC5Z6OHLxt9kGGA2SN7d
vKfRzxH2YFD1py2sLJUATSzyVZA7+1UYvaipmPdSHRJN6Dk6bgNGzpxrtPuSyU4nnsU4oy0WZHCD
yrCl3WirY/ZQEw2N6Fdj0Vrd8TGybpCMlN42AxgqaSWr0RQcdc9sb7UsZa4UenG0nqsL80NctzdD
IYyNKtZgleSGZTo8Jq+piY6+eeh/3v0LO8YwuaQjOCnCiXbFIcocxuUBYdfbW1eujCUAk/umni1C
KKU8H5jRFs0egN0/XHpWxfomkcpbQmxKMexGM2Kp6nDrdIHFHl9IyWmHIv2gfNF9j+d2z/BSGzO+
rT4ZbMhhNOHjDLYznt1g+6LcbS/eS0uXvQLVImq9cOHUV1YbviIXZf8SwSy9vXdk8PYwNygHe7Ra
2azgKSRGn78VcnwUgTKpKaQkPEaDOWOi3/RBFslaKbhk/D07qSDn5aCJnMCmEPYPQltBnvBjXN8a
MIri3Jnfw6Ywv+nJHt+TGC77nQM5RcyZDL79/y8jBM7ue0et7lwtknlhzEqBWWuoaql+yCjoj3b3
w7f14bP4cEKkbxa+1GMaDujd5UGv1lBh/ZBeBiNuO7S7/PkGyTjAauK7izK36Na22bI2HOGEQMPS
3vgD30vpIvTV9ZaSFRNLsVqOphuYkUk3k44hnq5HeryUJfoBpiMDOYtC2kiB9mdnWrMqdNyAIU3o
g6hi2fa2Vfm9xIBaepw2819RLRH5N20kZdrqVVyV7tne809CPMiKgDdpwnJYEzqFgzm7vcfpVDSo
DatXpLPsdb0Ql4hBJtsr7/3UzquXWCTmJXXaIFIOXnoHFwsUb+Iy4N9C66BkHoPmEOCd90OTwt18
5CHc6sCXhhT+snPTv9q7jjNp/SsC0eGiB8kfH8fbUkxIum8+UoIwxQuSKrs7ot4y6EFwUglNMFf5
3FIQUDuNf83rs+qy3CQ29KEP8jgcDgqz/a+HYBvdxMZntgELtO7Hw8yRT7F4sXrofIwMh2Ltq9YD
muMgjz9zCUP68f0ooVxoV2zMSnCA2/6Sy943kEhOSkUHFYGX1ODihB4MEvKQIpChgrdp8yaqRuTR
tgb1sPVZeYTx5wTILfR1nW7/USNYwHAd2Rs2ig+XNnhF/LIsRBJnEs7E7ujLqD38f7x1O1KWHYeq
Q3rzhpc629+P4vbaI19iX5Yp9f06Gih1mNYqoXx7EzJPpXz/VVHsWjcUoLvb3WoMmW9kDBUfpxGd
VJkBtBJ2/nlMddgudT+5CK6aME4U/qDv3hsSZiiPOVy/lSinF4uf/nieqBG5ayXFYVCbarzJJOSU
coFzh5QoOqi5XxZlzJMGKmKR0uY3GoaykwmjpDKxvpJTxvgMwFq1eYwnCIFsUhjE06y4LaAZnZCU
2JdoC1Dg75zOte1GFxlYUyB8zs9AwXE4ODeFOxerdC1reZJscVInx8pRQS8IAcHhDJXrU8Yxqs6W
Z5RVC7aDTwJqgddq2PkPCbXu5TtJvT92CJ0/LwHM2eLy0hGROpqeIJa2pDf20YI29rQ5/uuzUldq
WHTvRr0mPhaqkEWRYr86DXMnGuKEbBeCzCDKS0RZccBE4rko7A108zCBc3uy4E3BiqAXVGMASTu6
S6Mt+k3fYb38FiePFeA4vdgSvr0LDxC1JlDqerzrIwM5lRjcegbEzzJoC8kxzFgCcdK9yzAXmduW
gZFTc+CaVdYJdtH8s0KQu3hkibfuhpDaw8Clg42yeLNpwE5oebwmiFCxm+xUnf9bcA7wI1Q99ljY
s1n+m0Dj6yMBG98aQn/FERu9n9ocSjQFm+xCp5Bgz3YhfOM/nV/Fu7MM/O+wONjH1JzWLpOP/034
ZY1V+TvAwjAr0KNlcsE/hR3zctZkV2A887fKncLChV/nB5daU1/ApFe2WpgMNP0LPCpZB8h49bTL
HyyoqWlM9nx8tcOzVLF4UC91qfAzjVDW5L7g5Oz/AZaK3sOscaJyMQULlqVbgE5YNtRq+Jo3se8/
06LayR+su9pi49DuZ/BIXFjvUsfgmgk0e7JpIfFQEG9c8QHs6FgWU8enHa90fW/haQlwJIJtoso3
L0+AfxSLDw/4cJy646wMAN86RQj660uVU9X26bpspIq2byPGj0k+WDZq3Sfwc1LXDUCq95opRZAH
FYXwIL8lCQCpl7+SyNUH/7QWc+3906e05KVfGN0hfBvVEKsRyKJJ+ahp5RRq1b+OdYmatEQgCTGy
kD1spr3Gj8F/Ip61z7b/LVhRCZq79xs1lhHCk0e/OFtS3sMikUl3Dxno4L3IKI9ITChWa1PICloH
qo2AgzBWG6fwyhROEUlLMSjLNgvXfcqo/NsMvPQ/IlaB3N3lL87ug5FxB6vnhaNZcVfFQyHyMkq8
3Mb9z0Y6NQe2GUw83moiRj4jRJt8FrdPc3C1Mkyv+7PYy7PrK+M1BDCEBG4g83PFu2EMn9Z9eyEm
sRutoCYA4Me4h2T3Z2yrB1i1pWxARt2aaS4YZFMBATeM5E7QzCJ000YMxa5uhVzBd3wZV6nLLoK9
m7KAdrhvdINZjkoE8GbWSYFV6jW0t0J2PYuXfLLsROfqg+w956s/kBc4l0yzpnrHHE/eWl5jZuzG
1Bxp54xY8ZbXEZRFXn9UPKdDYlb94mbcgGSdctIP21cOcgzCW2AL5nzwiM85U3fPZikFB6A3TBLL
cO5Y5TXjE/qlUjfUF0t2SqzzqDVVzRK3DSwaMVEE+jYJDbnqjWK+WZMnVvMxos/6fiBmw1FZXGvs
+Cu0rLSzYTXZ0O10oAiwpKdTIOhu3zQ/J+O8+UDFfq2G6f8IlCB0RV3xGEI0QiG6Yhiyzfjuwj4c
m+p0e08fL1S/9VSyIlTYX+M50t52SI2RxEwNeesHDoYm6xAjkpyOzVvmfFtjmrFNMMRLHhAYW44S
HrMR+4deBLjj27xqn0LsnJLpW1qOz2bdoUu+ab1KMlKwG/QhF3iUnLlZ1upQLj2uJnUnrHgYWfI+
qotlPyrr0XmcceQbNiHmiVm4x89Lgi9zGNwD/hYBPChvq4YkvfWEY74ePX1mdlFbd0QkL50nFfvT
JO+RXXo9OR7+zSaUshGmoVl2gogO46UtE2l9VpKyf26Xc4AISA3avBFz1wmkwfosCjUE+pWqWmXg
3WQw6gT166mQka7Iaaq3cRTEIWDGGjXiWEbOpn7hUdwOMKhiEVAypUMh3+Lc3iiTqdFvJtlEHUNH
vja1a1DCAJ92PIyhPSG/a4GRYvwLvYUkdU8yNInizHmis/7TbRyZ2U+aPRLQV3LQOYnhQWSRAtFD
4bes9CZ1SGR7HMVDX2GwtyC4NH6CZ6GxhfnLgjkhkje0QMIBjbMqcVLOESUoFYnIET0bJGeq5JPv
D0g1g/zCXvSfJ07J6z086O188P26JPoFSja51WMm+dJ7ySAHfFI8N2fztuknW9qGWPmzDGj1ss0z
pUZ5foMIn+dz9pA1fqV6pi2ngs0HTX0ifJ9Rl5U7mrtiHmge8qVJC8huHk45ibMAeMQ5DWuaJFyK
emLbcgwldZgFWlbmq4yC9AVwphbnAlDh1YrIdIBTvQlVLMKwHTkS+pXumjfxKURl3+SSNl0Exvci
m5ZGTN6pl/w2B5fHThxMw0jEImFXf9OAW0WwwBqNE/ISW5HO5ToCCPKRi2wKtK9kwLTIEPACOeaf
mKiJcZziNTEl2f2aj+PfTdTBmQaUxEVTFegtOdg3NlAUMHx3ftPA1Ki7+i8G+9YLe7iQ5ejHLEu2
CR5lblwpqVcONxrzsDpkR2r1lyLHVAZHjc9DdjvvHgs9xxyybPskLFs2pnWNcBXRTXtYqZBw5qAn
woE3hRSjHwFI5HiGC4ThKEpHSMG3qU3ktA6XXY+mqFsvBDrv/0JiNgWy0fmwSxyXx5r9DrUlGFd6
QIRf+cZvN0CvIKFz57dlFHFcNL0UvTwT20X6dDaVv2cvPLqLq9uiXGHpEKcnE5zY4M+lJi3w1VF5
lxxGBao4I/VcEN0usVTSiQzMkDPfDCPcFww9Dm6d1wA7KdOfBZ+XTcKiJotV2fSxxPvUCgCcB8rb
/WGtRSHfB+xehGPv3ULmmaHdBa+QJR4XxOSOfHFYN/AWg39XLMXnjdDgMANicdN3En3MxDXEocEW
aefLgvT34zz63eUaXjG8iy3Dl9CjIVFW+yG3ibTPnvZpQKgNdmkBWD5vBRoVu5gA7kfcg93Qm7in
FTnwCTVeuRCSBcF0MJE1m8C5xWI+Kninwe24HRaaRMz+gBI2ll7brmSfbX9SFMOl8dv7B/t9Qd7m
xhUtjZDVMu6f2YdOWuDu21nUZQDt1tpOaMowoMsj8JCkcV18FuANfjn7dBtytRQPsCNqCdsIaBHQ
5+HBAD2xnPFKfHc1rQtNW4Y72NOOb9nYBzVg9qEkj4GIuhbkVv1jDTkDFbhpBsnuogBXdhnwFFS7
2YlopNlxOKU0fkzNEDBsTLmXqEgB1rDODQfGP9ldQNxKcUcU8rmF3F3gidCgVxQTA/h5B8c6qAEy
S708Wvd3M6vNt/8uGuiwb62fy7Yh4UD+KmzVvPsTOzlqWPzwTgweYNqgC72p1G9XI++IxANrapGT
r1C+Rxa4ZmWsoGXTc8+0fBpPBlGg5aLlSWB1bTwa5mcvG7br0a8LWtuF/DX0ISei2oEQDnhvybcN
30ud5SW73qDKRDfVOVoQP13p9d5LP/Etc8jXR7NG43/ZIKTrR5P+pYhH+wSQIpYwBuGfdR6K6gJT
ieNEJJTkvULRUdGv+EFAMcwlwgvV87+KJBziDPz/1Z4CdBDEyL0YvyU3wp/gutCb373zgi7EixFA
PlhwRDv44gLJD32Ec7JxizGalQy1okMTdTH5LZgwKQWp2TTAOMVhLFNgQCFR7d1FOVjkKlVXv9fL
iIbQuSHeSABZFXTeSRu0Xy/C7OAsLdDtsPkD7AcdxPC60DO6kPVtV1oOiE5KxK6UU595CjHrxBjo
t3krrqTkw7mXz0hvx0xcR59exY8xmZ3JO8jWelm4/7+UqOvsEkydZzZnUQtFWfpKnZZs+/sxQ2k5
8sCVJFZkqwG0H7JNz+OyK2Dg4BoGJlw2Lj4ry+mOMV+sJZLajV5xmJdrvOb+5y1Kgoe7iJ/dGikt
Q57SsZUXkwm6gX1U2ege0Zgr5pnDovXOYu0t8891CzxeO3tbfofQkEUUf6SCyx5VU7O0ITifV1Yn
UGQ2OJcR5d7t613yUGx57QBg16X8SbckYq2KAzdwjSsYw1t60g/TxwBWMtHwhMQmdQgKdN8QPQY1
D/32sYwZn1IgB4STkxz5yn1Z4oisu/T7y93dJWE5Be9zEzSzyMEvaMwSXvyyCi2eZXIbBi1LvLb0
G+BY1Mb/fHn1UF6gTHTihILFC7mA+uETskVGhoUzMNk4SGMpSjLAIuiGFwmCfWVhWZ1DlyW3XdEp
tRdwjCU67eTzr4kPOB2fSFGLEKKZVOxD3t1SGRpbigFUX1z74RlN8NKRwMTJQJ9fTFGTuXjgNibq
3E+Qdr1tkjfhrfsQ9YRL/AaSbYc6Ex2G9zH2uCELsEWn/ot0VhFnYmd7THL8AEkI2BmtZWnTJ0if
lEriTaB9LrIzHy3FfdzQ2KvOF/qX+jbyl3fgqtcNI+/mLOFP1TWFe86ajRoaRAR7SsrETFgzZNTI
zFacMnCH1XjELAoPlEXn4LifqRu3GaEagoiWEucKcZ8vVy9FkhcFOay8Gs6GJVR4WOREUrTS1ZnZ
KNB5FstHrw1XP3q6fd9AM2jvK30j00Eg8oOnd94R+0YzCH1w/3nF8P7A/phzViGrpcDamTS+zwb1
FuMwU9feEi8oLguiGq+vz5uvNpHDQI6pHV07yl7g6rnOltnOe96c60HgxAtLBU/6S2qZmR+orxN3
Z1Dx7fB0+WyMdekkNFRRV6mmROJYrzbQ0n7ZF0rS+DlGZeypX3MokuJ6yXIDc4sycDPmwV6/KyV2
g7A2xaagaFfyObFM+XHiFBZETPHgQdNqw3wUhXfEMR9htt2NiyDDM4kTtaBmfGmzPNde9HG+BQYO
NCHJsqmiE4BujI0CoW0vUMqsqurb+C6pHPVuELvazQQ0Jl0ISi1djGcwsZ8I1U0RZrwQTwfgaXwR
7g3QrldwfZtjA6uxMCxVkLgH50B9xhhlAOMWjwvHXSzyyRd1kOVsihF3VVX0KzT8YOWL7oagVnF7
SsJvdqc1Q5MQNrUm9iBVW7PsVTwckg9FiBiX2WKabF3bZ0EZ2nhUEUE4Sz+IR7rnLsHDAHPXeIwg
rPW3TqM8XnycUUZZLp5hLGQBLvNyGq8GyT2AIEYmEfp7JXsjRywyxwyznVgxumhBwg5oCrprg5NR
vaJpNOZInqZc3H2dmPL6qmHUo6UPMQ/fHDi+2Hbd5lyUPZ5G5Q0GFaAkRBGmPObGXesf0WQ8IjEp
LyfbZcjID7SU0mvEJpNZfh1pu7VdmIcHHq0WnEldvVroPZGt3bLB5rd1as7V2bCOLzVFIBUvMFC8
DB4AYq+l3w8hWMUIma22M8qRnALxrR/gp64QxcLnOUZXVCaysoNS0Y/gmMMalXWq/Pz0RgAww07D
/90jMayKcBY0Cc/E0rRCyPCyf6oqRSCBuAt5FjZiV6YA8h8F0y30Uvrzc+D+seuiiR8kj2mPziGH
R7Y7rQQPLJ5pM91wC0POpeb0mFi2ww6ULhIcwpep9XiB2L7zJFHHg4smDJMhiWTsobHcDB7ccn+S
72Qi7pIbF+J0V/mvwHf7bwSQ6Sb/EfVhlUjB5jbv1ffYdDv6LbK9dEO5rSA8g3X8/Q1ChPkJMxd4
2Y7pNut5U6FGqvxOEpGEGqaco5RBtHSQ1i9HFJzZbSI3SLVXc8esAtphZZwxGoNCWrDX76V6l2Js
J+OtKnnQxDhSFOROfPFRtAZT5YQOdsc0AZUuEwhjNHilUG35IGmVo1kSSVSv/zCklmtt7lYCcunZ
lIY6hsrDY7REJfLzZUGmxY1yLf89lwNX1Arj1YyYdpfP7vVWedeKnnLkrXED0oO9kHlgJoRMRJkn
pEQjDoW60tdBaG7zj2Z+vIPtzqmEybnCyB0QSvLJEvQRFgNqSWLgjTZaShuqfIWH8Nc0/YfMzHvp
OGj0q88SgxR0iHJrIaoDgquTJeiVQqXCWU8g6PpTXMJxjJIkmVa9DPKTBjsxlX8T7eJxpiRQ4HFR
WqsqoG/w3YNPLtIFgl1lKnH5n6VHFqdDDjH2tyGBLDZ5wMXj5S9eplheEgbrLvmbcgiYBFNQP0Yz
EA8t/OkWpXrDRyP04QQN7S1XYa8DGlu9KGDcuKok/KJS4P6TyhQkCy2QkzJ2puACuOzEd1LjDGNF
jdR0GbVsTEsBLvknQyzeuddkQUloZnlCBXxmaP1/nOzCai3TGIaqVxYTJWAzZW63CosibJHlvmv8
vnUrekSqT7H1+jdtvJQpzBotCu5n0LA+OXiA9I4VqZpcJzpKxmC3pqD7HA48PEKtvG+g491mp9Zc
oXT0LId6OYipBW/vPZSfGzOHev604arNr9+vKoaEufbcCDFcH+fPuC5Mi9DphneToCr4u1AH3kAG
WGvzQAo9rHB/Z2xY9wIsXlXdVspH4C7rMC5fJRuEbJ1334DW/sIg9Ko2mYBzAYWe8t7QugqqvzHc
UiwgdTFQXWw1LCuJ2jXBw/kdB3Y4sx2xA0UZeE6O9oOoBEKWnPKDgAYdLX8PeYMzBEW5mbVh9tww
g8ghNzhehvsrNsHzwdPCB8eN0eTu1NksRRCo0qQK831mMKY3hFHSjx1PtSgHR3f9JrY2WKHh376R
YJa+mDnWK0tY4qK/Rx617OI66MaY/Ml970IylvQK3sOFnU+HyiXusKcPw5CCUjVWrAWk1BKW4q2K
qK8yvGoyTINi1SpkV2i2GEfxyaQ7CF7r1SEXzsVEG9NqbBa47/Kn/S/j5qUtx7jXG4VxYMH24D5V
gVj1kUaXR3OAlrdbTRxNPWIY+tFDGHzHWh07tQ+k3zbIUwFG5eeq0HI+WLkSZd/znurb9PCFTw6C
UJ/idWe1JaSqWZ4Wh/PhkWBtAPlmPxVz6cpbdozgTnzzSAujKkAvJrQ2ygKUkIdwDDPgbO2pUHAz
peAa7ls6yu3mASRmElRBYmQ7WxCvRI5wyeznQwP83NczMSEHxDE5+uhuABXNSN/glU914oL/oTyA
TE2e/PRl6qydDAnDOl5w2qi+aKQBPjCc7CpRHAXnbLKXmmVDZXEfZh7W7BFUCxA2QJfnPIUplw9W
ESd1dX0KyUBKbO4rH9vaKabRXAZDZBsq7X9Uj303mfYQSp2o3guQrRc8xdzgSqNj5z8TWd2mDW30
O6qW8Uh8QTqMGOwykS8KrMqPBtgash0Fx5Sx4JY+keI9/VoYCFw6cFh7QeI94jt509TCPNvVfFMv
gi8QV45tR3vbTEYBKOrLyuk2Y18TAjwaGn2+N8g9ib9uiV09LsPAR5CyyVYW4lSGwP+UOSVeFu6i
5r7s9OTy+B4AeUglAfBKUX48U7Sb6tY4p8Qbrdn+GVkfOHa2OMQy67PnYVUicnXIjmUutorNbb1z
TZuqA3gYYr3jbmUnagPTSoRUKRifLz7yPZFoa5ullQ+gVL/FOmNN2gOWIkiVXnd5IcIR80uzUMtX
6zgHqBcjonIT9yQ/kVwQpQs9tdXbpBaDP75UdVitMgTmQgU56Yap+Fw5qNX4s0aHhieH3CKV9N8+
ZmgmnhiTQ0fd0PQgsjJLlKRtiU/uwzcgiZRsrTEvs1BEtfux3bYZ2NxTwVkyv/ww4P0IeJIJJ2r6
aT/HCp3MSFhqv2bpY0Hix3sLdJAPCvNdlMb84eeyn7npLC6ij7eR25CZE/7vBJBzJHnYy21pa51x
t0gPgl+ejmYKLS71PewiJ5r5m8RrW8lGfdBs90vn095ofU/ug4cz2J/G640V5dLi+Kipjb/0rv6y
4xxshpHhOKXIUu0t784KNUTZY1/43KEyucpcNu2zGzUneTQSb0wFJF/6FadvmayZO+9tPgC0xJay
KGj9nBy+qtWTI+3whXQV2jMsSx0LHjmP+eqJrRDoT9SeEsebgA2KVhHcsHqu54J4T113biPeml6B
qLPa67yasB4r0yYtL+1045jOWjbJIDywL4clj7OwWLF+q/BObWHcTYB+ViJNwiMQ2lL9wFFe6p43
fnZkqMS/uRFfV2F81Nc02sWawI/wv37j0BKjpMYhXs1KtgWjtBudqzbpW1I+BNfTCB0BME7M8luC
4Frd3TA8ltHGO1LxAIjEyRt9y67lDN9H1CWogkAQTqaWCpNYvALn/UajjQ9JuhHsujDPqFpl+Al7
3Xw7qnLBTA4iWUxPOMHmHt/j+Bo8Fupltg5LIiho/Xaz3cJKSuQsStuis8uWy1561lFh4gZFBWpT
AO40/F9StG8Ci7W64mD51A/4+hzm2e4EIcD8+e6Oc09RfDXEzoReM5CmLBK5szEDNijcvcsAdXE7
D3bQgEWOs8HwY7XsLD2jV2p//YgtbF24G42z2UpVXOfHX/6mLEbGArD99nrouxV0QquterDBp+Da
/vkz5KGXyd6zgMSNApZnTUD7AWKkhwPIJKJ/YrOw8HIpBUnUdbK+jMf5TAQe1yrsouNvy6/JYo5T
jeXI8tUGLU0vsrFU+YH2xfoXMsHrRu5pNuBNw9XQdBIeA6OIkYJnbtFbZSIkOUM+5cfNnSuEyghs
1Y8k7/Wg9lHknso8YJM/O7rnckkcRWAWKBwQVCVdKUYiv/4iqFK5yyuR5rYlvL+30+j2a7fSEehw
mlyekd1UGQ72NCFx+mcUu9cQK69pyAF1+Hsh5u1Ye4RtvQyQOQoeuWfhlzBCmgoV8eqpPaRaVvru
5n1mUfUiHNB2Yc7rtBRECQ7l9xLGOBgY+e/ac4tNIezJdTqjdZhppAg3ExSh3ZhbCma1PEjfg5L/
Dew7fgQEjPHuq8PoQYuUrL4wfNTt3zxdaf71IPsNtXet5rFiEIM8ydzlpRGxfKOmKKUC8yM+Ny5I
kTXX4qorGl0JeuaN9Wid3Zi4sBCV3nLz4cuu8OcRHaXYpFUQSroQyZreV4GziWZpoGHju5qZ1969
fUQoVWNSfWttHP8TmkLZrqlGh3CKwmdMuJFjfUrjMtVvzuIu1E982EIJVwws1FKC/sWX8ZT34Olo
ub8GcHdjQkcbo1NlgYTfzJ1GkB3mWGFG06AAJuaEPPCJ+mr/7BQhZFkL50TV0F9p6V6G2f/ekvM2
eE0+pVl35+C3oEq6V5It/qjRcM9I/MowsSfvMkJygw8LlHpwNy7uXHWkqfL9exmnv8JXK/9bvlF6
M1G1Ta7T3m7mYJylDNX3zCHpmAbAJBzDNxY5hrMaPBbhN9vyi2YsgcCUgykJ5QQk43b+Kouu3/Kz
+uFjycTcq1ktuzns+7mqDfkv12qeDsbPvQ2BA6WNwlc/PPKaWeGaPCBP3IJxPHCO/cBJJBc0YAFY
dL5Z5YhdOFfu6yFFBgdP4857ntgZCOVS8yHnX9WBjg+y4aPh+Nf9WfGtzjnJxnREkxlwnKN5tr1f
odwFLpSYepVO0z0f6rQSogL6kZTjcs6lQMNciRCCCdmpBoHbDmf2JTmZ6KWvVnJlfrQAfSjz9m13
pKwvLW8c2N2sWxiNCH19V/CjDh+RzadGVkn/vStfcjQPyKBOT67KtzGN3H2H2QQO34uouTpvWmV9
CqAt54RtO9nyFjh9xGKX2vRnVtOMeXzfM2LJ+3uSTrh7ySRw2orb6rkl5aq6dSWsfpIEE+QtkMtU
hnXdlqgb8WewQ8+cQMWInK66TC6GjK/X429mSY7/qy7cE9xMVPJCm79Xdxw5lc9MYtL05I1EVobx
2IJJgGEMNoV7IujrgR3tuboREymeN/bxl475Y4P+Yxj4X190Tz2KZUP7spIp9SXqUGxUdi7OdDbI
/wHiuCGnrlW31tDluG1mISDAkOeLrx8V2G42dsF8ijgRqXawcsuXeqG+T0b7e36rCtXiwidiejtg
pKxXnChERMzIQ2kGQUG3p3SY43sQAQ9ebl2sKJXuLYV/PhNslAgknqVoNOkbGar6DeTNMDOJVkVO
k0sa62UUOtV3mDLIPIMdaZKW51hZIvDjIKCQvyW4pMMmWxJCDG2/BFMS/kZXv+NHSNrtRL7tIbTo
sH5IwlxocmkzLc1KnWLBL5DenDWA5IH4n6xtNhZZ5ykYsIWclmbMK7nrnFKV2ncfNU30NisMkFPF
dWxgSxes5QmXo01XriFsdRJCb0sD/w9nK+FRrlAeNn3f0tiZCrhhSmRYvHxh+IFdUPcSAVTM9Y13
6DWliWYGzzPyUtjb0KE0drAvLhtQGw7piyiZnkLGihb7JKw1Gxi3jygHABPouW9JapLrr6y3JBbt
Fus9WbEdDp8wrM0RrrZ7qzYDkIVkHdwpLAXSesaGXXqcMBcVUWdIAmPkHU4Z/cUQGgavqKB7ih67
M+hVKPAhXKJ+97tQqklCbpxHd3COdDkZ6WOTL7H2ySTkDDEyAF6rm0d1JAYEzRW9VmAHlG/iqw+P
rHtA67FWctu+d9VPzYUluCWQhOrAievZP1n+VPeDCBNIUg26qhmsu27sbLwnFx4LdxLcd1sW4Gzp
RZLansxFuEsYdhhr1TpCgQJbrDf8spwEgxrftacdyHXHNNspIWKoGX1C39VBXDG6DrkcC+ZXGytZ
pWfsxz2ulZJNLauI9+hVc4+uO1pBKYhQCyHV9J5khy1hQkkLwgDEiSS4ODWHXu5Ue+nIl57o0TEi
iYop+Lc/6+fxlkR0ip0pBzYKJoWlWtqQsNAduauMqsZ9rcj3tZiTlNyc7zg8nOQ16QdOalvtfo56
PKA7+3jxSWKRBf5lzQJO8FBa1e8I8RnBzzUtuVPEnjBK7YB6txJq9dpuguGNkZurEU3BAhs0J/kH
/wZS7OgyFI+/Vx2OjS3ABfKIIIIxs7uE9nTVGmowBOF9Kx/8K0v/qTqVK56iWwbAIZRFZ9RHliyE
msc8I491h6vZCj4oZIU4DcBFpsGlkfJbjHbupifsdceh1FxsVG+dnfD2sPc2gcN/LBOjFK1s3SHD
j+2cyiTVmjFkLDAWDaCtkpVHdFRD2x5jrcQ3CwAgA6LYAGRrK1y5UdfbUFJKuhnE25OYxIiEQaZl
eAjVzMnqhrBLfY2Vf12dYZ0SjrP7okZiDHVxZ9P5Shzt7nA8lXEY275GJD4MiZ2vbo2zhpLpbZ02
OoOGkYGmNfw8g/9HSqDOiTMAirlzB+iWL4X1ot3bS4iRMt9vFqPkWGUc4IN8BHEIM8pt299HK64o
TECYMX+d36Hfz7tlVh/FkhEFXuYHuxckz6+GzqjtV0pdCA2uzgxhz6kjZSyVmQC/ajJjMEAwYizD
9M/nCa6gnCzGLdE9rd52RUv8QYjXuaaef622hxtaqpIcz2L9Fm+E+9v2IlgFamXyYxkTT2sZIBKE
B+MjZP4QJhWZqpj/er5KRk3NAzKEh0zjuUVGXpA3rW+TSFSs4gVHrkUZO8YiNhEqhVkeWuJJwsxb
sNZ+kCBnabXx+QyjpL/C9YLuLdvIglu9J9s9r/hkHmuJ3khsMU9cEKPBN7vPq18Ntf/bl5T8XRRk
0igqVuszgE4OL7in6MaoKdjpxH1Ym9pvFM6fdj77qMhYGu1KcVb6cb5NVgFKhJ2mgn6cU6hYebKz
B3W3gw9/Ezi3zY1iSrfaSjzKbbrp04hcJ8y4DnQzqSlb6I4w/tQ60pmkFRnWadt8/64WZidw0eGJ
ohv6p91IYf0oMYHc7A8GG2Y2zyELQ9i0d5yyrYqHl+5zxR2qWxntdMr1NHFdQIaLx3+2IuFyp6KM
TljWu6Z2icBBkMb43P7SHqYynBjubNZlOeBF5KLAmTW+tuuv/NGqGmFNVJimf9cJ0tke6sx1xVB+
EOfGn7roPeI9qzdfqoKSAluAjEKr9Df1Q024NadXrXU8+KwhlMFrs0qg0h+oMWAj3vuxurqWkC27
lc98kX6sjUXf0sy+W3At21oEIF4ZlzD5pYLSGUJPbw2+2YKzB5qQu1TKiE+tQYfzNDqFHHTyXz7V
/7S9jqKjAtgZtFKulk8CeKL9VtUyCDnx0LtdWfNfHUgx1nZqxqEH4KR1nDDt3MEZm8mKgEndbg/6
35hDNSF1HAwTc4P6taw0wcLtirO+XfRN8OB9fPvmcmybL7owWlUlSKnsLAvBVa9CScCUNyL0CEI/
YGF93Wed1QmXJjBkvmhYJ7Q4JOuKV7rb1/ikPXrTBOhUCFl0l3mavbF0KxSRjvZRLWo5loDOKsAk
dtekSSC2713sj4/Johz8eqpX0IFJi+dmx3bs7uktWyyAmi8EGJeE7pvsPAb2lF+hmeo60X/9DMma
pudxIxAs9xXp3cZ3c9AUNmv9N49uYWBLoQkS3bEXXR8KyqPq3lZLW+Zuf5LvwIqH5XhssOaBXqmb
aNPEdIvmJX5WOS+jgUA3+gYejLg5l8wXHM8JWUKhvAjvxbTo/GacD8odS/o4PKvGJX35GwAZnfJT
4HPDrai+itH6gh9m0vfSeyKxfXzy3S1p5dyHAHbGXPitvBobg02RFbuBsTN9cRGbQkV2d8i9cDBC
RC7tSmbPUeWCki0zjY0km1v2koP6wcTJYB/ydt41HZQvfWVwL67W4IeR60+nx2OvILP6ddkFufi5
y+PFIN2cfQ2yVvyFgoHjlWftGH0c+hQ3kw7SYkS8zdXIhPtHQCXE6GCHYgAnW/XbPbmhmp2Mj22t
LpCeSTlwNCfdnOV2kAIVXGgsV+xnEg8Mb2TrEXV7c8Xp3I+LT5N0wLG1g+sW2rTHyP+jNz88bcXC
l42HGAYI5L3iSLxe17XaGBlwUI4etndQG54MmiZoiPU3d/1AImACLDuKfZIkeWPwi6gZhMpxBViI
uQzJ6b4OZ3jokk8k6BmFHJtu20Q7HgkTfJKuff2WdiI1JInTlsWUdu/3ELkmSatsSOY3qpSfS/QI
QVDFbsvQz6fPbO30YMDIQrSuxcZSE4v3TCDx4w0Z6WL9W8wj2i9QtOls9xuChoexrn7yGhlTsjzJ
DXKlTkO7XXlKY7HoSJahdGIEBOGWQr3H5YDQkdfpoRLMz3Jeq7WYuZmOpL5ATPZVTKKbDLR4+Onu
dIwkOHckiJK9AYgWuWSAzeF9lhAu995jRF47bBr9iuEPnSsTz16xWDtp0Y3VEOTSfCH+6qI8P3Bq
Gq5TjaP5eDltGPz5j8WVH04r9r4ZiG8KtDEDUfrJfs4DWusX7hkm/G1hxb847/ZOqdevL3tKYVRF
62MbM+ZF3+xPj1qMeEQDtCiGZg3wJ0/B475fN/pZ/rv26Ab3fr8Vr1NdeeJMGFY3NyJtOCAfV7VA
EJvwoF0jFQZliFu4AeNoPk5mTFxmT7IU6TwHC0NsaEu4EhalXEtcWm/BDAU9srYXVbirfpHt6KSD
oEgZ+UHseQG2K+QwtMrQ0iOlppL0ZlsVEIB4IrR2Um+EP4PO7Bn3t0mEyUDDYG30Q+olZVVpf5Wv
CmprVLq11QiBT3N5HeejZkAyohac3LjbxbF3tlByLoMbLYIclQ7P7yWCLqA9378HsYZ0Kw7hbYnV
D4/HsFjYlsXpklo15N9P6Z/RN5cF/S3Z4h/M2JKHrJWVFjrEmRdSIPRJ8V1NNd14t5KASDewC+Rk
cd0U9ViXalWuWRM5p/AfHj3dfMBBXHIfkQo8A1Chwg0T0uzzjpuiex2+FN96E2tRHzcVyzyVVa7j
BIT+Wmo7Gy4qsSQ2j2DzCm3LhH/zeQq94akE/1WUKw1f2FpSAhlzb2gZXH6jtOZT1/k5443o4N5i
nTIbihwYkebX05CvEAeyXGWlzbHqtPzUqeC+zN22v6pQ/PlIsPS0q7HSS4rDP1vNbjtt617Kf22T
dpq1Oh3pYnLaGWKZmj5d4H6ndMStG2JzQQfhjw2c4c14XlFxr0ckZJTm2jZsJzo4GHqxOthJGFn+
zn5Yt9c966ma81NyPPS5zaEYadZACY5k7AobBhY6KNe6Kg2nuV5X7qvm1PeHv+XpEhxorp4V9XKo
qxnw/H+6LM/y91Gjihca44lmaMPZgPl4xsgCKg6KaCRaAbMzSYgnnyzyIQ/outKNWBIFMwXVys6Q
ebRQYV/lZaycGtyF5l6/B4q/zlbTp7o14jfCURFnPTOGZhRXPjM5qeO+/AevWY95F2Max+CtCP9r
e9rGVrjdMMZgYzL8rATML0DwRniD8+QvdICxgEObBl/dxjaS9HqH61H3k7YGw9eSU2PyvrhtxbM0
SJ/WfTqcJk3Nb6rqy0rFqy1Pjip24/e3qIhSTlSSh6pUmCfH6GKLa1q50V5A0CzBnNR2NsvLS/wU
37ewoaJS40PIbME5BIlfmnA4/A/SCNTroh/+Ou04tOlFJd4QJhs2yG55gZIAPYj/fDVrQLXxjINC
8a24YluA3EfW5w5KBcXM6zg55wt3hqa3NjavJxwhVRMF7FplrEdIjB5h26I82BWwUwETdi+hQSSx
FQn0je47nwkV98KFrCi7ZNYhGnRRiOWEqTAuO4Lz1b/i98LNLW8Iy7dy3ESG7LutY+SOFPiLTW7h
JjLX3Q0MOhC6oNESHhwdAOOWXtXfgsWJ68UQKw5al9rGL0M+WGCYqyLnWmRbMSsNLOuId4bvvRao
s4L65B4am7gjhpzk6o2Oa/e3hEsq7LpGl8CkEOOjVkqTHsWDC5BYinxncrndJ6aRcuHP/bOeh/9G
fYKbl6UPfp0wKGKfaQvCikZGLDlneMWdcZiY4nC3J70VE7le6NL4uq8mgm55kaP/NfjyJX/TZRea
qRbTz0gbqXq7M40mtsReBVU+dmOrzhZlD2iv+Mo1Oclff6k3nYaDI0Tn1rmFbJ2RvYyBoPSkANn6
PzH9j0CZOWDWj8ZS87FV4iUAElKS3LzRMSel21xKjnc/x5VY4c/nnoF9rOdDkT/uBNeiQLjVXChY
fsoHYMRapUWGeVX0SCnUI7UJTLCfnRbSw76tv31wlyoYyFxQvp/VreEBlZDoo3d1rZxzZaBHtUyW
O+BEBsA2D11R/T5PecvNtcNEuBdcvJtDYfPeBegmDxIfro8+itvSzO7XVI0NZSmZLd0tGQaeBv2i
lHWV0bhhYrSgOY8Wp1jGXUmMaYgCsivsL/XKJqHMyfqfC5SI8G8XSfEotfIHbVGfhJvMct6MKj13
jnI3w0IBx/NYNznZf7tUioLc2Vbn52+c8WOmlq/Gq6dBmZvKxZsoQN/AWIYKC5n7m68B4AkOArGw
arCzSmw9yzpGe35QIPg/BehGj/CVQKeneY7oeFkuGcimSlESKYlj0SB/UZs8Fvl/y9LyIlWEa3fj
KooJIl9PJRaCfgnMdGqYpHBhwhusq1MpQkv9pghHBe+jnz7PA8U3EbTJMB5OEh/I6FX9wscLarXu
4pXuQ5O1QnTITIp353H1gN122/R4iKF+SNkVQta0eAMpGROlqBITPAG31CU1+9+cuLFBWxhmnyDQ
R0JPdlMiqzywK1gUtvFF+c57cWocCaF/OzzFlrlSo3hSNvT+UCyyFlXA5fwUwccafd+4ElifuI3r
ErESRSWsP4loM/2ZawkFO+Sf7X8JzV5aAAAYWQMoW1XtBf5aWKNAlN0ukCloLMB3o6fHE169J7U2
f8TsEX0A8xIiCwM4YOTstTXLbW5fU7Bn8cZmYVME7kQ+G2a30qW8a8wWDYjSLjfMxq5o8hcyFz+q
hw5xNMJ8I66CEqQEzs9O0fMky76OhWFGTSzgT74+ozjkMjqFk3W5CwudharicljVqIhIi6ne9dX9
6EdfUU9P2MHbu5Qxm+iYsYnGmkd/Bb4N8JP0Slm+i0+pL1VIGr3J1OBFzP6v69tllbUj+SdNztQI
1j1WoJ0NDFKP3cAY9itrRMK0rptUZyYq24fuH4V4I2LS6tEaazoMqxjEFYiHuZqlObG/2z1RyAyP
P89h9CxTd3cJFALABp6KXQl6di8izpFKOX0ICGkKVzsO5/tBMqD4SNGUiXXpx6XKEDDeE5H6mjP2
rszwDizMUTf2XzMIFcx4kO8DtgCgssVDJOSwkGay0qXdd1HgDgyzaLOOfD5lCxvC3pbXtqlazkR+
LPW87FJSfGtrwpOY+QNwZx8YSBgGyIqkCBCwHLVFcPqwzEoI2euqCd/gQphWieTu1fwdQWs+Bu9X
tbZrtRNqCZcRMEEkosXWO6kB/+CR6w5emPbk5gn5Mn7pSO5JhTflhqZILPaiOMOyw+a8f3Gltx9G
fs9pK7ArM2bLXzxtOkCBsRCbkbgdsS4mXNxF3sosdTH+u8cZ5Enc8aT1gsofhjSWkYeViUwzY2Ra
45Yfhfy1vemhkVCGN3/kSRlGv/C4kdWamvGZU1hb9UMNi24XgrplGfpNxaJ7FSKCAGJmYiXPEwhk
ntz8TAxzJ6aAYg5wCQaR17M9KOOldprXl4WiO0Yy+yJxKJVJ/r6SfIpzEUlR+NueKabxjLsyV+/7
On2Tv9sz40fTNJ+6Jc6el8fmgJWv7jVoxno0LNqeAJPpFmd3rbT2IN22pyf7wrh1GqneAyKgMgu9
CrZjDPS44/EWNhCegW/S+BAN8QHRFUUNFjPQ8L3bkZJR5Z198KymiGPfrpqRqUPHyd0fKRFsOlEi
20Z1yINPwrXymjhkpwxDY+vJgPfEFvFYLlYw8Kg7Pj+fPuUKdHGuz9pmihPLeLbM8azuZL1dPFGE
ckXFctDFK3cP1pf0JviQhtLPWasHGzVVCBLZU0mrqz2dAZ8bR0rBli37kiaiXCdMFOseI9BGyg5B
aT7icUlf6GyUVeUcJ6KL6shPQZMmX9zJK6tYyHNUnhcsyMKZAAwc1a22Q9DjONAFz8AKEwBjBKLK
qafGf1QT+QSuQRjbK7GZ5yEYVRWp2rCOW4cz1LIV7cZidZViN7rn9mGNcgULVeMHhVAwVfV3GSag
yf/O5yI2Bqr53VVT/J7RvPIdgDgTUteB9cnMMwZQPiJ2juSCWlXlT2N9ETkzO8Tg5v9bPAIQvJfU
Bzkg/fbngI6Jpl3igALuanVPyIHHeeH/KXeL/rypb0FEK5DsoUMqj4HM/GZWWrSCitsPksqwJ4xk
yt10iTi8aJ/TK7pu7CjvMME/QJCpLdxo9dTpObfyq8W3zA3Y9yxmhX05iLJxFvh/NtgDEDV4qsRR
RC2TWK78cg5s81jdYvaaos+dXdDLGspwjYtWG/zuWP9FVyug79zC0IV3PRKrHARSoFBV7cEiya3w
girMH0K3TQKtnrnhcK0qwPAI8hxkxaaRhAqr7ZLGGm4dxlBoOa/4lpDOG/yoSv9Y9YhlTU/LNIuK
OgObrUD3aS6eClaVhVxrPpehSqotEM1ZwovCEbgl199xTO/dle8CDqOSeIWkIQW/6BtDnMP2Rqjn
oBQy/Ap2hhb3dcPCzpSLbubp5/6pcWJMo1ASBsYMX/gJn7ZBRyBOhwbCWYGnhtjbj4396NeJewST
SAC3ocMV2bD4ZgSj3H4AWe337wNc6TNoD1Pd1DlPdCk1WheS2qPQQCQTbBI0vMOrpMHcQb2mSWMR
Fd6ZMNRmfrORalpiQL86hTWLLBFvbpzauENLqqj9Sa0C8M/AjCmsLqmdBx4Ilft/2k7Miy2/u1uj
MOU69jCNCSJnuiksOMZRKYxiymi7se5/1JUnBUhbPO0neYsaafHzZVNGF1S1qavdB+wra1YjiL7h
pkzOEOb8FAi++kVo3NyBaYO8YXU0N25OI/Fg2LpfA87l8g5+jNzjUAcFK12CofaXZRqf7u5sT3gY
NgselCltP5dgasgC4CdP1F3/ioydg2o2Hc5OK0THm+uOoWpPOkWwNk+MHRLvS9alDJbnvQcuMYVL
nY1atiZRePGvI/x5bH6zT9gCHOwg8MYlFm5IaTzfhwBst3Fz6c3qYkII4ZFIOFo8iLVoihcn/egq
kPUKRAkN6ntvS41lnaxDxRkktnlcifIN/V5wKeqqUuMz3o55Lh6XITlciFVjBjUiywH8eM/ejAhV
EafiSNtA9XlzmHeHHdPerLNdTT3ogEwlPP/kxr4E9jMIG9lVmetgJHADgGOTIF/vx1DBXBiG64Ki
PAOQcDO7jTdLQPNyQpxGvbxtfHGZgYdo0G1hpMN9ncgpgRp4zI7BWodu+LbWc2Ji9KZXHt2KY8xa
p7QHCNo/5QyuffNvaZ7VkCUmL6lz9nqvDQvlegKsenNzj/oZHx77eArsKb+t00cEHADGQ6CHmDtB
IR49RajdKNYxcl84vF/00XIDbd3Dna0a934F8Gnh3DX29efeDVpo+blRucjL5hJTF9h0PTvPwXFH
PE0Vh9QrgzQkydTMXXnfDDHENnoZN3hKcKIdO5rgfIygxFPlcSwJCOB1K4SVSMYkUhJa5C2UQxKW
oIxr9RYJYtUYDyQ5Sew1kFgDqaFwD2Rb4PubEUAKGN4mSpWsPTGjnht1dH7+IUOEheKh2686fktV
7nhLTheYT5AQuiOzVOOoKZs1dlcCcejV97wG8j7DPzOcjRNvMBB0MsfI06yTn+6QRq/3D4/ktc8E
NUnXUeFxR0Wf+FcuOqNksvfYK5iqK3dckxrCrDcHtHO6GEffIbmfz3ikUVq7WoWybNH32+LeVpKu
fKKqhBotpiNaCTrDBmi3UzUlQJJ1QO6GYIqWOqCBHAkh2Sr9a4Vqw9B3z1c7y3fxHdRdXi9BQx1M
8EFaQSF1jncAb6lamtaPTQV0x9BBU2zqA5dqq+NCbymrgcYNIum8Z8ybaQdGQqPwAXU+V6pW0zyB
mjxUnMpn7G74fdz6PFjedE0D6qr47zghKQ9D9S1Hqmrf02qlimcmrvUKp7/AUmGheTMcgcDUZrOz
UBFyXmbaJoCeclWpx1kuhs2Ld/UYamANpN+Nz3qUF2lXN/8MhHjqBUXOmMhnMzbM1V5Dzl8S3QEP
6zMfZL90eaqcgV3SIwV/el+fXQUi4GiFM2ZIYw3tojH/obgQYLkw3wx+DnIVLJRDYBYkaUq8hxsx
R83b2KZEenugZbmx8l6nyK/rg5Kx28kPQ4f3ZBe5gwU6AYHY0AH5/rGYIlT2nDyYgSK3+ccdScHs
mPVNXdfrJlFdMW8A3uerH5ilJlmzigg1eE+QCIVPFcjMww20FxkjG6aZbFaEwJkbZcm0kjo/TKe8
/G21+tE8DmfoemVAAp/uUDMp/RAumNcSLYdc+N9i7aRDx3cEI4wgoK+6tCFQsTZSQvOojEM4v5HS
wwohX+NOCPqK0ItHyT4uPivigN7MFbfyEkJIOOP/IHocXHH3mULB4kETq/U9W6HzbwfGvegXP/aZ
JkRcrWy4Jz759mKAR84GhhTI85TSDD2rrd0aKojqQQsZGxSfZtgKz5fuMIw3z+NwaaTTD4NnS8tJ
K2AttJHooGucJPkIHKoyH3rOyhMt0OycifxyPIy/STchXEhK8EhTvGrf5gyuDb4Km+A3g6Y81stb
knU8cUKJGIPbAmwfPcGfiNSCkt/LDeROkCLEU+WaQVFS1hCw4IVXRUytEx+9ZdicfoHVqIV4KBR0
Oa+a2s+uBFHD+8fSwrOb5v5OQyEsq/i2U8Z+QwMfqG0ZQ7FSySljQHtwBVKKHsRa9e0Ob0hOSQq7
wGygDt68O7y2KdluSDHLV815T7yU3JpEoM98tsAFSF+nlDEsPZzxcWVVtMHHmNjO9HbcgQOJEKk9
ydBq5C1vg9KbR+Wug4tb0Sl3pLlaufkiIoyWJkFTGkKGglejzavzWrSGtjCMohRiRN0UViWqJASQ
G5qGoK3IdiV6U6LDSm63NjnpY0qTrnt275vSYkkdulBKYFWolcF1Mxq/eXeXv28e+G2xJrvPwnEY
JGVO9RRCqF6dDFb7290JH2GybC12NvjbZmQsmo295zVSd6W1uxN3oK4CxtHYGvltnMQ4fWfyb1lt
+UVMsVm+OI/ZGUkzqpqe+eZSNMEUMWdJUbbZ0nR2MhRWOy4MXY8VY8f8ffO5WDLPze/w0z5luAEw
2BIc97Qk6eYsjcMD+nz9i+d8oz9CbeDjprvZG7j/316ewResp2nr2vMW6fFZauZIYtdh0wYKJM49
wUC6xoesHes/SF5Cnosr27DkFCeKr0d6JkObdFjf+7aQuUXie/xR5My9CQhFZBqbzkXQmTeu6nK5
hseWe9sXG0afXGIC8WN0fxYiBdrodFFdpk0s6112hgEBYWfCn3QqYExN6FyQ7rmZta3CpiH7M6Q8
X1jZt6LBQTsF9V8pQOS29gcDRyfOBuCGvmM9dy/lWgWeTZR9nanwJFRRGInDVldtcYFhzQCJEp+i
Xl2zxUy48fDqj+OUZwQ+UhDbtfSkXpc323s+3bSl00rQlxDgL8pJ4ksS8JsoumHbLltn29r6nZzb
6rSlojVmMScqdgzVul1UWebUkFEzcAhtvdHQnb8TECzZlXjKPrsvd3vN4TEfm0OO2yro4DfUI5qz
Qs+1RCFuhmbHyDCKaMKYTTCk+72OiGoNvd45Y8gE0xPYx0rVSrIweVgmaBPkYcVQ19leIFo7id3r
a3n5KSQot7KP1vS8Nw0/QrdznpV4jWD8i2pIxg+rV8FZjuU26WOsCGsL7UVU/vT3mssZUWIEIQxA
qcgoU73R4UNWe7Cq+qp5x06OuLpcnpWgAb7HI/ShiAyUx38WUvTRhbWNKg9ixDgSQg5PRFD97uMg
upNOrGOnUuTNp0QEF9Q4qqvFG63BkF1KzlXFnZA6mtLdqxRW0KQxHesf0VD8yEDtthdGIM4E4yjH
qmcNbXRVFRruBdEDs2IdsyqqfG2SGtoomukBSBG02c9mtXZVIdR2yamcrnI23uaC7uO+o0T3jukJ
poPzJU/aOnTbGWhtzBTFG1U5JCFPHiDoZ/DsvFPmn0QPXL8B+NJ7zBOgMsMF03lHdI+REXMtslO0
9DaCPMCXMkT9aP1yhIZMZoOGtHXNBOKUJonWoc3XKp77QZoyFe1RXMupzyObAITiMBW1+C3oemEN
B+i2kC5SfPsBd8aeACfuoQWnoTUESTGskqbbF6jMxBIgu3ktXWJ06Y5QV/xkWmCXynFz4xeIUrHd
kGmPlwJybEo+7+HBM5qzuYvVQZ/leUl/yT/GFiPzoFRtiMRA7O15qm2PI4lAwzMeHef9NpVS+7jq
n0vOnXI9d1G/g9Yjb55kaNpkTxbKJe9NsfO6ZYWuBhqQSYltp11qtkUT3DmH7EM1W2A8Uwy3zkva
zKoQS5nskCVx2eXEAVluUxVWNd7AaSN3QQHzzRziEqVX2s6yucbxbeHOa6wZVk01fIhxifzdQUaj
6/DtnOT2GKnhnNjbKlYSRwRQqpvGDSYARRrfqF+R+A2hnH5e7asoi5zS/UnDksAwiK9/cIup3XkR
MdjgwrEaJwC6t6PPjlcoV1ZyrKkStylUcwmPLEpiaJNRy86pgqj/w+MF19erK9DyrSCm/ZtPXztA
qUMv1mdbROAhLug+XbXf3EOGSIc9kHs/Z05VqnI14NOCZO31P/JcULXaYNQnHHLrM3gdfDf1TEX7
oHL+dseu0uGcrHdWbN1Zxv7U8ZDcvkL9nqzOLLDMMHuy5BxaWHuWM8fAlatI4192xImSmw3fHJnr
RgjRyrq+J3cT4LjYn0UUM/H5Mqp87x42oCV5srf7lUMHwAhhQZZOnDl/T5vP8+J7r4RpPJAqzA5V
VMxce8RWf/XvLUNde4hXwtmU6PWQWHs1H95sTbNIODBeGjlpUBF839k99YBxTuVAF46nTXVuATIk
WL6gTLirNAhIQqP2wzqiA+FTFTBqMZHmweXCHLhGpTuKdAZsWn3kvXaeVVj+7AvKFiupQBrGvEY6
+Ybw+iMBVZPZBBn+kGmHldyzADIUsbaEAtjiXA3jb8aGq7YHz5ip6WIO4TAUg2Fw5ZIoDTDuZUcW
o2rKvr8PmkAjaaP9nmK1PxAz0Dh5ozaWOpmppTnnRNjDc7LmE6XbgqYX8RXxdRlULJwQTyOIDtbJ
wZ0KpJL7s8q/YjJ+rS7jQEbPg3G5OgIAiTA406MHFbpuLc0fJqIv3wezfTW7KNKOBcLbhRtjC680
mqOjKXYj7SZebErjomQJX1qY4MmA0QV8EP5IzZ8X+82wc0wANZJiHR4oywC52XEpqyTul0iKJxaH
PZ+me5M1l9TTFyCCidNEQwviO011Je8rzz3gVtuq5XuSh/ZQ7aFjPH+iBU+2YxZzY39vEXlj4Caw
dVNo4zFR3ZO3NEHA2/jiyGGOtFwU3/iPMfbAp3V4D7C110rdpiYSeXtw98n0tx36A6Dpbw3i1rXg
cxuzMIS28rE+OlwjrLqVM6ITttqmo0BbqdrYb+abU1XGNpFx1BoGjPmIBu94XsTXQvOP2UKXaMEz
0d1pvbgNM4U9P8eYdpq7o21Fk2u/1gkl4G9vKHzbJ31nLAiadoHWRP2Q7o0ZrM2N6UscqVP/BBmq
hykp91dFD6RlU3mK08J0tWpSmIs95aCOswz5dE8ZKaGuoeWGUG+u6xD1IwMo3hlGZvNiHdfJ5fYJ
RVBl8/IeMIyl6G0Eehthbyo+sBO7SPF6GUuq9lDNK7qnO/Tmb9CCiTf42xsKtGeqTlHG8hAvqgC6
abb0QYFeLN3eZnerb05oIcr3scUqKQ8fbc5FrTmskjwMvenKGywmoAlaqo6kYAmt9OGyCv+b1ua/
TmTS1m4AqTlSBCG1EE0YlsHZWXQYHT1CB0FfBtWySyLI+CxCQSHovlhaTe12h6TI8GbQff3T7thC
Yy/EgEWcDPEDK4E8ZrgDkuwMPTD33DznlAkaASdUsLRbQr6wJUPowqdLj4Js+w806Qdew3mtLw/b
UlXi7Elcxdnu2Olbq43aA1HRQiYZ3hfGMf3XhMgg/7mFNgaqNRXkS1XafFH5+agjpts9QuFAW+yO
cx/KNsMJgi+LutMffC93DlXwTwJGyv3O50rpsMtOGab3xLIqR24Fy01L5UxdOJwt8MG37jTa0KAY
Fig3+dETYHB+mAY5AyTqjyB6ztXR0cHAdK573x4Xu4xxr4lB0rW7RDKeqc/0bCSxuPTHTEBWwN6H
fX2DeeDpuZ5D10io0Z+o0z+Gt+EDsY96OMXPD/YL2Qgy1YTEl1Lx8NtI8ibrSrgGU2wYpeU5F45v
pU6yUsvXPEOMJ0KkdFRjHgl2rLx563wDCz5Jf3HXYYEbqgny3c/nUAMhxWcuFC7LCm8pB9bawnHU
09ZpSwOp24S39wGfllycjzecPgSPvOxnYcjhcLZiFIQX6f7ZyFDVsQCBstmg7vyhFkJwHHAhPPgK
68b5ma+WV2XCXoRWO3maERfAevCfp6poHl4tkcOCFOzF0StxS4uS7ZOTiPA6vbD6Wok3UBPK/7ES
JlLS3ZxB27hkk52038vsnZUF6+wWUBIaZFuTQ9hcfHto11NjBjf1TEB2gE9J9fd9vQQxw9ZOhLVN
um88gVp6e1cTrnE2Gc7+V5Ye0JGMmxulGxkmhQV/TI+pBSGR4Q5u1G8bFGDMTY/XYi3QO4I2c+Zq
DgsTqZ3iWOjBQMLYiUxzyAA7rrLScWfWdvRWgEaG3PR6QYYBjUBFBtqkZ+aqqUw5FeLy2hSGnojp
voXL8gehrN5ziM0I/ytWxMVZZC7yDLnMTexlK1C8PafCXX3D0ht45yo93WP8mQOxfqXvMb7XqwIY
uxaph9bIu+3S8BFf5/aJTWGMZb4ykZDO0PkFi5ageygR9SvFX8cL7hTRhn8hI/24x+k4gmNL0QsH
SVPgyMhMYJUpBtUccNXKa1R7UKkBEw29TKFqsDaAEFFYvoLOCpooWZ11gCqX8T+72ifKXcxsglSU
ama8isBHBTHdQpEnemDkZFJITXBsJ1h9clwskPohVHOTx88O/ZYgffnTPI+q4/D4GORzvbXm++Kv
YmpRmeLrlm6TKgQt7fM/qL0g/cJ9R26Fi31aL2SUBpYS27UbRElKNaVqzZXpmnoFfHSdI0ntb7pt
neW7AlRBs+nwOOA8FLTT0cTgOkv+WjD9C9L9mswGDD2oyc7u2AY+3yjJNCURqHc13yM3jyx9OFW7
MIqITqUXLfDPKepeyljemGRlFDpTuDI6IPIWYAy2X2TscvGJg2yBHti9m5zBYTS9xjMkgQApqizu
M9zbuP1T8MbcRMF8Qvhp8vyfdEQspOw3i5qFmrr1ybNfLtnZJUX+QGw5LlILo9mK+L/WSkfw0Xo1
V9QexwrhSZPnwCVNAb3p/ExexIAyn4Ja44Vnsf4K9oQwv7CTbsDI/RgZi1AlRFbkkTI3O9+BNleT
1nqPNiUGqpGgNt2GySTjcubb1QomeoMX2ezoVba2Xo83x3gTbU0Mj3yAYDHJqtwMUPcoppCNADsT
Ob6Eueh3Bj9sZKrTJSjTSfIrjLqt+HqLjr74/+3HQD6d7P7ZNu3JjhAREUnjSB1WdhT4LD0Do/kJ
jrxOizsAJRZbUhnyZi/PKMoJgsuIBeViHRkq6oTbYEizh/sS4hneqbmevWnmYn8FApAFE9Y0ueyx
X4BgAZXX7L2QYOcZ/UubfivisIR431H38XxkaLaHOp4jDFRPzDBrL/yTi1UiTyfQagTVO7fpLF3z
UyEJO4U3g6Mk9wkbaRoDYe4un9Attdn9WUXGn4ULbQcQTPvxFiD1axtsPVVZDXbUbSSWuzNAh4Ho
iX+UDtnZFb4vw24uixjXekMz4PNd+fpWbnY0GaLYVNYsMZVburOWtD+/s081+6UsHkIvytuT4+XG
34E8yc+jOQxptA0tR3T6JRs0ISd+GDshUEvfH6POe59f1f9rrqR9GVYPlgGiPb5Q2j0DX8UrI3Hl
OL/Mb/piPVwSZbzuUQs7UEEeA0zZeeQxuSYoovtUKtCTQ65dUbCVygZEkB6E7Ytxsxi0FdZBnsJE
zC/lu/Ogfgr3aFSKB5FKfzwcHtlBIc2gXzfP4GmpYh3Zuh0OpMovs2EKfJtX7QNjjv7W/Gy2EdGz
jrIJEzNAXIKejVudF5S06ds0YpI4GZ+TEzn+B3zp/H/y5L0AZW4fBQg1XSgZIolHQOSKGaa8qRGB
dcpjer68/7duJ5iz+iZt5CwWj/DEJHrM96zK/Cch9sPxstzJAb+4O/JmZeCmoImqw9bBp/Jmk5hp
pC+S2FKuZ3rEkmnkPW0xBqdzkop/Q6dmxI/PxstizmKdGwmvpGlS3XqAibcDt8qA+P2DfHFSecTV
6DOE+uF+JuZCNn8/LJ2qFvaAXKyiDs/4AbUXGmQGdkm+uPSKVuo8L+7oq3ouyrtVTiW5f5KW9Bst
m3ivzTI6l+y3V80vJFam57COrycSCVE2K8xW7psxltLfBmNH1nmNEM/SGRGwhKWWctoqZSR9U9/1
Xv2Mub+uEMnhTOCPaoGSf/SQ9lrw83WbkSgA7wDpOxiVxr4wedpzevvVbb/NzTn8ibqH/liaJWRB
7IGvWT5eHLxCS+lDmpUqHbnqCky1Pdue4xexdma4BE/ZeXCbasZhmv5OcTjBrmuDbpQHnFFhA6tv
O68KBWU6+XW40cZsXunocYawelvb699OXCcrYDg1+GlL92LtBFC8hrJivD3R41vX5i8XpQ3nhd2P
Fbbi5K+r1NAuUYjXT0fCJbQ+tphnThvQHtsudBiApKa849n6OhrabT/YXjTl1A57SBF0pI7UsuQZ
GzwCtWVTQErA0WDtWE7sCO1NSlqpNQ2WJ+c/P/KeaDou4MnzaFGTFuVcuIxUYO9V+oDKEuPFLsoT
9R/WApK+E0cLAsYHFsc+xEsMwXgjIaqxjKMBi1ZLFAJ30D1Y+dq0a2neHSSg7TyHuPZnhDFBZ2uy
r0sBHOhImQsKWgdyp6481ZflhSkkTSwVUdKCdFNhOuQd88pt6DDQAJkfRJFibvwp3IxN8nmVOHAK
CI630WcT1pQ656OqMIjZmwah3z7ehOA0sC34U7dR7WxhQH/OJGkWl/1iw8uEpueE/719IqN1vvLX
jXWVDZX+6nbT+U06ZBcUcRkqtEXi+5QHWb3sMuIAjqf/V/7DXg/R4/1rMTsRlndYu/ydcopG8zj8
g5JWiAZdsVcTNC5EWsauWQ8/SsLS3G8e4NclBwViCDYBQv2C331HVJN2tKsUy0ITH4B1jk9zT0At
24ZqxLDs17L6T77o2j80HETb+w+hbiNc0AIpMCIDq4QiNAMYqPwE2imNm0y2/N69ELjAYHr1L/ug
QqRfeJWMjpx6oo6lgQTLRntEkeonlw/Pw7DfKGataeEyqe5/gGWxhZx/Suw8K8b6duzOrRQcl4Ct
nt/41Q7tcRsnhhIn6My/iZ54vCipeCtF8xs5u030CoGPg3687A8Fkckj2fM3FnE1ZfC3hnRWNy10
FoKI8KqAntpU4MPmb3CdjBcFZWDBJ3dZJd10nf5/P/Few/BDsP//GNFtFsnl8t4VUeGcyVfCvCqR
n5lfiiiDG/+fz9oJsxndVcBidO7sOhgFnOia9Qhd7vUgEeYlGkGLe2En6eGjKo+u4630PJ0wPeT8
cfaKwg0vWUOM6qaIC5q+2v7yj/Y7HBKe/f3qJawDMSD0MARRR0nCg56JLHOvWqN3/TRgekGLFtzt
tw2AUEIZ67Nj6kN1081WgPfUMIT5PzHAUkBnRKWjbTdxmHuaFiLcVYEqEqYaT24plbECmSS0dIjn
zd/A5xcH16fG5Xg91ePzEi8Ozu97Rp9Q7E/I2WeZ7/OCAWphNo/yi9kyzXhc3sogIo/9QNm1vsc5
0w4nzGHI+1DMGocr9OTmZnf7I/fWEZtHzcI/rIrjULOEMyL6Kz3yOCHWZGreBZyaI9nP4cwbLIBu
fKhQTBZNlLOErFpGzh3P1B/PtPaRFk/LNSTJg5cxSwOdNFpZ12KCmwEZRMzIQAc6qm6E9xuTu+Lr
mG6+H4QkZbt+j6Kzdv7nugi0hUzHw3L7FQcpIiQ5sSFQ1P670NOQYxPAMJXwx96qtmJfX/tGCOev
WTbIJEIDdWdCISZvBnr7itnTavNvkzQopxvdkVZ8m7ofc6G/BUIsmB0GtTDL97IPWZo6sNmVlrok
akwVz3SzGqCv5yeaEshM/+oN2ClH/n047lW/gzxyyjruuazeaG6Ecr5trpggcS+svFFH2HqxdCEj
rvJvNYJKdSg2ARsl47uBvQBiNbr1HG2jNNsU7otQhxje8apSm/ab2GC0H2WATO14k3R9BX6yl+aY
9IUYtzvYQHnsXDsws9G42A/IgMjslwl1+5u3+T+eBJmrZmzn/GeQg2jBQrSIqmAUidIv336NdvK4
ssU3pAQE/SmXrw6LDXgjc12XnjI+p5lKVuhsFGy2asJT/U8f6wNrG8KzOhLKnAuNAeL1F8QV0OIG
ekzsEPYbNrb8MqBqrMTBQ6X3qANipRXgJlbpyZ1RgjxVvkFdv5p0MfbiTHUTH9AJRbzjP+BdiJ9H
XOuZF41KG6XYctKdZFh/Bvp1N21AUSEPHJK4Xk47SeZEhWoDMdLr+pxsfQG27mUfgsWP2Lmuees7
cm1y9JgqTc1Hop9m1cHAzvVbQkL/2OLO0RvieCjQ6vFD8yEZ7Xe4FHgFxb3snxCGCXNOXb4EsJ/D
VmLLL9Rw3ZzVbu7Eil69eVG2XJcFQBbsO1Sp8MCdyWfUclAx7fsoVSkP3lEnUvXuTfBN9/xPtR6Z
v4R5juoVPzCA5IYNPoGWeIUrqyFdmKN8dP/hHQ63UcNZJ1yc4wW9qWPgSZFzf0t+X4BBJzsbo6Gr
z0PW9nQl7IJeBd79SzfD27jBNkQynRT89w622GcrlU0eXCdNiSE7+XfTqHaoZ3aiL81zenUxX3S3
rf1N9/RB6sWmMzsyurcRAWidtj3kdy0PPG/H0FnCVkMQM5kkrGvP57pbwiFHHHJvxAz7nQF9Thg7
RaLIgXhIg/dd3jplUKBD/KRlJU+M44XBiO4Dfb/zcUF3Kz+1MtvquYDJPZmpL0svEasqp7QrrpaN
ldk0Un53X4HYMCZu5o6Om7qFG5HDaXEDTwJUmQrtVlPp/Z0Anl8A4ipADbOPrGaxnOKi3bo/Zo+E
nT2WZYtofVi7KyLxsEffC+xG4y1Xfx3pwk6kLFEkGPZgqqJZtWN31Ydxbk2rX3oBiUJsnU3R1mdm
uPTvcq+usAXidvxsoxZoGYKiaXGQRKjPB9O4IB3cflwu0u7qZZJKhbwMinXwm7wBL+GP+nkdp/9W
cDOiu85svE/Ifok51KB4Hsbufuhj5CwI45RPupYJw7TufisZmJXUbZZoRe2goAe8Skx14kSjIAnb
uIpTOdXYQ6V7+6vsG63oQnLbz+089iAKCFpyG5piT0DLVLyYTagh3rOaQ12KR9gr6lnmKMtPZvwX
EZJL8l6IoUj5w25KfVNEbzODysSZJcl5z1DXp70IlWKYH6zfPqFlpSRAYIoParCaccgT/BBm4WDE
HFt1mP+ECdUF0tsyOkA7qhETS93ZaNAu9YCvF2yRsUlA5mA38Ui6JBYUmx0oqYzI8vWoEaRzwtrW
ETma1Ejz1BhargwxlcR4K6BS4GrQbsZH7XuLKP1oTk2LF0bdMVaLk4c+q6QIeNP06b/JENkJckUY
ev1mJC6f8SCeLKRDPiE/bNaHTv+CzSnWjDbnRRpAhHyvm/IM4mz9xlMu8RxpDxuy2S7y+xVaR1Ue
vf5NBhXDO6rKQiPoqrX+krw9YtX1+pi5Nbp0FwcBcTzoTx8zEqDNz9NSjrS3w1U30iMuQHbtYVWD
gNDeViENhJpkzK1wILgHCo8f+vmm/9AjN7VaGpeWYKzT0uUFg580VMylfnf6vAE4QRltZJsgOqZE
LNKZqRAToDAOutJx+4JN2JA8IFoKnqfrboOT5J3JMe2/9O8lMjMAPvf1pcwL3LjtTzge1wFKOw46
WlLBoQXJygjm69Rnsixa8HszoxTcMLPKtOVkMzRL7EcTAqcvTHE6Q/CayZTQ/jpu+r3R1ixMa72X
eTkPmlEXSwlBIsk+hTigz3pGk3DzGvbRbqsDrDZesBguPrkMGDwX8j2hf8rTrBBDTzERpwiQRZ+9
XGWsBS5ylp+tWtrJtewJiqsTfnaJ1+rc9qyXACeVE4zDxMSvcoym8InaFJSxJEqiL+SDqkTYYeTX
s+wmo6KZDWI0ONoSuKFIZHbjPwiqdf9siLcOMhAC/4FDl72r9cBLbfmMIMIa19wRDx5hedTsEsY7
F1ii4fggwT8+UtgrOket4G8Wlfg/gH9wALsktPkMxdM7Cbp8AHh8rhufoTj4FP6uVvO6g1KnC6nK
GqjDW/y8KSQAvLS5ZrTkU47XmYbDVUEy4a5GHKzxI6MMtQTsDitZKUj0j+k3VbUeeUMxhJJZjGo0
d1uZDOu1ZWtvjz0ZoGSK8lVg1hM7yvBBb5rwZf6gnOmyhvyH5SRBLlVd6/XSH880BMt+/N7dxrYI
0olRJiv1jNsKKEpwnmyOd6B7psnMexQlcaCTjc+jza5T3maZBI2MdNHNOqZaEQj816mLz9DLQla3
t1NaFDlmBPU3HRriN8eZMHjyBJTF8+1d7kNO5OzHy0KBQL0Cztmv9+LXHK4dDYw7yBQoIQvKwUTV
O8NNRlN/WopiyN3+8Nl4DGhEayBjADrVgnrA0HFm9ZOERFmLOSymSz8lpFQjUqkTLTmrwSLx4wTd
SUOhx7Wxz8O2NbbcTdo7my6jHLNuUcZ0XZFgF+TrO8xh67dKeMtO52WJm/DouCWQHdgTWppYiqdC
0hcqxiyWDDxtDDHC52Yr6ql4Z91ftKZ22FAMK6nH9x3V3SqFronxTSL5dZaXLxxnpU/ITvSx7b/U
H45TtqPICK9iOfwPicDxST/M9IqynV7b56brg4rxaPLntR+wsbyfqkj38RDTm7DWYeKnblC59Chc
Wh/6hViYua9b9fZkstJ7Tbdmdf8ctFEG0TyuiMAPjW0H9CFjqU+byeDOYjlfbzEbqVlxkUnJpvpe
7WnGQWd9taRcar89dIzTqHYTYh89xWat1t9ns1Skhi844WqGA+pCwjsuPSFWp/k9O4t/O1clUPLX
ubudHEDPzeqObQ4uORZIEw+RnQu2yjE7BgHKFyN4Kt+HzCuRWH0UmJnma3I6gLtDgCrUoDY+EExA
hoaDGGfZzSZs8zXg/+7vI/z0uzR3vPY2+4oRBYad5Y9dCVhBOXT0+quCD8F8LqcDEx9c5rSTucju
W156Wh7BogkzqSlwM4PQQfC8t25Ur+3t/0WpZrhTZMPqY3bl2AMuggS7Bn8wsUuB4vFvKr66IsG7
J3eWC8LKW4JMSHi18ZBIyyp4Ag0fTPGh4kqZ4Re7BP2M+572OJoP7dutFsq+2nKrt+DWLC3JzE9U
2/i3sSWMHDSFWafN54+KOVYnyJgF+Rxu4MUH0AfHtlbBGCIwzWUma8sn7ZLQ2s9A9p3upjl1BbFR
nHP+dXkXN0QqIiPTmWQmzV26XT3Fdk+cjNvvG0TeWC5TTc07+yPmpiFzDG39ldJITEXMPyD+y7lk
nLaVZM0IhPzvIL/r20E5r7GgwLwH/EwHOXaEkOYEQwY46w3ztb+c9Tvydc5NPp3PjEVG2d6M6ojf
Def2+og4B18xsk10v/PCVCWfOtQ3jiGyqAuqdB1FRuayGFM09R5KWbUE3OE+9Lhby/1mEjgMU7zG
2pX+3vNQpAqluh6QVe2G8dsVYgqWwMe9w8qvTzhOeAiWXt3YHPCC3ZS1fIldz0Fgaqbj/fNq7COD
3dyD/r8aGrtfnciBLwGzTgCggm3OxBK+lgGE3pPXCRvjW1GeWBx193+qvCTjj8UarpAShOYVunly
0ZUVSXtd1nhs6/5qFxgTmI0DxkHV5WyeWNGF8UzA3xPJbJ64CVUrDiC0b40hnerJPFUIbJHsk5J1
P/zRqfmMWDdD7NxqyYk83sDlIXu7Oqu8nWOw4hZAHvFrMcIpi/V7+CGnln6WB1oVjRGGhj4AP2xo
fqJOkaRSYsVdrRiejTvCcUfZMZ50KMKNbXj1oird2lpMAjfkfOKoGuMLFCZBTn19a7QkH4uR+NuF
0wZv5t1u04G+Ai3ENJJau7Rpk0tNB9HlPBPB023+ZmlMNv6ZELPO/r69J0Ya4U/g38uCvGcsXfOc
hraEb+4w5ztqhRJcYlJ2BY3pzcKl/hhJbX1ErZNzGQ+Vt0FCdcLZhNu0cx412I5UZRWSupE6cdH+
MWIMvLrt21d3UL5oi6jZALjS8WXS3q59BdJuzCQnK2hu5IrQqbIKnGGbi8L1lkdJ8/OVTYh43sR2
/5gQr9kzFMvNldLdCoEeACIBVd13fJQpA4IaApfNT7P4LRAUigdIO3EBGL2Nwk+tb7TYEtq637h4
NtQyVvXN8Hbhyno5gNSIaiY22dMnC1HDouXhy1r84ayrsKURqDBjMnzrskJYmXCk5jMb/9yq6Bgf
7WEhjI/eQGcDH7Edr/9qftI0oibFtEFhQcau2dJHDfrJ1XYV1xprUqaKLeN2RutXs4VM0rHRPHDW
/n5TILsw8UE4TYPk2udn7K13wphA/eMt7N6KexpYy1eskawx73vhF++6EmNM6D1IpgoTwQq9E4/R
oIoi9i1LFMz2LbUBJgmfTogq0rff/AyN0xRQd/ChZfVb34xZ7Wa7FtGHGthwM/s6VUHTXYZRSkJn
h0Bjsz4ctzHadkTMUCnfco0Pul4sC7sYRt8lgFYGNCCricgzyEQqtsFm9avIp5F/1IW9+9SUdRGF
im13uXFmjENBpnoy5FoOhMXehEYps6W0AyDVc57NgmIOpDaJDti4mwcgsreZwxDk2XVA0kOA5jK6
Fz395z6yy7BAxZJLoEC9oP03Ckz+nh00myP6iB35muKjKbu8apZ9nn7VctWMucXqryjvY+Oazgs0
nqkVSJHt5cLVJrZyRUAlsv5vYx1w2pHcgSkQuqMrQBGf5FRpkAIjrW5/8vAaevizt5CynTi/uKRR
L5R+uM6rsq7C9xAsZhDjljcGuyg2GpMb8eOzvFhGIyETwXSr9PYwvm5+DD3Nb2PJiqzdYOVPTEA8
8tkUoU1HL2U8QWC5H0eR1Vf1DmhsbqcUNhKnx3z48W+opD6G54m3UiGhKtAUTpRac/hJd7DOmmOt
cq3f/585zAxjDvJ1YrNLyAsVFjiRR6qFNrA5q/LWf/QxMzaYFDffkawxElKtWngznFz3BGkC4R4U
NJHa1GwNOE4BR96z0YEvWm2Ark5CJyeC/CSFAnQjiSkqHymQQ16h6RrVzdCUf+DfyyRzvosb632x
MB+m/bmpmpRtn7hsdpFs24iUcTJBLII5022P18ydaeFW5feZukWHis2H2qcJysJzb1O935TxN5Qp
LVXoSvUbUNDySIqs6ezQ7Zx/Yx6QH6eCHe3WgE1N7vs/P/UeXynk4Onj1zrHTUBVSSabIhh/x8S8
XkBvDo7oS/Dgp601tMZGDPDOSfvQbRokcUQVl+kA0QfR7Tz/MD3AUYFw/hEcjn5wg9iGmzzX1/Wa
Cym8Mm1NJBY/N7M5VoWm/ccugAUovJ6H2NaJKiiqy2GCMq1W66Ds6geq6C8EvSs1sV1rlK+pjmss
8JLaKpwbKiDIWr3jlHzPg/Jx/YlGr4SR5W/V+SEmHMGYhwsdvYxoRr3nigirkb3zd6tEz4SYN/fW
DOm9IUGHofGdSpr2aJKW8hO/3rbRvIFddr7EKT2RK9TbajFUzEYgSm0aeW+u4GyH238gTIlrTmCI
dYfPVMYab0lXJTLe+XER5C4HqgPab5F1yf7oP1IdQmni/tMfnElY2Vzqiqadu5h4g9YGqsCBhkor
rY9Uagn7THqAF11jSIe9G+nkSImDiONTfpxbr+lSS11fSVSJnepYM9S2CPGAyGzNFGPCI60+KHY2
wp5hxRfgxmjqByqj87BjHMOY5XqFlLedtCADZVQO43IOhPbi2vtM42Aew314G7FyK5kwC4/9mxAo
eNr4akVaxeEiON3yJ2jBAXRpF6lsfYmXuSh3lkQkvvLSnNDo9DcwIatW4tuJl2pLBks+orkhdvPA
+OlM+6kIAhcuNYXGUgTxsCFhfYy/CCNrzKaIzm8dtyYUQPMGAv2jRk2vxSBLwQIozDhURTR0lPvY
umIgak0VjxbwFhiUphAkiQkJN/k6AD5WNJ0HMot3CiEQzw8BKNONs1rXTscqCUJJamBNNwm1788Q
YPJ/X3fbG9zOOoIL1g7nJMVGGdgeSpWIjhF4zKW3u6hY3cMa6hUI3PhvSuRzo8d274r7NnhQABBl
Lv++PAaNqEOp63dyJW5NW1mU4QLnWgsNHppC3Hr3F6r4I34Sl1lQ7zDKB7oMNh5U+VINFgF41vRb
j3oKEifTqiYY6ozxMkt/dym65e+YVrD73DPsB2oeZ5DJeGOUXxfQAVEggHJHi/c69DKn9ulE7bCe
vMTO+Lo7YfZKpCIoDGUwog8SShF2B4RyQszWlxClPdQC6XSAOB2eMG8/YSHC3pf1/9tOigxUMm51
txHTHssUTejVwjQDzksAZHil5SNVGojOv3Iub7Jm7BGk1Zf6eI4BUpazMhPhgc29dNJ+FBO1YQRy
ba726n/RIolRHt5yxqKWHJQlrYn5flKLMMujVBnHepq/A4aZecjsHGwzby9R9RmFX5xRTlTzFtT1
LrYj9WkCtQ7/VaXJtj8J98vPgccCr/xPBaOL4YGNMMfDV1H3x8SVgTcVTitQKjcEc1ocRMFH7n/I
kCYgZNwv9yhhQczkmFlxwoCl6Wu1x0VguZ9m7X2a/hQjmUHVO3uzeDWUMc5iLAhpKHE1teK4A9Hk
oUfaHDtfq37HL9joJpY8ajxfOWGA1/etLHj/hcGTxXgUqUBv+8w+WJjcdsDFLK20fJnmNJr6CZvE
5eh0/ZDfoSebNpM5pOP9CiTFdFhgAwPkUO5y+RYJQargHc4xZut6VxvT4NR/+rwQ+4TFJAtLqI5u
JHKO+v3UK68+DJtSaKOtopBf7d8vNErylw8Bw/aAtfyIZqlAAsUArk70Fv8aPNst+kziiZ+qN0lz
nvgTEzUcIWef0Rec01SoT2Ewa9d9vlwia9lMOUoVHvTqiOGrSST6Cy7gO52rHuw/7hvWqSz2+dCO
cqDV11iitIfGWArCQXMdc+nopCfeLlJmbNaA/eGwPIlG2QIAfT9njguxFCTaNYXghSKh1fAZeU6H
w161Zn0RkpyslS8poDfV15lRo/0UeAhw+lcpfTXche4Pvteom0gd0eQC0TA82Xf89NoIaDNo+0rz
g5OJi1v7mf2gGazsAVpa5AdRsG1AJkcFLVWbplOIOjZX8DEOUy6hCPQRBa6xXvUG2sdxzUaqqER4
0lXTU6EvTqFDOOgroXZwMySDAbt/UJ7IwXwe1WJ+5zNW90N/zejUMuf8eZyZj60iHaqBc/QMF64D
4q+Ozu1qWEV+2gg0EhYK+KlxCnLxUi28h+grcvgdMXr0AxFtbwVe1G8x14YamfUDG6p9pJpjclRr
6n7oU9yw5xNQN2Qi/DGcrveTF6S78R+I7InAs/pqJTnB5BscIA1GwQ6E2XAoGUgMkmT8cNUMJ7fE
3buTgQgNXXnFKPL4/AgvQ8KagA+HNqOa+wbVzXXfKUZ/pPjN4Jc1UovIC9bMBy6M9PMICjG1DnYB
g8KfUce8wmTEpZD+9/eojtFKn9EiQDSJDBewGHutTkl6kTw1iJMiBKQnwC98F5H+ZdHQGuAso8kO
Ieh+jGP6DUpeUyJKseX70OmAw+nuXUuG4tGdCo3N7FhIybzMpUi/KQ8nckLOIRHGCy7JYDrpA9Am
ikvfUGmfSbSNAhNuC9JYAQTlgvmrwy6vkn0nfBB2Z7V/p2XiYT7qEqK9S8fqgns7esEBK7FcAUMh
ACiVceQXptmloL3rJ9kDskC7wUW8zGw8qBOqrqwlRz3hdYeguPsZoFRf7S+MS1wbG1oQtDUPcl0W
feaOIFz2X9QSHyneUDRuNAP7CyD40bRLqBhCptOsG4+B2aSm8hjBvjL57nRMrOAYsoD0f2Aq9vp0
ZK2x/wGgfAD9GVfMNsqOnMkHeJnrq7NJpk+jRw5lani6ckdjdSjYvXHYNLWiBx3dx2kDLkc1MEgu
KNQMdqCYCHlSPl9UjcbdsCa8bAG2MrCFZM1QIO2WYND4ny0cPfM7JF0XUOyhBUJg2octoj7Fcf24
IT9RGDXGQhDX/qTwVR9wBNphJDzUCh4RnMAVwKVyooJKKSM7tv7S3oIEjS7fVYk7bJvwK1Qhr6fA
RlnyuqL7S2rkdlDqRAd/RAQFLc1QyY4EuU3WoAF7kv6eMT9OaUAxs+hK4xHVEdeVmbAQaxjO7X2j
/XJEc80LzgtNn+UGorbxwD5edzc/deV3uoijYk5DosVFqC99gpva5KJm/IKj0nT7GPyw6sEsiyPc
e06frg5YEH+/E/C29FsN2HJcSSe6eg9ddwz8g7hetLu3BCa69V9Xo/rlObBVbLqQojUqAEpUTpss
bUidTXHg8no3e0yk5Q6EU9HINceNsrkEGL0dnEUquUe+RD63acOIxfg9LgWt1c4emZjdOF5Fps6O
/jKNGgpBMo2RgCFphw1dRW2l5aiGGNoRHJrR6ZCrkLKHHd/JS+yRIZwA/jsva258bd6VlbMfj86n
aQIrmyau+sUP7TGrpj18P3gFuuv0ddV5fG+TKpoJmjj9E0YBSslm3FF0jQ8ganxc9fKsT0n//8T7
1a4AuWJRUTnRDLxaDoPNDc1u4w8IMxhBgw0tMW4QT2a0+uupFqhAX0jYRQW6r5IowPaopMu/+59s
ByiIq8t9TqiiveDRue/twlrSgeyNMhWXJA5btAtGTvsvbKMjQpGkVc8MvQegYoFK0kAtfZ5Nkp7f
fuq0/RQKTERvn83Yt5tClH3Sb3OLZwqlwycRtFdgT90H0B0eupBlkhWv2K4iFv9KvLnr2toC5amf
AR7i2ff4GwVcW7pkSABud3dT+9HyFot9dJr6Qxta6vdX676QKG42y8rJWgwR8Z9otxkC+5QZ4f7S
j27fBSJgZ/Wg+cgKc8UrZZCg9t4UjMByLku1sx8ARE9AHJt2+9DCzSdl3h2qy5Kb2qPQaGuwqkkE
+cGeL5qPcJxIb7eIQQW38F0sbRiczz8imKz8AjX3fkNTf+oP9pkEr/Swc9+jwXGEdOuRrVVaJ0H+
0aH0QoTmcPwHg7j9z2rkRz/DbubzOU/bXPiTLQd3r0dtYQS6sGrvFsJJs9rCmK2ZmnbdFHaJS+sM
DPCwGSy0G5wWfMGRLdM08bv7ejjrgaQZWV7RSl8NTEMydbxxqQQOb7ICu9/7vXkxoyet9J8dSJ1L
vgm48/tpRZAkBuRrWiBMLKPjKzgUKegA5mtCJBlmJ5uHB0Ero0H2lotvhn3SYcuJg9/Pjx88NWYU
FEWE4xTgVsBI4l0iSYlfnbzOMTiTTqYghglQwdtDV4TYM2CwcFKkGzfz2pWsIOS4nfK7E1EX25Jd
tLD9iLEj1ctyO8fnllcs3vpxw2oCb0qcvdMY9mvYFtD//BFv/UTqISgdVgLQRVZ+Hn0tQmOE/x+g
EDT/v/A84JYAC35AZy8CQmmfrlfshQ5mCIusNusQI8uNE+gWbdwF2CuZ+Mv3J3Qg1fjWyvj06Q/n
8zv2ikoShjXgUEXzjhzArI/HyCTPobHHw+cKbCjQwzunFTQJ765raI/dD3b4U9MbWm+qwEgJe//N
IvQ89QBftDMCbMBH7yGTu4W5SyatVeVJD0b9SdPB7k1ROhzZ+v2Jw1Lt+t1gYX4D+wZGqUNRLDFv
E1CoeBJu4Et47t9plVmMSmQUKSjtSI9nK3StirlZIwIv8mOZceHtyXDvYhVPmcaoNIs/2FwWEHm5
gxkFAtdJO/iJes+Oo9RmcGbNa2QES5Hl3lVP8vl/FU0jOA2YPNeAOVYUxo7ggInZdz3scizPfr/v
yOkVIZuasK8L0+1YiBT3tDmu7z51EnAt0wLkVTiHMWRq4pz9gW0MRwKY+7tR8CHTgEvGOQ6s/Rx9
m19BWgD+97edNhVi4Imei9w6+Yhm84M+NRYF4Q6g/hMWGX+euAC119282Jl4jujN8nkWSGyap3zj
qovG0B8SwVNZg4An3Ke4i6aWIEWQCnl+90rhVAwsV63YzjBt9hzsMedvngzq1zoYfsECGiTW7TDd
ZtZaC+Ze5VptBy9WgJ5tBxAswmTfq6aUhbd5K/LoGBDlNF7ZP+uIjgCXHCDZb7fVACagCkSbyIPq
qa8jgO7sLVG5HWZs604OF2ZT3GAkcBYiiPRNuwz/YA9Z7OvlC8J0wbT6frHQ9CdfkiB0mDs7oV1S
HzkZwxk+fkDMmeNgvCFST8+Qzy8MejeP+6IcOoRmfHS0f9Z3P5oDLFawOksEG5gB4Bx/7MsxVhKK
B2tsyvPufN1Gk9r45agXj8P7cD0wTdOSR1i3KDp9eqel8z/HXZvJJQbIFYe3W9crnlfxiQJ0aMEr
uElDhb0BJLYCy5qLZ9YSl56oUBOlL6K4XYL2nGoUSQKAuEfsabDLCXRXZsmi3DmtwkJs2DaJR+Dm
sBt50k7yMwoDcq0mZaMSsPxpHRqm7SwAGuKbFRLMIalQ2hMxekJV0UJ/LT/8XsX39U87ZULVxDd/
3N+77Z0w1lzKdr4Cbkzt8wTLJSkKgUXmwP5ZUJ141KcIb9zKvXNrSct4GdE5mW8a3T/n502i+79c
Q73iD7P7aDxkUsVc5uHCIKiz7oHqcrv6Mu0HgzsJ8iwDBbeWmyLYeJwdQmmRMcTSs3izn3cvW5Xc
Udg/rSyjS4hGvhleVAZP0zeGoqiM1HXKSV1Z+KpurEcDIrsbEVUhgPhQxhqC9GB9vkRha0VYfZE4
Bl0uK60OGtNJuUqs3a3Oyz8j6T782f+l6rwe+J/tUpf7ye2Dig/nFKL8yCS2ZBb73yf9u5DCh04m
9bS1QBWQM4e7MijGi02SKs0W101Exnh5GQ0pMWoAcq77+QNW12DER2s+Aoy542+D+TslRz3QMv0w
EnR12C1bKjNFJa3tezzHWC1wr29hRyw2mKf5rBqd5VTzJ+5xzv52H8Z37RAtKM6qHCI25WoTtrDU
KgrqZop1YSDHLPACy/Ion2ZzJh4wZ81Ogolr954pnvRy6SdzaECi7j6LLzfFWAeO8dLhmkIqk+jj
dkIQKMWGUbUgWNWd77i9Z4qZ9GsDUV+SYNfl8xCtdef0HkPr2PulVPbNka2Ew++eYFegMkvgBE7c
WzeiGcxZA5AvjOrkrvRZMZHVnw2r27JUCl0r0xAv/yGOX+8jnlP+Tvd2RogN3qdOkBp1syqneP+6
DENTpyT1AeqyGRgp2evLr2lWLfj6OvxbUVBA0Fyr/d3Q6N7yIzbkInwxyk/3lus+HWXsowrHQ6iP
vyqgdIsrBp+zJeq144HvI9J25YiYCC8QLNDeNMVAhGkEVMlZtd9NwJ5CBN73X+hwU8lQ8epVUpKr
OXnHpLspr1HcFTX2j71Gegz9qNFFFdCMY98jS6nqakO+aZxPcGgE4cBp9x9Zs0RXdd0GCVHNSGTO
IJGOpTmg1DnmcFe70fMRCE4yakeLZ2mGhriho0sao1xgUo4y+kjD7W0G1jg/56Bqzx/7s4HazMuE
aBEh2jjJUlngpKlPl3ve/W6X00/9pQCfwK1LdzxMq8A9H/EO1YT9N/I/xAXVZyphb9U52/jwNs90
+RDrEIy9PBqSv9PIHsqGEC40vfvGkBKlGHxykrlaPDTzG8Iul+jGTp2yBYBr58IfksOU79CSUAb3
rovFex1s1XyxXBvlesm+pkpfOGwcCqCHitkU+ToBck475tSiNgTvjKHp+U/8DM1xe7Puwn6VxS32
N7DErLaaH7A7lXmF13yHIny/sA/ryZ7Y9t49zHa85A5+CH0qC+zREAHg2DSp/CzbzpGWffgOUCo6
qcyr8s9ATk1MFcFVU+e0pQDSS/ByiW3fXgYy+PJyG5zf1wYlMTyWEu6wNKFaMukJe/rx8HDDoqX6
J4teHXCPTtZNZBm6ex3JULzZrAu+g2jxrytA/D2H25NhEOq7FxAF3DFs+rQgL1/SzVlFA7CW8tUk
eOAH0DbAVXtGk/UWaxzMcumFN5fj/poXM4Fp7YCSSfTOEbtGoJJPorzDVLUynVsBtT6ItFUpocDS
WZoAOvsnXf7gKoiS4K1McD73XfjT0Oj1mEokryJAMpElgKUcgwDha71lHvbyIW1Y/uLbGswFeEvX
UOAaX571plBYwPsxHjvFqjvRKsBbtflC67Kr6SROt4M3Ea621YpwxHgX0tACWp82nJG97I8aTQRU
CO+JVXdU6rBwBv3qyM9qJA1iBXmRpaKGWIKAu3iBcL9QckPExmB5Zo3tRw7LoiVm9RaOWoKe1my0
jGpO4zEc1PCskQZlQHBds54sPZcqSwDe6edjTYonl+WjYQNSXCVrkEnAcZdKagAQUGq2AWYiFNmn
CoiQgIb1sONxW0oEFeUwKaMrrwi007y6cYtXAG518K7wKyAUTPRWobCozA8HtWefODRFIda8At8B
HRuIJ7ex6+it1cvaWsIepQsYtCHjjavB+362OYdgxhw9mdb674L+kZ+So3D2bOl3VMMHjZCaKMva
g9JObYYnzwbxSMgYt+xK8HnUOudcH56yIcCpJYDmiOh2pQGAdfaGzlkRWXsfRJJS8JFa0w1d4VKB
Z++Q2tu8aUoRaIc8R7PsRv1nxTigy5WgkSFqunZyBC46dDlE+ivAla4yiITDExHA3Y8gxDF71zTP
mLiPyMJw2/9yHG9HaWEU+KVEsJYYI+rOxECBIsnY3LHMikMEyhudV9u/rSsxSvTDwGhoaDD4PStV
GqgVd44oq8NudkSWR8YPKocpHpzWAr4PAQnEfcGa7DFpOtsv+VKCfKXlo0/lPwc8olQLQvJZaZoI
oxl/lYNac/CgF7xuweCBRug9+hbF2IiEZJqDCTKC4MLeI7XSR3xe77WsBoBQGUw4sdm4j1B6Sfgt
CnWB/OMD1ILARb9vPpeXUgBTNG1AC25dGcvudH7lX5wbIXWqyzjCW/eHAD016/aBkhsPveyCXC/N
q6sVqwcYbywPfKIsoXrhX/T4rpp4t/k8poGfMhqC1q9wDyTf8Ewu0WLpH6TSC5G8hzDVzcQ/2z54
KAWD73TsG71n/V9/8L1s0cOgBaIm97B4Gl6TiWE+FtSq1nRrOtA3UJFb5t5cXRObeL6gm2riztmO
1To4aPdL2Mf0ikDqADymoEq+vghGOefoX91a/iZF/ND4FExYa6v0mb4SqoZjr8belaei3PXUbafm
R/9L/e0vov4vp0PAb881syg1IjOVrL5Zl4ZDF3xnUmX41e5kt0L86IooTw0+g3mfHZUyeJy2aulJ
2dQSmQj7MzkXyVDPdhtXeDeYUqVSxyxDpk/PMHNiyxZ4geOGnfpRe65uHLQxGXNP8EqaaCT/EGS3
uFEwY/yudGuGXJ+UZO+0N4f3EgHPV2sIwhJBLDVD6CTajTINAzM7XfOsCGMQ5OIgDLeE0q05fWnB
ufd6RI5TbSOPahfE+wYjl9JpQOxyJg8Axl8F+yohe38W61kqM6Mv0+iRDNSyow5pyw9ZnXRF9ifD
M89zNXZQCvAhhe1yHDMzvDdxTnaWPUZ9+MEEzF+ycis68QHd5jq3VveDh4yS5KTiOnLCUXeRdGzM
kd6ESxnRdpHWvKqVqU0PyPVVMFZE7U9w4ZUuNgAqFJQZwCxwNCCvas+kD0f4LEeHBa6deD7VWGC8
m1P3ozb3ySTgVGy84c8EV+ob/xgz+axFbNzKYCei0N6ZIOul7TY2FBWuhSAX5sby8up+UmgQbPW2
queDhMR/zjLGm4WRzhV3kT8lT67nOB0QCIXNcPW+pLig/5jHDuHcxgtPJI0Xb8qM6o/0PPjXLPvl
HE41IuYPDlOqPrW5NIqx0tSu0TuRmUEI1YKuodAu2sNvtCVo4PXW3as09TRdG+6v7ZanqgkUJh3R
ROepP2U//YafWanjOPqTZ9SDcbxx4eaeziAW7v0j7v5pmGJBbjHXw2K10IFP/n0pD35eoL6tP9zE
xlUX7sidb45SYNp0odCxPjkNdBKQ6pyZHscJXmsdyX8HFLNTs1/Tr2Sr+CvgoBDTm+rBzeQLSRsI
oR7AkcsKNfeIHUA5O/kZxd3CjTj8UD6kDcYyp+TnfRhqGNoutKPlsV5MXNRdpCvDaP5v9gYPxJBu
FqWXyzp7/H+ATgTrT0/akYmjd6NMAXXnd9/ev8/F7IEGuAHoeW7kn6LWYcWJd5chBMX6egp23arc
EsLBaCkCOeM0dJmb2NiXrKbiidVCmmaMsyQDlmRMYXweacxo3orxno4yEubZbSpYeyBy7kCL8Jy0
ovMsd7JgFig1+Om3ItuuvRtd/Dxjk8NM50BulZEB6qj8ngOJhoaNJuNFy269sg6fsi3S84v7FvPS
qW6azLftG2/ZbZpZkwaG5P6WlPGQfXLuINgvmStpPdHCGiFSNAh1tb3txiGRw+36/rZk5reQQC51
sGlkjBPWccpycayw6mTzmrxeFxnl2qwGusgLBuzSlIWEmsHI7heSTvNqrBcPuOz5hk2+qJfccWCD
hkqpX+3H1sYeZLvtzIdmsnCIQZpwxhXskHLTKICTuAkEgmFY0m+dcWJv6FtYOf0TfxZ2Js2CDCRu
3ANCtBWJRwecNesw5ImlArWcFhgzWMTi3ajbka03fMe2jxoM8AfV/4qAUSEuHL5NOJKn065OcshF
H980qBRfHm/s5j36dMjuOMHhGlgn+Gfv6qqwNl4XlmnqvclrHhP6OTI8BYgL1KnNfXaYZJ0P/h8M
22J4QBAxqdG47NaLL84z5TVoYEOeDUQLPtFRV4vTvHZzRT9aWssqDVJ1M+Vwkiy6N98p7wSZWxEA
JYTyxNcySHcY+JG0fsge6un9GndZ720B83FW3vRNSjuiiTW4pDIkuoMH9fmB6dgXwfs6C+MkJa2N
ZYlvAN7jLUJ5iz+IoyzoL4Qp0ZNuxtvpqkL6Iv1lzDJ9oN7Qj697XRcKF0YjmeyFrQks9iFzfnSQ
cr2nBzagRt2Fq2S8I0oCcdsBE3WQfTiJqGe4+LHW3/St4qO7BkOZgMi1cwXou4lSZhtTSrc2HdFd
GJcWjzqhJsQ+Q9QbnBOqSVGFCQYwNFMBcJn+KVzQT7E8gF9OUH2OnJptA3wX8gkGCDuc5Fz1OamJ
rRDwIUgy7gGZNVgv2jKFXCJushyFf6cOMxUF9R0J5JaTvZMBezacBg4PQHk1KaTzN9FfsTuydXgK
G0F9MeGAk1u3wBGQ3DTVpkSVI1vwIX9ZdEfsKWL+/oW6vJvpPeDVRHZUt0PAFQ4qKlvm+M4KbZcC
ocOvPZqdW9wvLPcJ4ELVThB6ianKfZMwLBpe9k9KB35GJTyv05GA++yrSTAGXt4Jx3bbokb9sLSF
6vEoeigOeTX/dlNVD7v7z9gEsUGrOElhvc+5EqkwxP7ZLNyeRHFpjXhBEHBmHOBzJ3SbKfHp5p6G
RjmP6tDaR8EdmvHsIA+/vd/SfAca6zIwhaTEWWlGgh+k658/kEMMKvynLzEBmwzbNA4A8CoPDvMU
LeTvY1VqRsKnVijwQv4Eq+pndclDSxl6vHu3RKas+tR2rEVL8NBfWrnVlvfBLbmxpM5VC7xw19QN
o7L+/Ik0sWGOnaqF67aQdrCtBz0J/HqITwFYNy83pnqx71aRzPWS3sTMsjlLPJJ+5fM6JTC1iu3M
zn7SCqQrtMkGbnbj1hJF1ZfhfUVTDO3M1q5YDYinZG0r4K34O+WxN5SR+CVrFk06SPid3EcdjsLq
d9fpylAq/gN9nMUDzL0GClxgjXrIObX6mWnIDquS8qKZi2WYsVf3wOMWpxpWx0dKV+P8hrda12P1
6LDNyNG5kGAF+whBlvmDbsMC5lRsAyu0OXwIaRdSm36FelTDK23BOO6/CbyPhs5Cim4dT8n2hTEA
wMqhTM7X6yHvgYP9Yh6H0lecsw1uXnCATTV9ATYQyeHc/0SqwuiA/SiB1V1HdF04o5kZRsN6lr8/
SOCyoJijayOTAhf7qaBBuMpLFCXqzc8QPhsgv2cLxkYmSyDn5YnQCg7fbya5eyeGjt9BiLnG3RG3
MbseZYGDaU2kz8gDA2HqJsdBRcfNNDglHNmeQeeit4AzeUeCrL7k/CIk2EFD0dc2Rjs41lmSPqWr
0S8/OdNrLj3b9t2gDo5MbCDztw5fiAoEwrNqib7F/JdgHwHk3A1zEUOgK4n1y9/05H23XzBiEuN4
svZ+eEXuc6y4vfLo8OblwqgCif6BxBZYOKLceUDMWK1xiDF8g0+Yxk26kjkyXB0YUmV85owaDmiA
xN1hRJ5bl9bwkBErSsrBoiBDLf/8J6siuFiDZZ9paVVs0Zytpi0aa5rDMcNHGZGZAJTbgH2Vz/QF
qLPgaRCcz9vs1gPZsner+HedMlLT18T3/sEHxEMXQ22tT7WsbfJm7ki3Dp1D3DZ6PLuYTuCunDjE
Ywo3CBNdV9TdotQQIBiivpsc90pz95QW50zX94LIATATRbBKk75f8yYZNN4auIzEQS0xf9GmmXQ8
mzbX11N/Xg3qX5hI/a2E/4lZUu7kzi2oNJJ74ipJB/aRK4ch2WUkA3jRvbiURtI4SNZxtHH4zybr
d/BM79xBHqfmwQyMIgVgwF1p9FBgVechR+sXFhGS6MhmGmfr6vldsWFkQou1EmUlg+hD6wOuGxno
TRmcAeoSe9ou37NyfSByMiSvBdqbUUxszbjFYZE4Y6bhwv1nGOySiFq8YoZUMMg4tgLT0K+w9KIa
LfzflTCeJGex3lZP4L7QEhCB/7x12bQ2N72+xSvTxGNRz+nCsDiyKnhfmQAq2xW8hlr2MZEq4Gx5
NLcKHKJxUFSWjPJl4y/LaDyKeMOzTujWSqHUO32CJH8YPjK28M+prGBmUvw4zqgwS6cf8tyMNSUJ
hm2dYu/lc3rEOBNNKrbxk/omAPtPFLij6g81yguQmiyUOQM8HhGrIwO0I6hVvQpxeIiAkg8l0ghl
NFQo/WNTBbhRpozz6O4YR/tPmUDAyOREyaQOqUy6wwJORR5iJOC1e6qT7HJ7WNgTZYR1DN65UX1/
jDj9z7fM2xhjhwmQH4La7AKuyEhNDnPAQUAkWHoGa+BdlYvLQ8zbF/HaskjKmPGDq7QFnKtK2chF
laVFvaKJh8hzjRSSJqD7gXz4oy2jhmvCN17Us3lOvu00d36GFBSFB+uZGya7yBuJha09WYXe66Gx
una5xu7mgkUW9H2YdvHSq9npEeOxa72HvbrT+IrSphICnuP6cWEfZ2cSOYZb1S8uoYsDFX69iaAT
zZvUOVmiRIAEdKYsF8kZ1+iD2+TktRruEtxRhT9/SyGbfCNbO78MMRfiSEXZod4DpMBBx+E0PqN+
Hj4q10BtIWSa9cuHjr13Xjo+6vmUFPBOixi2JhY9btRRT9RH7jdWFSu11FIyONHwmVCHjYsGGpgn
BHfgav4itWHn9fG25Y1Am0FBwW3VXb2Pa4x7J2ydeCpzM9uZOEedI2CA+vo5I55VeiCRe4yna2CF
49KBcwO6hSyj9K5cFFmooBZeTRxGTB+UlTjQTgTY6vWWay550QhErW++J7/CV1uOcbEHuN/q9+3u
TDQNWL0nsuqmwN1D4aJX87XhgHMXq1ca2yIb450AGV6Ziukt33MxaH7zTVlgKGVZJ5cXPcAWwMcv
sK6yQZuo6XGu4Yi/ZqXCK7ax+72qva4PbRQpeO2bhrueUcjNDvwSXk1S9WSNS6Nf7ihDlk9Djtmo
VEJzHKTgndtc4mpjaXIHKYx2giA0beYvu4AfXjUSLnyKAjMySFdtj6URvrF40Hnd077VLUJ8r+/w
XcZYo40SCOAZqkIB2pK4jUuTwJwNqBk1NMOf9lncd6cAYJIK0mOcmjL0fl/VNhHgExN9MJHXzzNB
LqPzQwMk1TGjA4+OPgPgRONYuL+onEU/7AQBP2qsxr8X2PuSyUBOyD8FIqySNVOEX6H7//xkKJX9
1uOSXPcfshHKkYcBn//FWS/JarQFahvFoD5H+nOUNF3VdQtALdEdw9O6KH5If6udtmsVzIQt1zte
fTBijqQyXGumAeD9aFSAHtXIAB1CdimNX2h2YSjQonHhFjpPKlP0v8mQk/mDiuwmU8Hwch7b5h/P
EC/sqvcoDvzyFTBRbS3iE6fyto1e5w1tDkk4Umo7RqlHwh3ilOp0dmdbqvNy3sJbmnkT2vAuLUFf
VcOb1aLQaFdZBaAPys+YeAS6ENGnBntSoo/qqjMvaBGj6lEivzGzSL+ArmbdRhQIeqFClBpqkSNW
BNGQCDsZQLsUi3yzvewqf0bNg7ZpfP7FPHTus75skWFX9R7GRxBTohN3lA7+4v3D34xMViMx0ejq
N6Nh35BnvSGYPktv6Hhtr2OmygRVjImzeUm55rovJdzD3V6nSBN7cQ2fXIJvIYRVkmdvcLkUbOGA
f4/NYmIIFTLpGBBBOnbqRs1eMCEZf4rk7nqRya2Wobp5oms8tnD0elE85lefNaTIGjrOZx/H2C/W
AT4yoVdBWXe6oR3gTsXrq/SjC8t4f7BTYUg/ngGDDfCh17Dlc07+Xr77oS6uo6OiN+4S3FMxEFxF
33d/4B00blHD3vYhD/Pt5BLsJudA75qLq111P2mk8nprvO/YFIX+UPr07mej+Wr7wr4dXN0b2DJ4
J5zD4Cu7TLMm+aVTJbWQG5muC4UM1/geUzRjLZjSteLEe8dimXsOUtSF3gymDZTJZlcOeVqpn4J8
lYSV2j8L5EePbv2d+JaDHduPNEHdApFeqocM0bI/fGmXggYUG99DOGywl+DT2B3VK64XtO5f2Q7z
gqHvLjuk2/58GTLrVxuthhBmUQDdrJaNm5DsLRcWVL8gN7/f8AuPCxtmnNn0mIwEHogW4LquFqTF
wGmB451gvt+ow8ACU7GjWmDGnwmpEtGtu3SUJTYA5e/y/eq02ItwLVU7r6efUJoqX7Lxh/2FoLQ9
P9UOjEV1W4Uu473Ur5UQcJTIfxT+CX5NK/4h0sWEj71nMg6rqas9ffsho7a5TYq2Mg47joL9cLla
rhYK3VQ8yiezE3QE886iVto5Fpvw0FjwQANnIMEbzdpgdlSQ5kV2TG4CDarHWffHsxYFQRg2QHmp
bUifJ8SPoHXP6uF5VmMizMe5HVXj6X1Vw5lXIq6CwvIzhydcRJWAMUnG4tLjzhL3y4eNjQmx+5F2
WXBM6gyJOkJkkNY3PBOMBFLkWTbz7ftmrkOlSAlc/szfANxBeYFmtHgKsmR/eAujKSfAndmalwfj
TTSIagicFo0oAMWPQCAADIaMhvz5kR1aCdKlTnBcO0CN8dOmR2rHCDJJBWetgNH6MLk0yS/Njpj1
jrd4ESQBvu+oguq1GGIevsc1KHqr3QlvkNOrnIwgBmt5PZ607rOZOF8He6AyzZJ9b/4u/hUqt/xW
I37Jd0jZ6tvJG6/T8w4gbdPV6RmMcBCCulL6vMS1/zEXxe/NtlIGMlMADTTmm6ZoH+dlzD3fEcNs
c2bxDzHbSo4EsLIzG7na4bHdUOz+zDasfUVJNEHrUH13OjwAFR8DktEq8bpuZCZiKjggEMiqRHr7
TgfT3UQPOtSA/58mM3q58UJyB9xGr+FJ9uOP4I0qcLREuElpkiG3jl0EYEZm9XTZkycqvQzLQZhy
OrGWjvtttBc+d8rygyt6yo70xD2rQe4vw4I+IYE4LZoUv+yeDbyyLDt1qiHUs/P4GOcDAsl7Hsaa
LLEL7phIL1sQvXMyRe7hHHo5nBfrpF81YFp3PPgViYiPmXY0Gq/69uXPGVsX/JlsYiEgbA3/Z8VJ
C3do/pML5enINJOaLU6Cuyl5jfu1ekG+2kK0hhiRj7CaAEphUDSx2/JmGEOCPGxacYtX05nmm4JN
E9eV/QHJu/Ja3Xz/yCrHbAwcV9viPXy8Z05gVhbBMnr6o9KBPOD0X6f9dd7P4OMHdWgX9T0+eSed
5vyKulNyCphrkovEEEdFnv/tZWE0nYNjb7K/SRwU+JH1f/rIfUJMZfLQxu0V1V/muDjJUjRMYZVR
q2SGNHTigO8+bY9iwUulghWW8alEOCiqkc3es5nJbvYr6b/1Fggez4Scug05K9B/STvO12JgZ7Ua
+DZPjC2vvL9b9ZJzghJSN7rLlsitRKRcwXjPK6aQMKQPw6BSz714mw8KDOJmx6oQ4/qCTZvawoTC
I7n5IpumtzPV7HKt9GfJ85Hvb0FqgYaeakomkHRH88scXWZL8m1u9iDSj3A4bhw0wAZvEDUce4+n
w8YwsPedttBdW9tSmhevzh2y3Oq+YPGNeDVHM6mCpIhKX+oMS3FWqIo5ynGRbkaMsnP1wDQL2EK9
5I3fYz/73Z9ByrdAmR27n5srOIMCPWLv0kWCwFuwOz5bwubhLfzboLGfTYzEU1vfqjtKjJDzJiIo
GstguTpB1q1tMKSg6M99ikQYmFgSXgPGuhs2HNCt4Epe9Vi4HQrFLmDmbxVv9ZL8iCUMmR4CJ8Fc
fttw+iO77PAYy8Mi/yRMLcZ+Q/MR6Ol3Z8jsetoGxhu52TY38AxUoimRXiAKhmx4JcDXRw/wjFui
wvV7I+YMFMzoRLgUW/duOGVUxw+suwbTf1pVtg877679kYYLf9+fzMJt+1wnkdkd/YBsY2jpjml2
xfC9hCk0K40/TTK68BuF0guLAsx80HUDsZ2WqmGzUJ3ZPxu0H0EzaUEtxHuM4s/+QINEy/zObidU
pJ/cVVIrRSVMjbzRH46vMKu4oQFVLsgURKyKLqe4e41wSpD2mkwmadwXa1IJyJQiTIi8jJ5Did35
/XlnfWZeKtn2BBOUyoZcm/lLabrQeGW/66HIRaptBuv9iviZn2ytCtRXzPSikrsjfzzgUAwRBRSw
Kh0Mh8oit74r5qDyq4BqYQv1ok4t5/tJ1h38H1hQ3Q7d/7QnbGO2IyZ7ErTSJRdlELsftMOx8CEM
F0fXTeRbO+QT/bzczHvmQCMTYKjn833otstJIJjaLNUgHjIExEqblzeTa/da0pEXB59gncxYEt39
X+Y9AbErTwddI+z0zL5sdRAU5U2GH4R2huAT0X8g3s45iVyZfCx05aeAwDIPVqVcuLnIiu6gXVyZ
cRnxnDqnMKQ26f6mE7V23amhgvigYIJBsIeeow5zXqIGWYlZseWxIytptHtsaUkpg/oRSzm40tC1
tpXzE+DKdohc+eGBaevIEfD6X6Lfm4ArloT5JOsAanhZX+1tCse60VlYi07kUstzL35Ek297wo23
fS2pbroVN0hqV+R3fXMLCk6WHd9fw7RJbbl8KFsFZr+xAM+aFXpf8nMHuMH4YPK5dtmgvXZeoGwz
SUbJX8/dBDd4R9D9pgNAnPwjgdrrKxLsppcEU4BS76DgIdknDDD9rj9rqyciitJfaQ3I0nTLdE+G
GahI+nULWlAvDMiIG/1axaQNIFH5Av4mzjzfUWHBw6h3RIjFGwAyX8QDwl95BztSX1j5pa0wcO71
W22Cm0zJx5ExSCLQsQ9G2EveNBUUZxeCLn11js4I/6f7I8FEyQnepQPXHDkC6XsFneMD0ztbUZQ1
a7Yg4lyGk3Tgo9GNqmz6xm++eRD8Dd3Fu4suhh6P/Z8lwbp5L191+TYAHv39VUlUIjZxEbzdsYws
N4TmrbY60Sl020kLBjD0eTs/liZVlWQmzKLq0BdXBPPChIg360rNV0GXU6sOzQBzZJNSkkkEnk2M
u7RcJ/gGubDswROMMdlW+xhPZ3+igUVc//CDWIY0W5DKXTVC/lSRBAesGCfLWhEmDn/YaSr7wkjd
LY66/NrIGMnCR3BsYbpIkttEz9upXeTOqfsovVL4739ux1ZdND8AbMp1t6Ofc9b0DzGg8o9OFsls
hwGH1arjSUxBMJDX9cBI4XK87QAUDaMRK4ZWiISFvwDxuUNn+cXVy9gQD4tdNwxIrnMl/Cby2UDx
IbYsJnDx6Ae0TNOPYXtwcKJeTHGlBgxqLGfr2hJSSSgCYIV/N/Ep2u/9y+4zENGvygJi4jIHw91r
Lsv+20jDZba2N1Pc15LYJCJspdcHmWsQFNZt/6JS1MxYK7ycfAMEULCRBLdIjr0w+Ttnam4LaPS2
sUymR7QV934envAll6h+Fwvc/W/jkS6XHNmAd+ADAWZ6qp7p7bXeYEjsth35Zi7LARnu1MasbIGS
M3cNW4lXt2d1IgohLtredl0GBBZZA1HuyRPVgTuI7Q5JmyWu45NRCWys/lHWflMu0Z+cYDe+hdDu
Jigf5e8SQCASXG1zQLpgMtX2v1cMOMj97w7AymuXh86YGQL1noOyABpJNGxz78Vmqd++MHurS5GB
nthy02Znyu+SdNadmz82oHpdCB0UaAHQy26sv7gBoHJMSKcD1+CrB1cuUktVGwBdFGYSqjWRi+71
iZL/KT5yQhzW0YahFZulWyECKLdCH+8CcOxKQ6fzIg88q1bn3W518P9D0OkOYoaQJd3LMIzHd3ck
2jb4hvYRyE80cPbUlzjf1mTRx6ELJ8w7Oq8p66htz2U/dkJn6Ud1wtRO3ZXmxZGfxvt6bYBkJ8Wf
/6w4LINXh96ickHtrSb30gFWnRujXNkDLidYXIGXvZXu/rtteFnQ1L4YDvtNoSp0uokfiPZ+4mLn
SnCdbWsm2D/JqxU6UoZkinFh1n6e0CoGlmVz3CuR6tLIAN1B//1KNfZGORlAf2PUsN3lLML1DOd6
BqzSeMvfUrT1R5HWWuWDRf+HiLkSwW0EUYR5G17092T9WBTHhVWdwW2GYO5wmyOKd/1dmAGPRZyL
Eh8ORnGLDt14ywLPswzDJKp6B72Z4pZQ64Z9L0Eje3OwnuIzYSq4VvrzoyqGyTildsUj+HlJWcXm
wfxPgOPQoMSu3ESZUpvUMToMxn6Y/JoKtLyqzrECLxOhrjXuuOLD6FhmrmVkF4cdwwK6+xKdCBZj
WlL0hB9+3zR2nK9SDXPDca7TkXXHu8uthyDsxMRkekcY7tCJWeEFKUfktf7nEheK47690Vba6NoB
sOSopPdICxDGnRH97SakPQwGTauK+a1UJMBzRK+F444IS19s/dMUycw6Lf/tdKL9DzfCIiwth/wF
y60G3MIQ865AWXFSM7PtUwk4fuWzgHa/9WhOG5HpDoEbM3jABeqNany4klygkeKuesXog66WjMJv
65whuohID0298ECAoLZPARB3xReeUYqCt17htyB4ZLCT1TuRVhsy9R73ACr6/r+J/qWs/AyWz9AC
2QE8UyVaI8I+t3vz8sG1vB+zNtfhN0MSBdQ3WyS9zb7QpCOpLG3kDRwqqeKxUu2ksB9iqrJ/O2/b
9HC2go8HZlCAUS4k4VJohQBiMfNNqgcEtCuonBSjnkQfhaJfrLHPPld0okgggHOTWhMl/EVId6aS
4s1Fd2g3hn1sh1M8fo15rLfJlETuLmZR1v69dYQWJkwUq9V51foQVYgLTtIkjXBaY95/4ia/wJvR
7j2aTiq3W65YSmWzdLXh0M1UViMkjYx/mYkbPZeIa/9hizL4Al/FKBi1F+bMHwMg8XQ69acbr0Ma
kAC3QYVVEt854+ZthQQ2PxwLa1546+UnLIGsr0B3sMK+H3BXl7ZhLbPOW05vF4S/L9NYUD8qjXeN
B3qd7ytJrWTRbsv6rqprgZHNdTaPG4BulWgDjrt7CRdvEud693NxXr3DjZ4t7B+S6AiEXXaHda1H
WXDlxEf3W7zpHHEXifVIFfw7fdQg00hBVhif06ezF0qKdX+nla4tNuMZcL2pz42uTd+8ZmV98oQG
ZXX6pBVHzfpf/47Sn+5i0FOWGp+0w4/qgmWggD6SFt8HYiULaOHqr5Dff7nsGCMud95fBz23EioN
ev1ywndiKQ8JbhObCbz0GLkEWBN3IVNklFtueD8KvWexnLCuo67HUIScwQrxYU8gwWfknXI7C5xL
/NnHdLbPjfN30tEzsv0DoZWRGIQtoWBUxs+htEX6XPzYek+2ig81qy6KfXsa/E5zWRQl6t+whB6F
jIGBMOwiokRS6nUTeANxDR9cl1xC8fzd2/0ci5XknQy2U6xDPzZuc6IDnSo5SnZL7tICijyN5R1V
RtT7wc5V94BvCiXcnrzAm6niEbF10VYknYm5ymm7FXnLWc14FWKwsEMeZcr3zFELS1eNYa0Dz+9F
gaV2fA9KIOVtGlULjimgeRzy0E/oDTTiBMYWYLxYj4EEkC4pEiJ3YZjogRexwgCQ4EHX+afr+8i3
Yrhha4OGArBGYwniz+a6jvWYQ5viL1KF5UaNLxKfFz30WofAjKm1GIbrnaFb7wf5teXAzBNy3RtX
N7Md2PHrx7z4myOnEf2xfHHjyZA5/DhPAgoj7PqwGUM5MBMZe/NS4m3FsOKNokJf21Q0COT6isxv
Fbdb0rQ+dwduC+CMaQRlG6v34YAH8mScrMET1mNP9eNKWIonwUQX4AHkAbAP7xYhb306AOhX5VsY
GotYZ7VtpUJ7CUs9nrw3tjOLlN4Iv1Hfx70jHr/weUmnfcPgv//oi4JO0M/6XOleYqfkUSXFpl++
/hWv6vo4Ah4iCvvH3cyy4r1glIEQKok227MbhEJ2REVcKDUFcnnTPVw/bLGp/C9vobUS/p54ISgz
DBRNt1I6ta1bpb3EScJIYhWQ0spKjaITyn+Dvtnc6Hr86KJqlm6S3iF6fF7TeXbar8rSiCJHeNYU
E1nT8pMG3vJdc2oSryIpalv5lpc0tU0C3C8GPqGBkcUMeyk0ZeDqWZCifjKKGRsEOxPHzT0F5omO
WUtt2tsWGBu0nl2NaY5D6vZCcOr0PcEwY6cfPF0qFvlM7iGQBh1s12tW4UgXoyV03nweoCUbSaul
/NBnqMil//Rw7ebigWDcOtzEbpd4la2YGx1MvZvB7BNQGjsP7/AJF7pP7c1hu7kn/ilSLpUKN0/z
JFS1r1XSsI8DOgytirsMR4UV4f9RN6eZ3LqnORLCgbdUoQj08PyFC4XNCZ58f3ad+dQUFALa4Jrf
BH7tVOGDlKN2gdIBdNCGeDZknvz23mwKq+ijgZobO3kx88K6X1aLE8iKZM2Sy0o75AMl9rs/8wA+
Zkb3utVvDdCTsrIVp7pOJkU0V34wyi0Asw3iL6hl768zb4b+JPF/MFh1cTzzpqflwU+vf9qSsjjT
Rx9PgmMaaJHKhIqIYfdTEGM/rHVGsQ0UUWGfJ0Dqx9qiovvJcxg14typju1bD1PALdAsvzjfrTqH
HDs5rEgLpI0jrcNmHahilbGIy7vjAOOVdlePot0LeYlQhqLgoETCWPZeBEPWjIQXwmC+tFpJuRMD
xHOsI/0cRMvChQc9cyREVOMTqTcLE8szmqpNTxNZYuNu0BNamOSiJm6ZNNHQAVa2cC00AKPpYXvC
bP7+dG3DO6JgD1yhvB0UXe2qf2zE467VI30Fp9TAzE+g+wm3wWn0MD5NIFg0r9bVYeBAeRzTON8L
QgWXdWCaGb/vv2LnTvq40U8y80fI1nLNm4TpQ108JhYQRNHenJo46YbmKxeOio8F6wT+qqWRPf4t
jquzOC4h3FlzVNHgzNDxonXC7lztiOsGzHVHDf9LQNoaUp/9kezllTLHC216e1pmtZuZvC2EuTRM
U5QW+i0O2D86dbqU2ESIMLL3Ae2P2XTq48MQCzgMlJqWibxdNMoNZpcv+X/F2EFWnrh6GKKsaobJ
potaY7/9wIBhB1m+P569WwjfcjG+PLoI5QnDzKz8oij1L0Zb6gwgXHfKdZVULTmP5FtQK5vihQ3u
k0Dmq2sykt5DeqQQD/Jq7Yyus5r2fa3RHjBJLa+NjSP5TElkG9NpmgGE3fg+5OsjmFWaM6jFRtCb
DGnPRWC1Fc+ctYxCkSiWfGNled4Rkwcev815VmOB23T8zZPwYbSYkZi1cnchVGfYpVRSqxCCyVjW
GMmxW64O+P4hR7JXDfzDA0W38sr65cSXhxaj1BFtlAyQIoROZjOM3u0lx6xkqS4LGcZpLbibMjyH
6mKeUy7zbcnTU4F6kLBMaiH81lOJpy0yc/giLBIc/DyxPQ9Vgu7r58m0VFrEx65hVYooId0q7nem
cVeEi+9bOCh5fh7ZUNvLqeSzq35DPNJA1K4lhsoGnGpn777SZM6gVq8VTkdDROQUuzeXkex9Y85S
MiRIOfy51oP8Kbc1xY3ge311gaxart39DDE8u/4/eTlllfI59tIQuuWt6lFLbvMeQnuTLVXjAGxY
QdB5IqrzsKkW42tXZQoRjEU3Ml6ZHMKFVl1evpkZm/7VQhpR31aVMEqarE78Qa2LwPfTlloOKSSy
IX/E+inRcmpoCkRBGF8AERBa7Gq8NDKX4D9CA81Mro7oWLT7tgs1P80YFEdXhMquKFCEiEIbleuy
2euUmwaiLAqoAu2BSkILXObKddAE/ZN3CrHu1PN51QEKCg08kq/Ns7zz6rJ+HkqN4Re60TX5k5VM
Bz+TdcPD7r4XrlYTRD+LD5DZGpjK2RjhEl8s/4mLY13q31sHoQn+tHcEsZWC/brnG8rQMCMVsQdi
beWA0NWeXaEP8+hNc7fyWPUrBaQJFddyS8On1UhnCDkrRYSPisXHGoEctt6/Z9sKRFZikHMi4wd0
vRQKwatoSwiZ0D5HOJ+grQ9UfzZaLA8Nijojo7Vtxxg0qcHIfoetFPiFyLb0i23blkvpbc0IRVQ1
Cii90iDYYsmbd9TCrDNfs3B9Ai5KuusPd7arttVX3sgq2YWyFIw8TaRGxvWX+yWL0gN8aeTBZn4H
CgAfKkUJsQGwoGa15xkpPgLKTE6tiWtsFD2ro2QDxqmQhiBtD6qG7dIbMeRIKvfpRBUTA6pIYp5i
Bh9xGtelN3G7ko5IBiBHJl+ruV7xVo/22pyvFDKkbxSSSs/o427i+6FUXOoCSJ+FT9q9p4btOJKV
xp+LD4w9YT66c9FpLLjXPMGrdzHmSJKWHak+yUI+XMVnaEbiX5/0tvvl4uD1vWDXjK2oeyJXVUFO
INuLc9OT/bgfHeHQ9E4cqStuQ9Yl4rV5bN+A6E9Ta00Ef1LvNoIIRc9fGhWui67ED8VsRXQ0+IJy
UYlvtU+pETJNvS5Welk0ltLfFUIryi7YhJHzzO9OHeR2IEhmAKHMxl/N59ef5vjuvwXwxU7IVDOu
777rpL5ERoC7xS2GsuFTWTLBrP5yKJIAA9ore5Ppf1w0mkk7irEJUP4Eb9vle942anX3EpcREnZu
5swp2cTNGtFXcwCjZQLVpVM8hXRoBvU+3pdx/+2zQJjItAtG6TRkkwHCz0Xf/NskoAhrgjmrVZD9
lb4nrUtC4Xm6vTTMDOZNFXS36vIb/L3J/pWV6GB+UgRrKQJ6gmFjEPwU9B0aSJhvSUzAvzf954kA
SGbSuzNZxJpwAWfc4agiXLNT8dy/kQFJc7gTR9wlQ7KlJVeSxYNzk94lhSJjuihXntGucM7jVAWm
XkNLDFLyKNkgZFilDtu2aHjjVPPHTAGpi9NuWy+B7W16EpnR5YyE79+8pSNxzDkdR6eFSThlpmRL
dlwGEV0xJSo5DbrOUqH42re2eqjVwCaWt3QVeKtsOAfr/OII0sDw41qT7W+VywQ0I8VDzbXinMLi
Me2moaaoI5qz2ic33Yh/xgl3ezOmlRo96aYM4eXba8NrRSSerAptmQLM7udA5zgkivab1r7t+A4l
1AS7vq2QBdnY2H3MnleGLw5wgn2uyjyoswzqGOYtNelBNSYkbvbOHGj0uJFaoyF0q9BRVAkKJ28W
9siOcixQpaLm9XjoKKA9A0+/QEEsCLw9tOZqESlgWe2/rNDPo3298PcSICnKV1lmMkwZeu6XBZQA
krBaw7iItIkc12PRXSTAeJX+ezXwwLQmOCV7q1/0Qi7bImhIEvy+gk1Xe4PCRJortibed89Q5IOa
/RSbCYE8StUpgpMXSvidApYhRFGSwIoclbvbNSCfzkn6jh98azQo17RPbSFsK9ogV+TE2FZkusAM
AkYKc+TptHGPWzSkNbqiwdBQhQwgkwg++QpQWojgnWi/bQOHFikxZdNZ3IhxYJ24+vVXWgi/VNrL
uP7qlp/66VBEk+ATFbpC1ibrV6Fq+H/XhoICIBzgnI46vtFKpqnYYZteme6QqYaEJlREzeRuyHEI
yOJcdzmGB+xUZ2KaoIfgp+M/dp/DNiGulR/j+a7e6vV48Aq/mx0zZGZ9X5PFW1FdYUlJA7rL3c3Y
wXAJmodSStZRjQ+qpv/C9OOpKrGbNdyKN+gu4Sc1esgXKrVdKvvIIz3PbhmhIEXqa77+N+ohABIS
pIYS/Hs9HkIPcPw/GzedxEWIWw5hCGhWENFTGDm+NC1zqcPg1AxaSS1KltcQKoXrzH2ZZNyLxmAE
uag7XLbETl4zU/oiz+yQJxKa6ceMOa2rdxxpjNnbbU1sEEtYOAoFPKb2jPX57n4UJTMwcma7c8CG
/lKMsRADiUN9PhP176BZQX4uc1bcSS5JNaU09tWqrlDMMA2glLqvu2nBZs9m9o9ssDq/7/k3jM+H
Z8DITwtnJFlDPmdP9NVosibzwqaBADCatLvd2yr7FcoY1FV7R8Mm6y7VWaexEXZsvk+jehcSN/Mn
WAspF/1eb217nfZFh+d70t//g2wIJzRwAhmWjN5NwkKkfY+58psGmbPd3SRWTFIf6Cmh1KI1gVtA
RY88BQCsfU4cf+Q6JU2fhbYTcFO+B9KuXMxefQX8DjuFy1xFlcePMnSADWvXRNdQGI2ZmmBbUoQn
VPHukEn4fQP9j2/+BE8IBkgPnqso53jkDRvEqKEaYwOxTdouuTgAq7zwAPswgkpb4tlHe9LqhLzu
8th+NBbA6R37LZSBa7gbTQ4r52DK5hEswXrGEWerpoOdpYyJhqJQvJKtsdTGDVxmOuSYBfkgWoiw
32pdLMaycnU1mxbCN0EasPzkAROmMcwKdlW+5h1V70Bt1jN8+yfkNHdG291kVHrLrNy/wVkZ3D3s
6rN6s45xwDUQJa4T8cKHvl9Ei/T1uUrXtL87FkJ3x2aJlrx0QUHFlvGctFlg1wIiD6k+Zf6P6iMb
tp43UETd2fyMEeWXgIOGMQ5JBZ0FS6BUCFN2+EBUgJtFCqRF5+D7h+wNordKJ1SGzdla2hn+5ATn
AF9wPsUTQBAwCVioZNLfWG1zoHk79r8Rx/DTUBdBuwJkE57OaZff7IeZ9V9YEFK8Psq+rI+N/m0x
JMXk4YSXyg8qTseFMHkRZPnzpg+9Gpq+sLIaNgUjeW8iBHLkRtKGg5whbeGgAFxESy+kvqPnRPkA
+0C/d8sZ8/PbbDTNCRD0mis614su32o6TsqhAGuelLYDCm1DykeZuChiGI34BHl5CQW45++nsgdV
J+qCcAm9wbFXPoxFQvOp6Ih7Mbm6hR+RvpSEyTlt7dDulmsYe9LmpdjGOAB+IBxT9L7LYZh/8Lne
0Vwmi50Iw0bMaW1yWQtztD+I3q57fGGjP7YGWBDlFOVmZkuuKOWyBEi1p6mnSOg6yodI/5PCi+3K
k87EzCUdchz4WKOpftnrF2YIpPbsLEExrnXe4KrFyUhpOm4Vxjlo+b6fbWEaKB4dmHP7buSXz5Gw
zRTG0nURiPSS+kIMITkNXkF0Vzg5YmLfk+aYoitFx0EkHEnkdJaIpVNZbCxIvwzM1S3zfOuTopYg
52xlt+JwnczsCptjD2gr9fAkLOklkaWXFjV90l/0CGFrf9k9sC2Qekwwc2KeH6szD047FKyVLyVD
hy2qTFrJO4vhe7f2AK1VFdMUYi27VUcEZbPnSVHrV/JP8Y9XGRwyVAtibDN3udE7NRHyC2tpyr+Q
1BG2Wa5I4FQzsRFZs+bOe2tEDSx6yqkzXU7MVH2s9TE/LWUQLjykZlOXwvNjLUhEUBZgq6Z09pJd
dc4EZvvjmiVXjVM88EDTiL0i3SUIICe+QIXJ4mY6eDV0Q/H3KBZYgnCyxJc17a62Eq6gpLZCt/Kr
oq4xGGFQ45dun2x9a1p+KxpdEXC1B71sER9xTscEeiuMHZ6KQ1QWx+pi/YdcB8aG/uB7dsquOITZ
IeSB6OU9qim7UkmZhc3Kz3wNog9raRulurLqjERhUv5QYssM2C/Uad1a9LEfE9lHQAePMmRch8Un
98kO7QqPnJh9myvXaoPEWtBmAfcuh1dn5PBnPpp9CaqiAonqD8JpaVU8KySrpQPACImzok/N2+Dd
I/dyfdvmFJo4n08PlIfmGNvO1Pmrmfd7lQ3Nbay7kZMmym2ihgomj06WNWmOd9L/DNqlUWeLbKKf
EZ5QL150IuoE3EznZj4ygDKdiwAqbIVhWcRZZfoczrPWQbpQl6lenGBjLeO9cHYRyqyIut123zBw
h47Wf/cj8kEdD9O4AvUcKFywH6U8qT2R+FWJKvVlkN5oQHwWZOh4+xzycbRS1IFv4rAt1pPt9Dhi
FEWJfyUnNNhzzQTFi16qqd/SxeVgsR6QK50hXiDVTFUJ5RIfnvoc77AqRiZOrfum1Bcn6Ig2Ir2S
bAxnPYuDFE1xaBG+BG/7LjsNlmpSM8gyr+k5Ym0HrmVmgMa9I+ce3iPK/KkQEXIu3ZjXjFQcA/9W
g0tjh3ZKP8QNWlYHz1TqGw94Esukkamyt4i3qIZ07k1v4XZgUYP7duym8OVD8TSAmknRhEzTh2P6
JPRTlN5tE7RVhEy04XW8nVNm0ldIm6GONS1YkIX1QiPMW5JgXVj1zJW0FeXYBkFlozSkt/5NvI7w
5cpvQcH7ZWDocTSbGB2TUPHBVjH37ew5OkyQQ4ba1yySy3mMhvDHbHYO6WXZMmaWX2+R/ZjlG9xi
r0bahzHh12Mh1FKdYNA8+7z3nkYcJYDhBqEHaPwVJQcLJOi7OhWEFsvqN/gNiOEgPXhPXTtaqBFh
97vrfx7LLwzTL8i7vQnwf0KQDKkQ+mjzMTgR7ADR+84d3l0BBR178eg01l2bnQMO5m8spdeNZR7m
LGpDgWIeRaKdEht78jxKzyK2vsuyDf3md/bfgCi9hX6n0Hai2446/cuaWbBsMjCEZbtTwd/b3YS0
p0kJoYAJEkv6w08gFLrdPvEqalbB7MnMoo/qCK+jN8e1NubwJmLw6RyTy4DUbsm2+D4aasNTkCbx
zvdKnbuj24dRMoZhNXCi85lX7bqbTusCrKvBiT6JYglgRReKeeXbrKjVXXDGZCv+1HMLSTqam00a
5BxFkWWoP1Y+FV6AWxEt7A6cUqml5CrY3l+y9DwcpPKYlDrwexRLK3SAxQXU0by8sa19xQUhuocO
5GYXM5lY+e7vQPJoeDpD8hJ7XFeifuukVsWxCuIfVzdnDDKWroFzZJufLrzsTRIbQEbfL06NIenY
uryOkSUKUJZCrvX9Ajg2CvyybgAnMMrsgur0NM1xL566J/8uGElZb4cqBLDTSQ3kcqwMr5Up1ham
d0l1u8HHopdFT3A7+3L1x7Vh8wOEKLczcN5+6aeJt2EtBpYxipRP2Zzt3yFQJ9b3ze2myRZR3yYd
9/gQL7i4vRDXkXqVBse3md/CtjoU08Psv8OQnIU8QR05SVMxyRP6wluyQ/I3YXuOM5NSGowQdZj9
kqycpvp+JuuUEuTzSpY1GloJndbxMXoJMzp/6nWUIPJFdXfMgmhJibo9lLtUXB9w95oeEyh1+8SK
UbFq4dPzVfxDFMYLdCisb2eKUJtAoqajVVt9Rq8/2VIdiv9Ld8+L2n7XDmG5ekw7kWItpJ2PSkM5
ihyMnMqu377pyF2ed8w3vPSCgrY+UI8tYE0fToU4iS/9RetGRMmFndN8UjwXlTGSke2FxLa1Lw/a
5MibhBxKaKExxMF5qiUQEF59LPKKGUuqu+o4S6ESSj+RsL1ymJf015+zMazdMwVz/9ybQAaVj1I3
1OaWqNNulFu+5wz17ZCa4nCVmm/9ehOqpu4ruHdsVn2ebG98XSZe09n/buK9eIxyAk+YAPLpLRqs
TO+g/2TBjS8crJA8Deb6KLMNPNiwNfEHXlYJKSxUMgwWSnSqYDWqnnnwXU71qH8s7+BRMUTIyKd5
bcmH5zaJbS23cdcwA9H8JZJU8pcPrxG2S081oeBRvbRH+rEIzwnBBIKXbxDC4s/gRv8Z1HnBMSiS
nONbvwELd55VCe25VcFOUO7OVeXK/VcQQe8jqHZskJFOuQBl0wMYBaFAOluv8EirZfPn3NcIBlyF
sI94eOjF7oBuK/h/QWLAzzrZKqUoUydLcvZ0tpADiuxhD2O5jSLuUuC3D5R33IUrj6zNE3vCL6kt
sizp1XnkjAmGFKQMHB0mU4dbtu9hyyRivIsqp9pc4Jf5Ba+MaBNrrVZsoo3R4nWamJBEi+vjRTMl
7CQ86feVE7lDmLxOtO6xEa7gUeqOjS9NJEbCh9wGIjRTvJeehl0QwzXJhu9wymEOsSIZ2vxBdAAw
q0oFJTdpnvCTZgLYa7FO+GYDJUg52/HkdDIir4o/AX79NfzmuC8RgWwDrpJs3HSSHFM9iv5mN3kT
gNgcV9cDUbQhQvBFZP2G92GDArLJ7VNF8X3cNd3L/O0Co42dVZ2An0XkhdStkit/TAlKfIlTWJuF
cEyp8cMl+NhvKTU6Z3iw5vykdne6IaXdlHQkZV9IiODLYc0PXSB6LsFpGBHu/7U03Yyv63c/UCVp
VayAmj+Fhb4yy0HbC4v8UghdmwyGiN0K0VxJohLi7k4u7D8kAPVlTs0k9alZkrP9xmkdSQeiS2Uw
MoOe2LkZtW1VIwcca5FERmRmCu843HAJFvFVA3kMEXWjQoReOA2824xV1enEY1e0cMoolIaJQLSA
wObsQIjYYXHNuqIzhf+uY1p+v7uayG4gr1XVN+v7mPdnwX661ZSqKxUDDESSuApHN5QPFVgKQ6Pc
BUOpX1IABxveT5znck4x6G9iAHZZZQ/cGwSSpbwYj3M0gwwCyv4T/L3hgvYDxvdhHVfztVsBUqzL
/RZZVOKb4A9K9y4qN0c1hPZ7UqpGWrRthgHFL07FBxBKR6jWWpIaZh94as5Tx/b0BFp3e8B5d9FM
4Dqg9OWd2amsuxQlyQ7qW6BmVadxGr3frVl5TeEBnIM6639vKhhLo0l2gtFIeCKwKZgaoYIkjeSP
Js1dVuU9S9ZYwGHNIGj/rvyyNKSNQQhUS7D+MZWg+/8o+pYAZHw7iJN2NK9ohH4XrxsNk+yWLlEN
hFZm0qYWjUileVuW9N88asW8Ox7eDz5DBT0P/YH1sMJzxaVEzBV3iK0IxGtutS/zjcZqYR709EH8
yxVLLvuQF1cIF89ydYRUU/coAzSI9ncf6G6ZxZeu45PiRZHoj5glpW1HniB9VpNHsovTYCCeCGsw
qA/4cN+SIxO8tfjxbhv+sXoETDWWGL8Rm/kGRWY+fY1V1txMz5O4n1buFupPkLwZQtKxE8wtywDL
jXDF+a6SvG5I5zKZgjrQ8DqdZXiPOvjFtMeI46N5o08+dCSsIc/ts2QrzMeAk2Pp1aw3yFElUhTy
W1ETt1EvdTrucWsHGd2X+tQk+W2/maIiBix5X0u7k2Ox1yuwwCm1cvPrH9+x5L4Y84qwBIQGNpop
SFZ1IsGJHthJBMWAOyjVRMHDcaZlrYKjiM6rd1Hqvc5zTRhexqcpW8rpfMcny447BjUgFL+vmfcW
QAANZsylMjG68QfOEe3/V82qYimqY9A0N+5aRgfsNdENf3E4RAVnwTaeuiDJDfuaE/O3bH2Kmofj
juWlFAAU+OjccVKNIQPBef1eAABQHCgKo6q4AiXx9VPaI6ch0QUC+ycgS8CLS959m9j321mgY6os
lzDKBvOIEb92Jsm5JFC6nHj74kkzUbRP/qqlgPtFfbYjNtmjp5H5gt/7kyNvKwfZAXWd0GkXNPBP
dZsiMl5oFMit2pZxUOi2FJQXRJXi9WK8WAE1mv7zyNff3EEamc5GtE709aBGkiq/51yAQCdYGQcL
Ly0i0ndpV3ei2o+WAl78LA3n3V/qQsl+HOqf7YWsfBA1DHF1ffhVUgAWaSiUx6Hitpa8EuCctjZ3
kLv4DMN1T+jE4cWeoYL1zVMms/fdxoNazXizJVcpzmH7e7zXwlrJSBLEjv543T88nluqxYAdnmx0
R/02Ysji0T/RkpyGHMbDyrUteVx8ONny2nofwLI2h04apAXgSclshwYC5N6HiuE7ko0BzlR3sUSg
C/gDnODBHt9AjeqL/bw+B9YqBoTxSs2rzlxnEDJWk2+Ydqzq/aEx/1IaplTILm7+sQlDDs+ano22
iK4f85g04cf+erJcOcPG1D9VDhBtdRVtBmGjktOnMINGcfao3obckMXWIx1A+1FyIKxFxxGbSqr5
rT6XUAUGNE9Q4KBu13X9kjK/ck4tMwoPbFVJC7rzQSbNm97P0GTHQg/LpGZUpNSoyMkxd4VT66HZ
OZ5G2xmtW6oo7taLzYDv6/v9tolZqsMrNaxuib8nZXPSGX/sozNxat2DABmw++pt8mEVN0oFJIaC
TltQZvJepmqIWQPY+MzEPapjd1ORtJyCYhgfSoEY400ZDLpB8j+wGIukjC7wjo/WcUls3f8WD6uf
QQgXBV8XeMMEg8XsxBt8Jq7+NpK7830PnpOsnH2+bOblCEGzdZGNU3QWWxuFIkI3zOFVOKZ6jS15
aoqmrD+TAHbL9N5ybMyCKURa7MX2WY16k0NEZYAwbqaX79Tz1IxoPpjYgF4Ds5nn1y1k4rEBpY2o
0ihP/0zTihkK1Wsqi/1MLJfiEuYBJDqObb5ky8zDpHrlBwpPPn2UBHihhERHgvh9n4RULLpH89yY
WkgGBfxLv/Q11gGxRmAMErodIC8LFmSDyta6JZaZGRi944uzFJhjR4nAejg7yIM+ixSF9KmfuvBW
+RgPuyRD9VVjvmDBt22QqHDZBmN1DzKxEazj3o3wVRU/lQGsZI1sHoE47bHJb49mOiNwSvuVa7Z7
9yZszlomzBnK1rZUeVNBwupyVUU4Siv0ALrEwwbsCYFoyax0VFaZ5I3KvHBJwyw/Bo6c9YKyb/N/
8qIH7NUt/xr2n2xtfpVkg2DbWqBRY8vobVaoOiqLOa5KXnjHTaDw9q67Jnr08jRZkiGgG2MsaFdg
hGPlsxnVDnOiXSA7VhvQmHa29wa92XSD9qeEMGZbWCd4tPpmDOYVKz+NO+5wcrX+l7KH6Ro8VMsw
YPmDOHE+bdzTuYMPetZlH55u4JY+iGeefXIe7n5qAPCmLGgZX7E7E1XUg93FrJm33NSZr9zkditH
8L9fModHAef+WPuuHQ2PahWWzmibyfyR4x4uEXwZxQKS8wQHi/ug0KS4CHcDOxncK6MHVJnV7IJX
OgRIy/UL+gFfP2cgGz6Ym8HP+2lCbr2RHte2IUWMJszXKsLazj4hpEse5MKHLF0OADkSYM9MzJ/n
PPbQWoZfFik/QNQXrsUeTNo3QYPA3OIDfoJ2clC/c8rwNYFAlhM7cwyKXG13HG86a3Mlo7BipGN4
L9coBtvSBOQTNN2DKEz6a2Q6e9K+8FHj6Fcrs0ESwHO2aa+YyDkoK4Nfi0a/8rT8B3XL92y4sNWH
P4M37OWe2TjPwfpbwW/DN42TXX9wGLNmKuV/pSwVg+RdFuClUZ+FmNOfUt004vO3q1vyk5wSMH1F
C2GQy9YCtKGQtRZlSUr6C4cT8o/5gpp9YpnOAZygDXlARYF138Go3Fig0TFNh4b+IqkNl49fGo6H
n0XsH+hXqP/wvdY6GfOGlgLNznM1KQJMjQ5KYmXeSfG9ugSJfSglv6DUQb/ATrTKLCPRzRw8VHGz
G7JgDeXzS3NWVlMvkNoVpa53V1J03/Si9+rFBnM3ASjM/LN/hb7XjxmzpiORKkpiE+ypLAYcBkKg
hRVQtL6Nhd6LXemjFvUKf+yFXSAsZ5txUPpGdSZwcHSuODgbXPYyGF3OQScsx810wFLq3RwEhvYb
g9z6qj7MhHyM4Glht+FCh5e2sHnZSYxARRmUcymS/PYvlrqBsE4SMu6KFPi2qIjoXHq6T70/B5FU
QpEvwYbpCbMsbVUk5OgSAngwa8gAHjktdzet+sQmsFfYO6Ff5I9YSdZ3XpdWOvUyhoo3KgmjZ6kk
REv9RwZ4uB8R2nC4UBKuGWw5BplO6ruoanz9kVYLBdtxr0U/XKYEBRbGiDE2ndK+Tj4Tjk5Xwkgd
nXIKdTM1PjDvvadH/97LWKanasKTY10eX9PyIwNCKTdtIiKGRiSIbngvahXJdbdBOEZiYgHd3cFQ
vchMT2K066qP0zmXPLEIIbfBFJ4nG5FnUQKf2krSyp0g7OY49/lx1Ue8GLuDeqK2H3zZQAgMQpzW
svQRkgkhFM/TmO5v1Rp4Vtrhx+MeoVyDW602LyHvRX7Rjn5fyJcce1jhTIQjGwXd0aW1+b37OkjN
AqXN05B6tYYPJr+TmWdJYRhTUyM9mP++8C4G5flLpnA4qRoyY5okJpLZstK0y1eX16Li9B064doM
b1IB5yK9Ma6pAi5s7C5OYFSmYMiIbav4E5KawmD5ikng2u5zUlQFfe62LLLoRk2GTm9iVf37sssR
RK0J80sT2kH4Qn8Qja7AexWmt3sGhjXkRU309Pqegs93i6jtPKXdiBikzBWGeATRYVNXT7qPS5yN
IUyS6DNKd4HW9bGJGSt1Y+6At7YYM54LrJ91HUVK1U5Qj1W7P35LbwHLWFhlvXt4Ha1H92aFOm8w
sgHVTFOHnr6SfjFplOuTGhfLvYGb6QrkdZ/L40Jvww/xA3mOqMOw3Uut1Qwls7Jin8gszZXojD17
bC7979vfbfK2rJrMwOIwKeGmNOcrwFaTvSXs6rspvYFODqfh29CrwsET65hWR356ewhan4QlWNuM
ASpg15udhdV/dciBn3c/DYd+0iHb2v+GfJZ9LenbRYEaROfdAZxsLBAzTcfJnAAP9GEFqMxpzLtk
Qp9HHA7w3w03eIs82ya0Legn9WwDXgWY+5RATBnUW73zdVuVUbjp/EprtcQ8WNR3Rm2v6v/vVbRp
HVnpUArknIOKqIKSVDhbnngePZN3WvgAi0NuJik8fMwubu7VZmoIoFe1tnrvlBf700YZdyEh0cUH
ML9hbeS97c+2N+XneYJLf34VC9gyWI1manlOtYWuTRHDQDieQ+26u6Bt1Khkr98RsLLWQX2k/gx0
cMJtYeW+S1g7qQmehqVuUPIcFSOer11Z/GX0qAW18SxKhraCRNyzrWTs7+0+zJ56Xq65CGyrwKzY
Sk7eb5VTRkLSa2jLs1wh5IpGF0K0nqpRJ/MP+M9izI1yktkaaahlbTa4OUj9VYfRlPHhtSGuMlj5
PBwxULKekwv37N7lOb1rDKer5MaljGrgEpElXrgrNV+BIHlSUlBNki3asqa5XyvQZ3WYnIaT0N2j
By2tJXY+AnLRVmTQjjwY64S1kqf/+0wA2lMOJDhVb9nUQQVqlB2B7UTWxJfSBgL3FRyoxSznK87A
2dWMOXIATmpAPdDW6Ih49A04ld3aYNoDy0Q4h843twjSuCIdQlMax5Xg/fWLMKNdtXUt/V0nmwmf
DVIgAEl5VNm1D9iA2SnwRf6qbAPps+ZDBn+FSVO1SybKqdpJvuaqHizQ1h7r89P4ZdEpcU3MKqKi
OiqqmDaj/4MrTAeqm1bHm8ghXuJjkNkU96y8AvD0HIJX1xSgnr1oE8tua53Px6uFCoyotTFK9wIq
cLqrcAEvLjEXQbp//CA9FrhUoBGLTskLaN+6fgwGeNpNiiMVjRosUPbJ06IZIWvxEDOXZMQi7j17
QUjP4ihor7LnDLa8p/Q7AUd66p2zAqpWu0TDpA6HvKGauqcQhDpc9c46aP9nnlgXWPwqnRc5vIgo
1QD4mcHqEm3Is0YmSKoY4HwiDRyDkbn0ZQxP/ogJPt7Z8zDhMcUoqx2ZF8D9FCy3uNFTaGZrcysT
Fo7L0lCxl/xjgHzBKD07csc/utMnNwOkSdeu7Bjjpc2Mf5oV1udqjJZY0hnKuV1/XEhEbwKwyevp
rOK6WC+y7tJLyJzjb3ACXDthIGEtt9ru+N7lvkoHKyJ+iRYf07gWtGKZW6NOOQs9DCBga+Tb3bKk
xzuwdZwQn+qC8gP/g2tivoI7tSv2cL2x+fyqOOKq6/wxXOhN6MiJ932m7qJ/wS3O/fpkGbZZZ+mR
uCwatiCmIdzYfj782DIGoo5aoppxEL2bY3F51DVPfRgKk+nD9D81wns0jZjdRPQJkMJnxQJV4aaA
7eR4+VObifj5r37tFhDIF/cZJ9Z+I1Vd8eJub0VHhu+3p8xb/NwdVKsKNHM5MRlAdbGbYZf0e4YJ
fhZ0mMr1iGbyvqZdadK4a1T+HYBZpFmlqj8qiBeMEHYxGDNf4eJ/DXUCfEeGED6nhpJtK6gapg9f
dsAnzmaVs8CrRTnLollWdS+ou9OLnTn/wI/rVKWM/dpfiSyp+CoB2MzAb//OClsWO+FgDIpfN464
bMinVcpaP9OUImUZvV2iH274wUitzye6Z74IljJtMR86PYQ7EPpg7W8yhzlicMXcHzfYoS76yGL/
a2J+d9cdgEy71c6dPgxub3WoWf7cm8RhTj4adZrZoXiiJv4CvkzVu/+OB3hvec8eMsDDVBa6fAlp
Q/14qP4wBr8LqaGiIg3ihPJY9ChzSiWpEQUW/QLGoKFzroUZRfPbpD3RPT6ssI1LliCbomhQ82jz
uMtR2jdXkFtrNxVdjrIJ2W7Xuj+xo85JoArywJx/2HA5cWVec5uxT5reb+VBoDfkWoVR01jTRwFD
slQYwbuUTIXe6LlmkxOWeiX54iGt/135HPfUpsnbKuAEbcLgugRhdzpRdnnq/AodtSClUPEohNEz
bz107kiLJ8X4AOfb8ZIkx4oLqXo7Q7EFe2gPuI3vLRY2xechOa4zPzVHSeARRsmtwUsHMth8IkvS
mW3Mi7L+Qx3zIfQsLZWKELo5ASebePQOsdBE6H9tyOkAQunggW5gamLodfJWsrTJIGTF7vm7WSra
Duvb3h8pQMQ1DkYQrT/63IgdecbtbelRUWN+2Opfxp8L0TrvDnge1Kc+KRxBJWYKSP3Xtptcp+oT
Je+rpPq6dRnpop11efo6zuEEtvxlTNEwrhyyJj99OHLa3XKQSjdpGsAkCgOEYvzAAFTD/FCRoPii
SAFsw0gn3OzXXJ2b/wBWt1qI7Z05kusMiMcIRBT1thq+7U9YMkFbOkq8WUfZztVca+ceOPww3ZKg
btXc2mQxfAXwiYGIMxev6EBmqzaRIWykK59I3mhpYIr07+IbvIMA6GT2ZhhdsK1ZZlM2YjudlxKZ
g0Hreoxr/98C6CENxQFkJ1VedcbJXXJVlRCRZe+8zxHWThNUz4lwFKofDtZrrxWnv/oJu7RRE1uH
65eQOeeNfbFojb4GcTuISMJlMSercKBYqWb3bJJeGMkcghfbXmvnDpwJ26/iNORyyEyus09W4DOn
wzumDojuUZxILNvNLNEhAYY+oJU/zBRn/qaHszS607dzrR0SL3io/by8ry7cCXyuyjEBZyvvvFRN
uihbtAHgnWXkg2fvRVwn4fZ1r9p3kLtTvKuFQt5JH427c/k1rHIUZLRbLtQF6b3+lYi88vGxjZbt
LiyJgB8oY/B+GtS4a4qhBUPtG5JaRD/fQILPXijae3bAsCIQFXZB2WuV9iUhDToUNWyiVXypZzCM
e3E7EM/eQtKih4KLB5nP3WRMMLHuVnEsh6IrDSWfbtGLEplLIUDLVPlHwmzunDk3aBHuMv7jpPrC
TwULiV4b87EXDddxB4r4jMeV9dCzfFdXJK2W7AffS/yNGmrVyYWxyuk/23KrLYY9gyo9cux3Ysb5
2VP1JgJv4A31NYOEqNSiRP6/pveFAWjy0sUbC5z3GgmRn7OK3F9662s5s3oH2aORyQJsQyf0hHLe
IOrdJkruF3zOUctapTXkH9+G7y9aGWmZMKA7X16//yyhgU8vpB8lL/P/KDXKEjpyVBMRAW43Ku0E
mfs4PPRVtQphz3FYdZt3DA+ciPt87aHSeTpBFMTYqhOK+B0YvHJEKZbbtKErnFTXfiwctV2SJKvw
kRnp1OmV/QUl0WE/Qzn2CR7/cHYMSpZ2ZR9unjQAI/567ekdTBW4yDSvsYTyszrqDA8W/Kuq0q8+
11Qzd5ydIBEowZuA5UJporuPAIzJWt/7n9ug+DkdhqXWkKFd4rGJEJj5Q9+PDRUMu3yO/aS1CCTC
v0VikYyH8RdOlBQj9OKAuFiVLlmXUrVkFO5zbjliKoaeGA/0IvsG8NRhN3YFZ3oiPSXfcgCrihYp
ZwdtA2k/RuanflvyfTuhBhO1H7Ow3sDhCwbOVk8Y+66P2KMZghRUkv4PQnRYev4IGGv4EXtgBoAt
hcrJA+RfNpO7ZmfpPpwSSShfljlTKw1xlb0arBuu/6DoqCWdF6qfFFL4AK0wlysFVxT61BU5A9wP
R3e0qBBCw7Y6XWxiJ9ae7GLe1BnhjaywjRCar3cmFo+6o47KHhwOwrgMlMuZt9MBv/u9yHBWoPOt
9XWVydgHhSTNmgkS+xB4/k62AiKazMFsvlNzHvICFncYxHwTxoCgxq7R8iFeqoMuouCoYNbdH+RX
+/slTow21eiKOBslnQ8k8Ceam0+sPLp7N26mbWgv9CuZuV87DLp83bldiTbDKDrjxnupBaiwG6Sh
B53G66Yk/V3zBliUilk2QieU7H7RmlhKe/XJNzNOpL4S0nFGoc8kcdfGtGiMai8hTTdybhHflrBw
J3nBjBkjEM7oNFQZknup1UyMk9XPVV+iSTFf99QYv7TPZlTC1hFY/sryR0S9mEesQ0OilrJAEOQn
s70LqlPTvSi+9keYhgv7b3uJoAchlteOBjvix4m+KeDTCPmGeptP4/ogUSs0EQYR5Z1IS5sovQBx
fzp83HB+IR56yX2sSxrwRwX5yfvBzo2Yf+1ZCb4ldDuVAA4ReAe03YEnVCM3Ou2dHpCDM+abw39E
nXnobxJOXo2FPPv5BJ5+HEdKVHqEcPFGbFly+SELi895/sxrwZiWdXFFEsFWtTUT5MhCoUF7fUvB
D/2hf76JcgjgD2aq0aUmgVCDOHItTysllzW7JHEQ0v3zYO/CGmRzr61QzXAYQP6idikth0kAiksL
w5Qmq+NwPfMJBMsFbCpNHpQf0ivXz0qo8IeB9kw4qVGTAMkdRwIkQSGHkehEMr0kSuQ8Csuhpr8F
jHCZs/0c3EIrWcDeDAhDV37MrP6aUX3dvDul2ARypjrSh432/+lLdqj9bXn1vROehA/7WqKRp5gr
4dWdzJIG4YryVf3fY7rIO7JYVXpBEjL2rnXYtE6SqDgzsCUYeSP5qpYAaZPbjXjw6IlLZfnflRlI
O6NLhglUxa6xfVtDsPKETHZ+0wVeQQWodmiBSJf6nnyrP4BQZMOWTFWxcxeIV59Kalu6QiqWYOAP
6p7uiLQtXviAxWkbmfRhKTN9jHjoVbzeHaQAl/adzVgupy5tb7KX0Z0QSEX5EpZV2bIwIiJJ4IxL
YZxrl5Zu46edpE22TuCvhqdxnElRIxXwH5vtELhLyofYw7tLzVtqxn61RtdMlqhsVg8elJmFj7kj
kOrAP3iVFUC517CPtfuxebvID//80w9Bjh+c45xydkn6BCAAdEqLmPalOeVXpPjqYl2vn6JL7heF
aph+ZgOKH/i39THF+dxrbUJzZEf5vwTAjNbsFqwT2DdeyFhLxXL1c+8qA0GyEo5u9pbJ0kT0Nigt
AXPMxxHvtutN2UNlaSP5FZ7o9/qdzJo8IRnRdEvLSILA8vLzYYsLoN8Yf6NkbOdE3C4mC8h+pCNd
Q2F5VodlKTg6nF58ixI7WuTx6zRvfEtTMrZgw44hlZsHGclFOS+4tpkJ/KZRpG4D7QXoDYx4yjza
ATqNKinQU946PU8lR+Dj7AkJ9vDVTw37LxwRU2TO2/liq58uYmXX+0nRTGkymVNUq6YL/d3sWMtt
RSWGVzotwIqZ8tC26n4sRcBohC8YEiO01mWPXpznrpH1iSYwxybQlP0QagZj2kLvyuX5ey2jVHZF
um/5Z9A1cUzfPWVyUf8o7Ris+I0DYHAMswGja6bNM/3VJqHgJVhohLBwey/kLI8PoaWhAYSHm2hV
ieo+MoEwb2ET+RhhXokMwQCRVON61bFaX8+frculkY0lxY6lADkRI6wNH0LLTlpI2TgSGCbBdhFc
LlLFYIB+s1hJCYH9zW45xINcGhb4f7mB0s19E6mNQj0vRzBpLLO9h+LZoeBMUCpl+xiGq/gUwYa1
EHSKQJCErT2QF9Y7pTGQfxfo212lxRql9yCYHj/10AuHz+O+jUMskjamsvF4zIRVQtmS+5CygR3g
QYRuCYt2cHwKc6eCf2IH40unyMOsBqsyF8Wxvv83EVYYMGO4tYka3lYDDRXe0csQ5WCChtj2X1uF
H4pI3j+qMK9NO0lMCxYWGsZBg1H8RoRSx+apnNVXELMCgpIw+z75QlNdY4nA8diiBQQ75K7sc2la
CLG162VZocaV0S0qmPm9bWSFCmYfQumZvgFcRrDz9mzcUv3ipt2YweszGGPc9s65H1hgmqgBXWnn
I+GBy/+m9zqEkiWC7csptMjpWzluCAfj4lg9LAQPgUWQqdBhPLPjjj4XmCR3MTaTrYN/FHmdCizl
xKK5t1jUY9S1RJpikEMCcKzcudNSrXPDhYVWvBHZKJhMv0r1Rz/nkicDB3KH5uaeLygM25BHfMCo
POvHuHqX1Z6C0g25tHAVWraZcnJv3gNec/SWkDo8AGUtpnTaNynpNGjozTeG9ezCsqjIGNJByI6/
+lTpVPz2yL4jMe0xXz1l2rfiSDOaXyGRzz+nx1/iGTW3ibfnl9mO/dvlM/8HzdTYYjNhb0VaFxoz
04w9AOIvDsVXxYOOQ5kv6ZSwtKbtteZ2MWpwwNtbuLrKSnuNQ8Age14pH31q7MqHMjf6xTpLKzU5
+SXdHJ0xglVXiXzkx88Y2GOJ/uWtyEhv5Cw+A1P/JV33WQ80mClhVTbVgQwlVk01o4XMEzLLCo0B
bLE6enourKPJISXhb4B/e2AzqxELxJQ1tghIB8tbJwQZlReMxSpgmkI14Y+X6q5KT6tiqb6lfPDY
LrajWbnCwmPEEMGJXRJAvQ9HTa+yIRUFOjcboh6VALFCvRgRE4Cj9nb4bqVEL0HVmQN4f09bJvBa
h4bSA4FeA/cJeT/zixE5BLRnnoMAfKvJaewgFzCGLt26twnHy6TOkhyp5eZZqE2SenKhnbsYmaCX
TSYuFBaeuq+03hVkdLJJeKMHDTasAgYTIYhmfPE7M6S4JzenwS7FfrkzQgFV9UgYj8ZLY/jXKbiv
rRjU1QU9x2YjjY3cgtvklHjW/xxqCluTkCD3mbG6hoapO9CmsiNEHrAUajLvOrO9RuC0ThF0q2Jh
O5i0jIC2zqBnjLKbMYhAknWqXu/CzbQDqM0RvlgM3kTCPHHl7xj/2lKQQRz1SfASp70j7fPheZCO
0nNzAJcInZJtJKMnSrXJSV1n6ASQc+t6vdrxj7w73YpCkuMqXAuQ+wD18kylKkt8ACr6XswexC1S
RDtMEhlsCaO6R2ccVnxhaDHdcPC5sBsiPJ7096M/iM9lBGWll5jXmqI0sAJgH9tGSDm4N8877glj
n8RhbN941N8KzBFirY+l/30y0tlkh1YsEhND4WCjTZNzRyyfrOS+/b21Q9V/qLBNW3jV4J7Ywkv7
AKnRsvmtaxFcjqv/fc0Ehq0ZY+B4UvckZzSNTMQUnWRvuAo2UHpkwwyysY71hYTPMuh6PpOov78t
x3G7eqOQeY9wH9pF+8yC44STTxtE9KF1drF+jlWNIJeLgEAVAnVk4LlwTIjYVBjzGWjS1qG2RUMt
MDNba8imVbnd89cu2x/uDVhtR5Cg0uCY/RsmNQWaC7csRu4UOLTeVu7lD9TkOONZA3GzByYWY1dF
FucNvydy8o6a3CAPPQg5wJBMjNdnRB5IfbGKzuwthW/+EFejqBsYl+WnzOhbb0DrJuSHZQBacTgy
i4l2hiRtPJ+haevBjNJGa/0WkySLmlARfE84iU1xSrNGzbAvKgodS3M3iy84g2iD/1cO1iDcSXqx
Bq7aZHTm8csaBgNhWcOoQOxxYFiaCisDa48EWDnY77dDYB2e/f22Ku2KF5sKcVg5fqtptur+VD6L
aemJS1zgTtGKrZ6/4jeM5abKkBKGndQlFycdTq6/cmL9p7y3mrlM1MVqFMjm5HfcwgRHftU23fpQ
xteYPlC4KXQlCRSqWkWY0KxoL5c/5XGoTi+N5NUBZdGk2ELIMLKkzU0eDSbKOIdJE4r9PZZJWZtm
stAXmtg7srxa7SOT91ovsfH6yltfZ5UQOw9Xbg/EwAdre4qLLZ39OTTkE2GeqyUGXUOQQjCWcVpy
OMogxykyc1OWOHVnFEPPtOjzsOUa/CK3ZllpC5tQHa3tNDYtId4ag9QTnfE1El37vgylaSsHiAkI
hjkrvBWilSOwO7PVjw668ZrwpP4NEcijAWRwIXgaE/otRnmBgvP/AW+2Tm7I6VhQb3a6QXqKjmSV
lJ9JnPbNWAz5z7TWNmkiBpMjpWbDn724IJUziFaF0pBlOLkTddUXWbyBkx4Qbjjea2nzC18BWEV7
n0ekOATyEFhz+IRKQvMEAjF9TZMA0TaMOW7qeGWY8uLsgqLbdgySOEjdvZUYZ5ywRsW/U3RidqEt
p4pCaPrI9Yxqk+E6P9M5xnDX89Qsox/CgL5s052pAOI+N8GYInWWDTu57YSzUxc0qWK8g7wkomxE
QHh59rsNF3hgFzrKrDT2B7usYtbdHGGYogrSYVfhND3+Ct/mVSxL3iuT+lu/d82xmc8c51PPEoze
ccsg3QIE2p+pQF7qQsmjxGcYPb6V0PVZIVTRRNhsOQu/W+3DXGcynBeoBAZaraDKFb+EE9fEx98E
T6bPUeo8ZXHttf+5+3LNgvzlAgZEcUY+0ORt2xWopfS8wMnWUYpmPgCZG8Rj4wpInk1SA+XvK+E1
ERiA0v6xgz40AYO8LXONSo4OOveqVxSuHh9dehW+yi1kUNtIaedmpBjZ4JojquaTHifShOBskHr+
ZuwaxUv1OcznPcOsBJ4JpgwglvAfRz6v8ERgwLmuxNYL5OcfCaSjvgs+D2+WHlDdHJ7DKWybqIDD
lxPCbM03/QG19H3KEzObulyUgH7shWVzmxxzYMtbp2y5P4kGnDmorTTZ75egpR6soCm9O+tMxEQa
qx5AQqeoiPRkEuQnhHyu1QDW3XCi+zBCRs6XqeHBVpNah3408ONsxUINzeKfIbPpfRoS0qfC8r2u
f8Gxs/rAqP21Sq+wzWXGNXwcIGRl0xGyfkaJ4112NbMACBf5GpFTYzoGfdOpHv3m+H+hjyt018BW
RkVGRIVTmV+2GzerLm5wo3MIGfYwrJKnYgjlYdtSnAz+lVNex4DMQzJq4dxYkfpKdSGLRl/VVT+o
7juHxeykxdsCSFWYW9FcQ1zBVdJcZbOm636lH00jx1TTtnUdVfyw+deWWxAtFW31nebPm0iIEYYH
NIjTe8EFQVux4ficDCbYEHz9h2M/GvOBzBJUwlbX7frzoZio0Irc374i20HOvmOoqkgAk91SHabo
p154RzY3Z0zKBSg7oNYr9Hojjce9upHdgIyd4NIwcGWc/qj0jK6zGoQpmX2EY/g/d3rZHW/Hdbnw
54iFePU3xDZVl8/I+8bHstZpdPjAOzOLFXdtbouOoQvqPuqFaDdFV3NaryclaCOEuA6zT/aBzMfI
THGR1mTd7aRZZ5NSNOMPjuHJN4RJDO3SjIdk32KDIf/MKrCMFdbBFlDW63KUPhX+lsM7edXE2Uzf
pkBexeWHnO2X8lywdkGaSds39oTMN6GfvPfGk14ssOPr6AkGxQUr2AjTRvAZi30Byx5cDEcr13EW
7yoh7uiDCdEIETLNOLuQlfnMHRJRT8Hesib97Ld7uTsh736sJjGeTfXTuiLYfjM7eUGJsMNJ80Wi
ZNPjqxvsuQ+Tt+Xrx63dSqbVEK/Ifhcq2Xf/S6leLVr5Ht8bWCS4DBx0nYj/HeGrnkCmPVsqzEjk
PkMdOQ8dijIw3IG32Z8OZutqPq2/GLvhEJjr7De3ifRafnwvvCnaOG82Vm2BmxAMUOgO2V0u36ke
Uey/00ogtZFlA+Lm77H+N7klKhEwBkjWjIl+58hMVFlhkGBVsG1JyGTRQoPKZmKyKKtt6ZiosScN
19eEwmWbPYJZYMNVr7zw1rJBUqAfuqukD98Rmcm3R1AtlRjLCqf6CUjXjyMJ4tvRgGjovqIUVr+W
xigkrUgDAqNve9ZZCM9wvL6oMgGeHcu2FJatjaq/HcQsSkwpVZs/JbmJxBoo+zf/nmgaa7DIxVu8
4cnmIu/uiJ/9akDn8AhPABSsSmAxw1IpwQeCaEeoJRMo0eqvtwoXWdA+hwb7kwyqlHXdBl3oOTdq
9BY2NWbT7BmVoRfUcKRVWv8XJszkV6veGi9IzG1mQFVmABTayDqUqYSVY1pTSv1S4HRPeIwn+zfW
m8rXDB2tOcdRFF32dNVUa0LIHZ2tLp5IW0/NL+95tKrZiUNu5XEU6jsAkOsyVt2ypQxoXFRYLZ2d
XgJkq4Ll0otCNAFuo2idl4QGCu/oiE1trfXA7g52fa6Q7Ss71ZmJ5HkOUEVc+82G/4oR4g6ht4sS
0Kc17G5KfEiZEYHbSO0fPT8EyF5koFBS31I+vcXY6Mdk1c7ptkJFoFlysuwzU9YOx/238K+Sn4pY
MiKlXp+Knzs5qlGIPoZdxW7XFb9QNNHvsATKglXapRRgfAQNlJ7NUdWQbL8XWQqf7IScTqR4r0Mn
ITD90WWQmGSuIcFVXX616BevybWyjSHYSQoEdDDFK/Q0u99134GNDK51Qp2HQFnGuTJ9NwfTWdF7
ifFyzZ/NkNYsRt0Dhtdr/IrIPrHqPRiriJbNxvT8HyGI3iKUFDxcHfsAojSIOgg6F9GaF9oW+3HB
vV9gLjtILFNlY1pbFW7BJrNk49gU+xJ3DJ4VO8ecI+jbTt1ANHL3KNfmv+gYdhWNDrlj8RqUx6HY
9ropBUQj5ELsuNI9yS/Wvyr7NAE4UnYfK/t4P/TdMB/TRY4SdqFqVyNFEWiXn+FZmFiS8YyBiuHm
nGT3/BXwv21F259Bf1MWi4rajOmfHsG+3MOclMKiMuJ/JJyIxosmjus+zGOVEm4OTkGKJrDpI39f
sf1ebAdtYseGyEZh/HeqAX6Y9lP4WCQS075bN8agOTwKdMF+amyX856PTXAgPPk5RZVE05vgHqYu
iddYmSRgipcGvfxsN/Mdmc3TCEsLRnak8y/Rt+Z0yXGHqMxwF8x+u8e/kpNGYrLG1bkhGmhIfhjP
eJypVmr3V08hnMk11ikgc5jH/Q0LSVy2Ip3s2oLajyfazocp0EIrTgjQVt+AGmuoTxkyHjtxAjZd
3eCW4a8T1rEjZgiaqH5eHkHPlMA8+hexxgzHUsxWpD456f7vr67UOS3pfQ4hamZlXQDsntmnGyMm
Z6pSrD7Mpf79DvYRITo1Y3FmpAyznEFvD/dmwRen+waLQHYi6xOm3fWAwu7y5b7Lddi1OqTTe75a
xSpyEnhuKiHsHU07S7ZLBA8yiXHQRPnTTIBP+/18WWT7U9pjLVvOpiKX4fNKp9NST/90HbxyiwEy
8EswyjGsSAHsBsj5wlQgLPIJo04sdnd6LRtver3vPkiiTDPimLjumWMJBKaDJA4/AeP2ImEk50+D
oshLCI5XREXQA+IN1S52dFiYiGegRcsGpxWCtUqCJdJDaBrZw5p4sEAP3HuWfn3KFDhSzkEc11Jw
jzthoJ9FbdY+1hOtwm/LlfCtQ08+gltbjKOiZuBC/946Esj/JC6t9w6ssGcc6pTYKuBRBucXl9HW
UaL+hHg5wwakbrCVqPICCeXfkav6WxkQECDeeQFvoQKFACosiuOlNG3MkH5amWj9nOLGIbfnhF8a
VakAELFEPH5Xe+XXzXg1pHs+8x9JY54izY4D91Opb9PL00xPYkHBd7N8mlTkro1QmP8YC/l7i+yS
ek7aHnNLy6/QQ4rETCGoTgN6fFUZMYTQaIPVXdRBbzqe+GrbbWJhZe+oofgmUV3arwoiVWRRhmf3
f5vkFUAZVmokU08Ou8u0UJIbUNseVa+XGmnBAbIQiZt55TQqgMt/2b6F1Q11ZObcVcAnOoH96z8W
bXh79VALe1Mz8BRxiQ2hT0P08+R4uTHrTfO5dIRjUb6C42Xvz/p6mWI4JmlWYZpMLGvh8QpaSQit
L5esvztuJWKAZ2zG4OUPXz0kWkrlNfrydIWZ3EpwDvsMwiOqSJoJmThx1TCoFGGL/bhgAtM3BOtU
pquKmPHgnT75XmFkEG57dFz6oJ2XM+GmBI1aPqjpNhCGBdDsg57DGZRMwDQhg/1yoKTSCAuv4CSc
7MAq0b+82RTsBb6B+tjPMXbnJkq/s1xap4keqyD2fLjmzEWoyRemfH4HnHl2iXkgu73nZR0MxYhj
E2ITxaRQOegPUasAdDWU9xIv0kqzI6VMisKiNrajb1bXVPgKi7atKsM6M/u6NYF0vfWyEeMsyLmi
oKNh4UKW14Fo2zvg+CCxSn8qB6L3aFY8F0ycFVDmVrb7SLf1pcY/rMPcOIs/gVOYWqtcn03ACFFo
U47eMg4qV6mJtR7gitB7GUA3u4MDpFNJ7Rs4mGNo1IR4wS+wNyXk5WF2Yhbe7yjsLVlULTcmmbYE
WxnmsxAdDUDA8IaNYSP28s/Ln0tYt90Bd++1LYyOEWMK/s8zQt7tORiGV5UlKDEl2/rUU2mWfZ3A
gUAh8tuGsx1EUUf025/HzaCkfzF0LxoG36fsprDSkMZOO5Y/dNOznHzfq2ODep6cJNB+c/hE/hFa
87+WR+y1l23/fCuI1RADd7J1mIYDWVMsdcfS5IK1w8IFR8uqMehc712Lk56hDfCzOhbc1oLtKRzQ
9iavrP5V08HX0JBDrtYrj2Nb/iVPGkjRjXqz7TEyicKxU2KPSak6jJsMkXKY82NkQIkd2moqqByd
xKbMM2Plgryl3kry1PcQYhM+NUs1YwurrWetmp0NlOkLtJEadxaazlgzuigoPS7FZcLVgXCtKGca
g9/P8Ch0bLabpUbkKeQVgXiHvoK6z90Hp1Y+btz0Ljs+DsEBnL9+xITjr+EYo4tE8TTaIaXrWQuv
pV1SHCU/MFOJdgKhUzaWS/uJ/DFhLCqSG3oONdWkenPMapiKcy1ROmtBzpFo6mOSByn182+33l+j
HKynlxkmzbwDyNqh00bF1fCUsnX0hOmEOlWKET/qmyKyApsew+KPTMA6IGUDDNK8KxA+LfsHOSGG
86Jt4H6zTWoadOgjxFGDPcmtYdczvr0eZDvE1o37aO67EN3YrC6qi5sDJVaEaPQfg2hyLLN3rV86
NewnkKJQudap/BHI4MiFPocQx/1MD3v8vMmW1mf3aXF9ZKuAtG60ucmRspc1gVE3Cq3mAOgOeLBS
bpvq3PaugghU7Xym1Gm2WVhZsTtBTkCmrdUcfF6zO97IO/x38jAtY+qcEcfKurFRxYULfDAg5HU7
hmDoxSSoV5mSm1MczaC/EFqiH0hQV+7iY+KP2pMEnJvynxys3xPiAsBkI72Sv1uDiW9mDUXmZcrB
lQfEEUfISr+5NKwZE+N91tPgtQqIVHES0bXmaCJAfnfObkLhu8LZzWyhaf9vUOv1HN5WUEfZ5q4S
eREM5zotMXYWuxQOZwaFbT4dOgo3WP96QkpVaKmTn76WqZZO4cyEMzWCMCtYVtL/GIneju3AwmcB
q32ZpobpKS6UXn4ptUAqa37jLunKoRGdjCJofYmYuXuJQC1qvHMbJeiL/h02SH0vovOSwdH4arbf
x69aJTDzDxaZZgdw+tss6o2pjZLO3FIzEcsLJSpZIQhmbR15yOvQBJorJc2Qv28etrFpcHkg56PL
BDaP10IyIX31rBzAIBpK4i9n7ok+v1Yav+wg9Pq6AjPMFvJSDD0deYNdiol5kpAHWNky5Kj5oI/1
q1bbuFNJv5swyajTGujnGa6ZcnwkuHXfmugAzyG6aTGiijQaGHtxXvPUFtExBbJdqCoCLrKn9aYe
2EfDaEbGrvu3XOZc/QUW+MAwyUvDxnMdYxxjRFedtJR61izVY3D7aHgmE14MidLA82pG8WjHzwff
2HBzgb+j+4tfVEBlwao92PHp0uR//a+hRYfkCU8fMXl48GPdy8TyjsO+cLFhzObkpGqYJXnlrLC+
mXFXYimQkKLSlmA6FxHkVnyMnypJFCDWw5+BLFh9z1951N5xx4yx4+3etXrmn6TlkAgiV69t1PVn
GDohErM5NbVuY4PdnAH6P6Q9jopV9cHPaYWe1WGqQSZT6W/+mkskPUfhhtcTk3BhjBZxujfUbsnH
CuCNh/OktyvOwh08VbK+agLUKnBhPCcsFc/IOArYGEdQ3fTYftfeTIOUF1FdB9r6jVSIHhb3Tqx5
gbJxj2IsIHb63pzzsXrq/EHXjSIf1i00n9ZZ5SDFPSU6erSfYiraVyl2fuYpMEEt3s5P727mAL35
+HdjAemT5ZhjnxTeU561/znYrZYTQIa1rzZsRdorHEYPZiEXflIZTBp+vPKMmOc0XKTczrtcgqWW
pRAO+GA5Pxe/QiZGDHg8yIFwk87dpkHTBtJeSvsi/Jhl0OW/xmGh8UYTHFEPtLMrCWpTBMYb+ObD
RqQyb24if0lioEReMHMV1UKtAKLO4CBlZGMb7y/1hfC3bAzGjym3BXdoZlQOi3vnd50BTf2cpQAA
DVhw3BhHz7SZNQcZpjU0r+JtiXO7Xl99EdhHZKB3f8GY1aasFkSpENpHEwsFZBfIx2VxgZhsbuqZ
d/nVm/+8e3bmWj9PXljrRj/2aKjPKS/9P1yQLOzprwXgz2JyM0eq35zw7Cv6oRwk4TBy/dKrv35a
XKR9/YdVCNhs1Vsqwf3oli0EGh8AiIENwF3opFZSAoCreq4H3Gaqt/DyZEBMfnZLrGms0JM//SNl
Y+gjdduA7pWTl/8Xd/PZownHeWFM9x440ko1eJuQ2on+0XrWIoJtFaKxu1KmmXSAGelQsNRlnu90
nk9RcMiKMncvG1Ge5eO98NSPvZJLLnbD8/qN+lGQaqWbTcK1L8OBCw7agCSXyOrO7XemsyMNjQyp
HTMkWmybUvQWV9flervqmODB0cS7ivXaDi9zk0RIDnh9LfG3OhastJpfpHqV68jwMZwszZ+AuL6K
y7ACpoIcacg+BFLSlxra3u74ukmIPFMpmlEJ2WrRmyrVCYu8B2gtUNDAOcRFEkmelQiirANPCL4i
1sC5FTfMDXMOJi/ahynN8syRlm+nfWCFnYb+n5LC/duio6MJkJwh4V5H9iG6Yf+Mm+LQGjdmaBCg
5TxE9KomsW3S8VyZ4fU9gixq7+X5kYVJucoRBWlXNtrn+zDurxIn7YpkkDlxr1lF19ZLYOBGUgnQ
ip63l6/QIa9kMoe49ZW8mbXi1iM93uBJ21xZo6zZYAvKD2asVnOZp/FHEDpufIUumSLguFkat42Q
yfLVO+Kf0dZAnEciXtckZ1vrqXtiBXCzbKFvHafjnUQY8Dw8tDSBhAEFDapP6S34eMrX211r64Mq
X+aBi1nVdV8zruhzkeDdufmczsS87BRxpnxwRvFPQyNeaF81oUgYUQHxIRdzUxxLeBlBhTQM3huK
NskqRkQ6bWkT4z0PkeGXWZbCxH1mniWFWOBW2MpvoeaDmpFrR5Gy/ajkeK08itQvmiwjI0JQzY2+
DFmwBzqz/rdnIKFvkP37HCR8MXNH2qdwZPFVs/tGTK7Nb4kwUghMbmbZtqunSO8xWt9xVLgG3Dlz
YvPSs3AGTUc+4rOLwYaZumUlNHSHadVv4hDgSCIXRsH4Q8vbi3DHxE/TgtW3WX0vNxDT2Lnq3IHj
sZG3/MYfDqstNkhBhFiRQJUWxVDS3Udc3ozF5M5JYKOo9PPKIhqHQJtQV1ynA6GJUYUgZTfwD8ZH
NowRWfhto7wOLbzUlf6XX6ibNZlfrrfrRUp8QrqRKlsP0siIs4kIqQLPAaHA+JrGiApWIRs4c8d7
43A0CAWnbU313BMx+NPnGniVKbprsNihk8j+XyvR9FEchyXVIKVGYg3ne5HKqrdfT2gblDR69SNF
aZ5BIgND/w3aIxxu/nCnbcT1l62JxiJ3fVW81P2tFOHG/tB18/Gt0uI5QhJoi+Nhdq4d1Zp7IbWr
Ol90RiW8h5+I97tEpKJMi14PbkBPsj9wX3gImDM9kp+jfw91fLVZh7gUP6CVlmYyAgGjClYFx0q2
hR9IFM7caE4+5LS718DPcCbDZa0SJlV3erhJ4LpdU58VwNObFxsZxVDPFHb8uoc4vdbsn+eMoSeo
9bmtRIgdEA8uOIiECtz2I07EfGfPCPivRu1pnGWipwf6AKgoWFr8BCMFB0mAEeDhLNqx7SxOvejD
y74+dhMG+iTrPuawZBL7AOyrjNWU3ZbKdjSFbBwx3+H/or1ozDM6Z4W6AxcJEOzec4TK7er89lP9
Wdmdem2DeLzN8vizA95VXncdxq7kLcw71YI/QLBsZkbO4FX5/AVAexbVFZqLrDYH+JsJRxRS6qhX
jhQaFs+VyfeLJw7gEgOUUC2bczBMLBD2v4Bq6TSN+tWEykpJ+loiWmfW5+lZUMXdjly/O7MALwVm
mNRJP/hMz+rF6nVmx2ZefOvek+cZhXl7ZYEwvK0DNdCrUDyS0WFbGNMoLb26icUyz/JmUpByeWsP
/Nhv6H2MmX++mo32zgdPAHSBDzqRzUzP1NhnEWl1zA8gojqvOsM5zVpHmS0ayvGf/mzQ8VjDcepq
42YQK3tm33eGZZhc6JUdTUTt1QuvvTuAqDuxaFK/wTV8jaDBgfZv6LlmDQjWyb7oUifT3/cxZ6hE
57j+bu+3dua4pAFEUmdBAZhLrd6fDvKeM/UbWGzCTnMc09QT9hRsxP649kQenvrWpjXhhEF534GY
w31b9cRz1S2ifHxDDRojcVdZQmasdFPC0jGVUq4Smu0WdPD9VBlkEx2o1qITZrE8JAE8L1fKlSZO
lU/ZEAFjQegJk9AgFGVNC/iJxCCfpE6F5/be1Gga/y8m/ViJ9md7kEWEqPRAW9wj8bKEJRQZ8qPh
llh11rcKJBDwXs1N/YszPHFJ6aakyHI1MsnZvloWQw4nme5TM2+uzY4+EHAwb1TR0Bk4PD4R91cI
nz8Ja+OYzRhs1GyY+LPCRcjXszAHPlIsSpCDKkdfZVqg2dSkrWqCpB1bpqjOPrUAhOU8Iw7TwHyo
oz/O1CRf/VBeZYLzjRTZXpWNASoMOOO5qnkA/2hEYEXS3xF6I67DckNx3zKT33a3xDOPLn0rTIv8
/xhSc5mTgL6IIeGXNnNSmOKbXQrNFG4Qadf2UPqRBBEqNO3RrmHylVXKZ42YaA6k10g+/bG36m66
Xn6BkF9J7L7uYGDKLvRkdtJoTomDScvdzrwJjNg+F3zex2Z9It6Rk25Mz0+UCYcVwl+jVjLADLzm
jRjvjnKEZA0pfs9OP9YzNjRuNyzWnVPsHhzLsDBoee7BzvtB2aG7hOmjIZVA6Zd5wdZWh2Zc3yoS
+h+D5hmgd1OWvqE1FBAGqQXYpQD4MTE3gp9cHMKXXg0gG/Dvx9AqHcKTMTDASjWFm9Wu31pX8g03
FMY5J0QGvzt3MkQB7ad7IjsXwPfVGpEuAk/P2Vk+gHGB54GVDpmQ4UWCxzq9DFlvuJjTcfq5XKjh
t+IVLUNEN9rVIInJu5ker4OcljG8camVlGTN6QPhEVJ7CnBrjqxRhtQ2o/iO7IySiQrD4+yoW0Qc
D6v53AMVGsEOZeLT6nky3T7maK2rwqIpBmPuHJyuORuJHObnEuCS5+wxdaTJNsKLS0wIF5SwRgmN
lXWV7IFxiz5ZLKi9WIesNxAWYpHKBZA71vajMBhPd/27mrsbmvnowfhvfPkU7jeIp2RJj7XQkFCi
5L9e+Lxq3qVVX6/AKWiPVTOZUd3ncgFYWAJsNy/P1s8oivAESPYO65n3eLcETvk8gOm6KUReZW3P
4a3Od6xSTFkRoyz3isifSz/KvNR8+5kWweFMoZQLciSF7nnR5+MdaJ7rQbbMWKSBxNQezUkHjP2Z
tzp/vFXGCmULOwzg4oinR+QvigijYPNu4bW9OgdKWcYSJlWK+itJmJ+6oEiypH6pxtFR0ucjgogl
TENPxGtcXom0Ub3mAaWU3OYDu9m2ojayFouNDeFuJn3pyxjU5Vyr3xopbCKNy8V5+wuWnr97AUgu
s6Tu9TBmJ2M0gGr3ErJ+LpH2sWWGPuhTK5FWUQwb5kM0WlmcCN95iS8rNCnet8q851ZxzvvSZ59J
pAPJ8EaFvVVjpQuE9H4RE7G2wmqR608eykGUZtguFDUaULNEbeLcpvxwCkDsBFmQYMdgk/Lt4ull
6qaxBjEf7y007JFHKboCMYM+Yq8dyC/7RclXMy6DfBUEaF3V2OYz6nlMSxE/mfMF11OUZ7811B5I
k2lHU0lBcN39GMMtIB0QzTqXkVL/nhjBRCWEWcCOvhxa3FE/fsdQ/eUKhNC0CAFbBQ4KOjcaQuop
XDt1dj/hdbd9xP82jPm8WBIEngeAOIv6fFQkBJce2tKQn8ZQH++4xGpeRsX/8yTnENdktBFYYm8G
JpL9z5/Q8iMSQBtlIjR1+FEdxbqAvbfVbns96SjTIJv32pIXX0rk/lD0v+Y1jFLojWMWMON2Tu+M
aJvIvk9ptFVwQ/oXRYmV8LtY1P4fK+a+ef2eWanb0o3uzLJznp5oRE2jMaLxg11JTk2BROTOtRpB
v3B+8FRFvrl8Ff1rdPNJSMzC9XOBTcTAXHGH4kBArauFrM72GY8OPtURR8KmJkB9VkowLiRZ0hW7
59vd0wN7tx4Mvkc37Czd1uoaBNoG1e/ZpY0/M6lDTWBEYt15tD6HFr5wTucI/ucrlRICuKPHdBc7
tXOSzYRVu2HN4rUwFbG9BsYfiMTTRKxSIuVFVFZoj297ZpKynr8Ijq3DMDCIP23QRYLvjgqdzorW
78gA6DLcEY1CTZji8QX4qHbab5KclP7rfcSGgfiBoQEoJDQ1ApQCByF8cJa/wJctW63rxwMxC+Ck
BZbVdej6+/Uw5DYFV5FBKMHz8aae0th3P+wIY1XQHqd/SneWdQRmuj2d5G2ff7lblwBXcBD46+0Z
5WtioZg0rXXVZH3adrcN1rEx7T2tOjPhA+fqxpZ550no8Pp/uQFbP4lHz5xhgaWpI/YOQqUwgN/U
prUAXue/bYRHTJPQa6982SOg8VwK1pruYcktf4Dgb2lM5jiZsKTEpyrdSjoxYJhOdwwCubci6Dww
h84vPYFtFizt/IpL/o5XicSJdGw7JWjFWJyMLPBLZGfYlZKffSpIol5xcnKHJRij6g7PrITwSYKd
CB5Vexrh+iFzR3vZyviiGcAy9r7pRIHuR41ohUOqm6cJyb6+I5CWUC/OlCdSjpOt4YK24qoeKEf4
2JteyzNQDMLLD7xspix1iWjEg+xlB2B0MOZkzww8N8gy0Gs3q4os8iYCJONAW0yKP4DnOgKjwO98
UroCB75840jFjYON6j2QTZ8uc8/6+XC6hP24OoNP/gNyYYmc5fLcARfCwc4RFR4j+yUEWvHtvEjM
AkQoQaaWwVHgDNRTBChaNsP9nvVvJZS8DvDpkGZpfr3NWZy6OYlqkRlVguOY27SfoCLweqzGircZ
WLMYESlzamr3eZePbQ8Ck8oQv7lkkmR0Vp5nLzGw0TduKi9s4llz6xZQGH266rGrSLOzGizCe40y
TaunREnQPU3ULbCfFCPUJ/uL2l/7rQ7hxpDArNB2OK8hjmvecEzwnUUZspUVM+1SSm/yApOwTO6P
uHG33GT6J4GA/SgAoBUtHBodYoTF405Ox8uVxnV7gq7w3uKPmj7Enr/XKXv/s+Y2ai6SUNT0sNLY
wKWxdvFT+rWBkxivxnoSj1Nvbss/lBGU+Ob9qi5fO5ah0jia++aDlPDLd8Hlcz/e6EOh1AtedxiW
F9VtGRiAQ6O0NK5WZhs+lbCVp56sEt/7hkcSLCVei22AI5go5C7N9LCYvFhf09w4wpoQAREBDMX1
MTW+Gmk7mzmNL05JP/kAXPCLomGKHjyjMqOBeUukKJbtuv19r5IZkQnaQ0o3udVDBa9+opRrYPHq
B/9u4kjXPHNhYPvyDW5oIj6nPsp3q56g88hZi09GWyyXH8MYBIwmkidAl5C1xHB/ifjQDHjpyu3L
S+CN5W1khig9KCTg7AENEc1xiXlckK9r3aWFgO1U0S8ip43/QCDmtFn192s59ebDysflSItc7jBZ
8bsPBrJf+t0FfxswF18EaSdxCS+O/2wZ+WpgOpn6lLrKCuXlvaagC8T42flTH2+BE7Y/t4V3JuSW
JhIldlEoXGxPozn2XhI7PnPpGk6xf4KJttuiHFzqF0WdA3dEWlw4M4ItRXlg4ecmFQU+pfjjnB8K
YJEIAkpX6j5kFEm5M9g31kTHpIhvZxzCfA12p2/99YpnPyOICFUxVci+pon9yo2W4DsoJFx2V+K3
D+EBuDA2V9/5D5B0HL8MFTaYtF8vqrUCJCafQeIdj9/BxOkCe8b+5OQhnfDfLudXXsYPxvWe5HlV
THD++CbUROme2wd3WsnbCxIFiZr3Kw3thN0iVHk5v9Asb4vDW4zL17xa98PUlUyph+ozP40+Sg8s
EwK9D884igTQMVNSIMzDLX9IhwND0dC65C9zdthd+F/gvdmXEqeN4NfGbx06CpbThMJKI4dyr53+
Tc1MivguL5ROS8bztIDF3+DN1z+PX61U5En+Inczr43q1EM9gvlwML3LO9NkyuOTfiQv331LgBb7
+bmWgJOnRE49cLLyLjDgQTh6Jcr02Q3MN9OgevYP4y40Uv79xRql2e17Ai7fdTHgAW5yXOifaOJH
y6OZJQBCazyKULG/TGEYsItEBFO7ZPFcJ16Lbq7ziOf1Kf7gqf6Z85K4Yy8O28toDA+hr6BP+TSb
MF8ehD/G29eRnFEdrgLwKkq4H9zWme+0Bu7ROzuxI/ryuUiACNUm7k3K0+Kt79xKokaQdwtx4j7E
kFjq/5j7UleHH6ED6+RCVKN+44TdcW7doIjrpI52WYA6yRPrND9s5nw/ON2w4Lo7coBjw4ZOrD+0
4wvmm+ukiwUD963meUhGYBkgQbExpcRViGxLO+46XRuua/j8JnZBpUJo0nIi9aslfaEuwGfmu8JL
5zyj2uXoGTyBs2ufa6W9sEyRTnPNiGuFDQkZLhmmETZI6nSiOdPIVYq9XHw50Jkl+OUqU0+JPqSx
JuR/clP/5ZCuG0G6mOoivaBrJdmGVYrKsmh4xx2JNLgSZY8gASWV7qLVV5KP26YWxts8YE7iqVLK
J4PpuVspIcqa64++RsU3cQDIlp/R277xXR+Jdnhel82dE0ApgdS6j07YnXgd/+U+tLtxvmvn+Hnf
b3VX0sr+hkUy9Ix/a57hoR4iffKAU2gxCF7IRVbKPyeKQiSpzYZeeM/GvUyNO7E/IKD6fpb3kjfZ
36kSj5+pLSN9Z/GKVyQ89BKr1zinLWmBe7ojVk20a+n2JcXQDjJcH/rcQ11hY7FRv6D2MDUydQx/
eQ6J+/AKIcujsq4qhEy9UE7cmGb+J1K/WxbzcucFXrelS/vhesFZzZluvzAU+cXOpmFD9wx714Cr
ZV04c6zRQYlUzRVvizizLtXFvxeBd/NzW28QOfVy62dzGCRnmGOfaLsQysNq8PW3eGk7ltGNK24j
vtB7dZlGzxxDfAWgbjsArEPL6ynO9hQT8V1SRyUE4nUxM1wx1KiBXM5Ka0Yq+1SVBmSIiGU+3EVs
dtCxdqfTN6MPMVGdEz1G7hq+TsVaihhC4YfvSNbFru3B/apjGqYsB4p921Vxvh+YzTLMnaaq7Lw4
QdS+xBcJTRSWQQenrI3hlAe7H+QkyVQojQZtQjyggd5lpxH2bGPjZwJf1pUUSfUag2488ZY3gEqa
jHkShkr4ZxqJOj9uARDTGTLJrweOt1+aIdjhgPMHNlsPpMbOhFOlX3+ugZ7r/kMphItsEhs2rxCx
/ZZAM1whhPFLua8TqfmuiLjKlZ9Hdn+UCU1I+Sal5M12SLYf6iFLPR6YRYI4dgCV2jdeuIUGLYAY
cbIcu6i81mnpBl0D7uaYijzvExuGHSR9dH6UyEvzuyV8ys/h/9CW+t7+AGwiXRMJb9FsP+ZZKJyV
yx/vnR2G4ncfmaLZ4lbvkuGwj8YackdS1DWom3YPHG98a1R+jS2GjkYoAfQDG6u3JYFe81l8u3oC
kOH9LpBtPODSliEZvHCWmn/THJGkOY8ttF2isvoI/BVfXvJbsGXjZ0A2DD8Cayz31FSXLCf4MOFP
je2sVFSfe7tO9hwqA7v8fwL7yBCmKSH3DoKuH6vfwX3A8fRHKXqm/GCFbXgm7tgnYm3bl4lK/uts
Kr0jTLF4YCpqaB95Kg5i9URu28Hw3TzV4g4tVpQPqbWTKt3RsnkqbRcn0xma6g/i2gx7uIcC29bL
/O8ZhW6Cc3/cUAZTKufppB1zMGdrIaxHQF8/eLY/T92YQIJZiWfsLKLbGQcw+5PxY+dXL9f4dTA0
TK1NfasqytF7PaANgjIyVa9NEBLKwHs/lvfoZyIMhsyoXpOwYSoQ9xR4ef9R0BtVe4CECzgJFBly
RWUX9IUjGAIjAaTb6Vng8CvcPO0mKy6qxrIjzUN+kSEIkWPMfW7RLqhEA6N+lJb/uANjYc0sYmXH
VQJDticlVZmSxk1z5eupaFO2a6qMfVwmlptAgXmGh0znbfUeh3G/iUh0ekcqFA8Q08f83vNoyzB7
cI2iqGmzrmE305rqzocAfGLNlICYX1YQXQ3OW+bI676yLKJWZ5VscON/f0FU7mn9sELN6ZcUwK2a
Djzi7gxov9U9bf+5OSZ92dqShzF8O6HMMVVNPKQpCoeIMx2GihVs3/HG5yGvnWW8VzIvjN3v9/Si
XHQYgHBlC1MyR4CZyejosaFcipIz+yvtR7pPSej9oHjlb2w03jEfQu5idxPAmaJCDtgDBwA94qfg
NFpxaMR7809wviC3iznBE21D6wllrLAOYns6ICjDSw6WzqxrWyoBIyKASkGhEy3i1tXdUGYi1OsO
BRyl2YOdwHEJnAZWXb+iROhgASWmR3mM8Sgz5XhS6F/iU83DOZuoztfv3yMNAYPaUyiIVhzHZcXA
mUlpMLEhVCLzlsXageNjElMyYDMJR5P0s+KKuZbflij9s52aPkLb8PZVdb0/15lGkPT29639CyAG
BXKRvfj0wJa4rSCI943IcmiQZ3m5VRwJlfwXB7WewLnrc8t5UkS4YBN/Jsg9qhwOCuhB0UFWRR36
Oo3GlfvTK21rl3OX/lhB1fr/tH8vCwoXCMinOirH3z2LVDNNsKYUCR3G4gZtQabLiF4MCX+H50r6
ExGvy5xGhIEDFqLnLgXabHn33eRIKwrK+s9NQheecvbe0P7dau6IXx1MwqodP1RdrfLM4QKUmk0R
+KW79UagAXkP8phUKwC1N2XLE5HIZFezQU8Gzfcw+QhT4vfqoezaLLkqKluubacxiDC86GhE/Mfi
vE83NbXC1dGb4ZW2oDzYzWhavc7FcKa5RFLbUk9WexJ3XhsB+y+g7U8nluJIShgyGxANTChu4JET
szHFFP4gjvdDMsFDIqmVOxxYYNB9R3WOTBp4+b9K2dCjuyXlukNvY9JjIL69yRcUPqVO0fADSP+V
7eOI4JJC5wZJ/zMSS1zso1vj0T1idrF7+OXiYuEoE5DyhFxt1LsKOKUu67pVUor/eRm0f/a4BoCZ
yEx0K6mX8/1SQhaF7JsMus79SjoDgV3yA21qXVSvpYpBAzGVq734fby+OmuLhAKsQPAHO60SYKLh
IkebJnOJqwP8F4TW4Q/i+2MAekT7dXizghU5aPHJqAkZ/jPwiTbmUOhe+cU53wccpbM6g/UGqSYd
RtCOaFATK53nsENLX50zr7QeQssNjTlCkmWiXOiz+j2Jj3tpeocBRt4oiKyv0P0Cqnl/wRIFruWi
fcFWBowhZofdo2RqiVQ88s+aQwosVp8b2cgtBZtZLLEALaZh2RLA9eYlclNGMA1RH0WZxVnOwVPS
JBwRZbAyVNJKzGjn+cu3V5ezMpUvBgJRNFLTW99U4nfUd/G3ZfDiAte8HfbW0IBzodqOQ3wuqhB6
mV/PlREmOzjSGC0zPDTigfd0q+tQsV0+OMMCY6eJSqu1li+hoKkoe2M1r6XGCfgoOtKqYjNw1zJJ
fOjrQKm15E0+i9JUV27VWvRM8MH0gqrwfFvL+ceh+9+3k4Ld1ZfE3/hWrgEQUSIAFwbPE5w+ES1O
hY/myACJFyPrCUS9RDaGAfgWqVXK54FIwOt9ZyuT64fOO7lotAaQq8jJeBkBwX+Ak1fGXJ+Ltp/V
tx+cJxy3njHyCRzsnBO0hplGInqXE2yYgcuL7P/kVoIyw8psrUbFrdvlQ0qHqSc2rcHxmp910bwj
IewMRItcjG5GAl6tjJ0dt+bJwu/xEPU5IzDbFQjI2PqtfoZOzIU9kMNvxT0R1Gkll5iXwouJt+vD
fdrUSUZSYKxMRY9ytQCNIWPj5S2K7TE53ddNfsSLTEychhmNuF5HJo9ZBt/dQw4nbAT7dg49QVL8
2H3wzT6wNJ5wYEah4GDCZqjTdDtY7ii+cexRnRWL8aClLDt3qDyyj0xfDEEh4h9KbmVLrIeJdqJA
U15ie1cTpYoEJRuCxjpJDi9axOCLx9Fc6AWOAa14DvJWctu/hIyggNUQ0SieN3As5qpU6Wea4A8v
47x4/fyQf9VBkamNGtcMvwHPRJF81OWrpXFyjRhW5iqE+nwMIDrcHKeW8BdMWPlE9Hov3j/tBoOO
Duu4AiTkG6/KllbBYE0ntq4STXXA9dilJ1grszGqALI7LNSZ563EkpqWZzJ4Q9Vc0dbJiGNEdglV
iL5u6OeQHJPT1INKTSfxFHmDQzwWwGvfE/K3lFNf4SBTslJ+zXIHbkpA1ZoQo7uRKwVesugwiu95
fzRhqC57orZaLcmEGsS9m5rSoyamWA6Hhm/uoN8GIWTJDrdyFr5tax4zQkjY85Hk0dvY2W4O8c3v
/0mA25MTqqfpcyciaaMYBmeHVX+TcG7T5TYvZ4x/khp0XBd/fho/goyjGnZED86SMcpntNHhgATS
+i2zBRcRBUGgY9tch28X0wHePPyor2rrs9oI9yhV/DEYRarkYSV1v3QB94Nt7pMWuFANnCNSggxp
2T1uarjjIuDBwhlq+c5j1hrxYq7onNeBbO9qhrZIEPO8fKBWpIx98eQ91lKrjx3qEsLHj+6jZvEi
BkcVqPn5r4caxjLS92f8C9+2g8vUcyuW1n3CShn21ZYLAG+cm8sj3KaIbDrjjNRalgCZnF+687TL
nJ72v3n+KUFwknS9BXyrQixb4NVUn0OkuoVk0NINnlKNDXnIrv8ff4tI97iWnQz5ejTM5ZXIHMbc
HkAQ3Aj0j1L4y+XIM5x4x9lrv6IgaPtW0rlL94Nxx0N6Dlmsf9/d+gBB7k5G9zVQANejSegnUVKp
dZmXwXDG60RTzBopiTPgkLFN+HKWrdxnORgQY0D3j0KEbzLmQZbhefzmCYQRp2y62Dxs1LDQ5rAs
DTYozUxZcekH81oYUYRqLlwHdozUCNo4PSlV6dUExWLyDF0EghHQILiEh0ozmtjjrBTrv16MQ1Yc
bvUQccOlJyw+Fp8jxJBPurz3cFsD0NEmdN14/Ywu1sT04HDcGc/d0nGj+A1AnI8b8PhiLg1M4NOm
opNxCOTs4tX9cAAAEGNh8C+5YhiSBf/CzYQuSakRh1jJARiQRTGGK0aZbTSypJFuKj26gPX+3wK+
KcaivS2BL0QECf1h9bcw3BOq4yFjTYEYKrQPBzUzyZUgw3bXFtNgnSmFCvA/jhhzpcrtoEk0GOdK
11xED5UJoUUn6CQSO9bWwGuSiMgXx2kzzt1FCUVceS+pkp3M05HHfveJb1d5XKQBk7fakL/LJ6hN
SP2H81/sNxiukIhvq/RrIVE/27f633jYZwTfDjD0WFi2/COXHgWg2khK8SS4sBDCVgsLLbAoR9iT
Mp4FdmpmR+R1ve1HotCjDlZ6GZRLkxVIoA4XTnAAG7ar65heuSSpuBX3CKXgSIgXJAZHaq94Xs+a
L5Ye86MbKq26WESHGcK+xI3lDtx3UssU8O9wSMyrBRI3hlgkg007RwQZ92s66QGpvaTzJ57mSP4g
ua96/sztDVfadQDEAgT/lJxHu1CGlfYSw8BpTFL44rJ5XfJlMclwNa6Aa1OnjvNQshLK2o7f7+Ec
TkLO6xxusqHUMjEpFsn4r/jlTEDtA5PLf0LGGEv2YPnA73p2QmiWcGlbB9QKbswOaUH5gA2WfYWo
qIWxYUU0c314H7P6OkU9Jdu3ZfpWA8G5MhoVcJD6pSw6XRX7BdDaXzAigwWU6LAMOolbUhYCYaSU
K50S686xjISNwDMI006vdTeHrEBrVoIKKGIsgPVFYjynsGHTHHO6yW+fHvbmhxxymmLBQ6npemor
8H3IFGGUlP6AOVMdjyzwtWkjJPwh9CaSx5n1S3YR5GXxXQYohj7qo910DXvcc4R3E2OKq9pI60hV
/QWrH1O+K+jDp/VGJW65EfPt76Hfe/VnN6RVhStJNlqGZDmBo95vymUFSf8QWTMJJjNyQlvtMviT
WrF7221Hbf8ZbG6BKzuLcKsfXNJk5trDx9dQ74FnQqwAZcFM0N/bs6Zvqnti7thHfkCdMb6/vP9I
mDqhZk0pmJ2jCc/48BxdEuZoWWMbfJ9PgnLySbZsEneaQnIcOjWNsV+MBlHjxbCWiwXPRPuBE8dm
/VMwm/GhUtvRcvYuAdra30JNAwN9Tw6yzr0x4fQotkFjmFqZkK/vsRdkKcEwEgAqRT5Nq91BBr9D
j/hJ0g3Wp7D3lW8UUKnn5+vvVTI6/HxCRERaDWXx3zaDrDNxEEQ1SeGte7Dr3dsi7OY/dOVUReUo
9awTaihjUIFvY3peQZSv64znjIfDFx2FYCghAObrjfzgXovRjnnhvP5YhIOiUXBhwW0iXfkOIH/9
lHCfqTziH7nWsc/DO7J24CQpOjpDzlgy0NAjN2lRxLO1XNnhEJ7kDAb9IoIlfR69hyr/lEGHbivX
a0gpD9MMcrKsC8AhoUZwsdEJlBpKK2FV2JBXLXWgXIwXIgZsWLqWMvrRQB7Fnmgw5s11E2/llcLa
Umi0e8hTXnMnjbYcmAai35M6BJXp1z8Y8TKULcUA1Bf6bjF6Su4cLtaFnrxZCEFpt56iq6dE5zCv
lnD4wc8LhfOQceqi1dWuEl56i5kZmKbQtoIi2IP+Ap2CikOGUicomaDmJQqDS9cps1AwfpzM8JgM
oPxMhMGaF8HN6B2tnZmBo64frMyRE3aeC83SnqRkrivg9bx5/UWGEgvXnJJpDFhVqt33BS5lqEkF
42IgeZbO7C4dKfxWzWv/jz1y04+HjDj0f7ZU9IvjRN341P3pnDag4Q4khtdBWlcHND+qvYFbIms6
kpFqAea0t34tWJBxKGZ7ict5N7fpJse3dUjHeo0WnIIbs4OKozMVecuRbrguflTC+Mt22uhTus9n
Zy7k10MRqDSYrS8SKSysI27D9pTlJoBVe/tPm746f5Va77Yjl/OOsHnwBCCapJEUqe2VEjk5ol0D
uv9tjJHFOuvYhom1KUx3ETsri4ZXZQbwOieLP/DJI51XSU+xJI0/HZPcsj7YClz082hUm9WNeny+
JMRQJiyIDBmegKhaWlEhoR5DsIg65uM3zjBlsQ6gJeIGXk1Y1o0Vwy54xxaFNpOYpYA60MI2Wdqc
+DjxmQ//Xqzqd59j+neDmnSxHj+ZV3Q/XmAm46ySq5rlN4+CAQoOmIwZxnT1q/1bL7w6NpXyvJzv
NOd9TsG/90sTzN3IwZn9PMCNxr8GBHMOR+0k4obR5b5btGjupfOqRNBcuRDca8jTT/ZqyOdfD1lL
sSMpS6ke+AhhriGR8T3yLsThE0uwUUBprC1zppH+2fkFacS9IXK4ykGw10Fo2ItDTfZ9zmmkaPBZ
g7B06m+dMf0HiLlmfV90lAlRs4MBlPliTEW3n7+gCM8dZtXggNpiZqGUP9rO0pwyZo6rNQrRoZP1
T4ibp0uJWLvH67ZKMxmqmB94SmPY3mQ7I4+EEZ4PMwqDcnbbhY3h2FhgA98YqKJBXmdGO3C5VTGh
0057Mkv0uj/u9T42F8FvQcLtaGIkeOWXPTcPXTPJwnb3RYGYNprQ06NHX1SDJqd5YYqRy0QmjHuL
XM63sPdAHg4lYiFeBQ6YVF+ir38wYBY2cJWiA3oJMW09yfc31EfYzZG88tGHTOninrdHSWLOfMyq
1/6lkyMthCdqlEZv2u1Es/BJNYUdnydycrajMnuTA88wWlEkn0c5vnTT66ndSO8I+1egCqTyTi26
4y9so6+n1jE28T4mVoWXM5FT+qcr/WjI2RIkKAgoBTI9erwGf/qa+H9N7nCVQMtxUb9ibRZqbC6q
ayToVck/lHZ4lglkzVCaSMWSsOD69MBE+Z/HmCZzpbMOT9ulyRbCasNJUeD0exr0CdMPPyooA21d
O7HQfsnBdaGPz3GtsqnG6VIk97nFqoVJHgqHcg/ojYGoOXLaPNpca6bcuOkbwzZSj+GrpY/+xQk4
e66h4n+8YNHq6dGprV2jBu6083WM1nnrK6OLj1HjilXOzSPJz6bGTGCxR3mztIXS4gzyxdtBr/0b
HsAiiOPe6sgC1rVJBydJNXRrsQ249qt+qc9GdXC7TN+ndCzahdiN0HqEg98gBKsSLMD1ap6X1w18
1XTUY7sGOj7AUyZ94hR4acaY76sV1ygQthPCrmKpuYQ1k5GuLcyTjXbc6IC657WOUgeqWboherRU
liHTnZVlzfAlyNHvNXZ5NawYlGjNV8on14l8GSNtMxvHKG/pUEkBVEaLLVV0qHf29IcyV70d7FYS
bBm8t6dVTIknpFu7ciym28xL+lNctziKHrDMrSQ72MCFLdDA2L9yKaCm/pRGxoD2bKpoRqcL0vOs
UEupq0uTbZXSUzNTlPRktd8mkOF3TAsU6u9bh8D14Ha0vR3Mb1sDxd5WnBi6PXPiyyeDUOWsXvnt
YVdwYFZ1LXriLc3VTqKpICfgD1HZOkPi1d+2vYVFmh3ckvI19Ll89z8SsoePoOxl67ZkTcI9Jqja
gtSg3xdPKs8FMR538KhVRWWznp68fKXJUXe1bfw2lLJDSjwdfcB1gW9ANG9zUqxXhNhDIr2+1GlM
FCrVr7yWUvsW4DyFt7vHN58RVeBvXPJIKxoW1QoWubntDpggUq1FI69c2eGFhr7jmHxbBAFQJceC
mPIBMleAoZf7DMvKvD/b3pfpZjxeZTD8JtlF1/+xV8+wioPNwA0s4/pxB2aESPuVDZ5/YuaXsK1v
jQBkYxMBTo/InjnigXOfB5Sb5lUGaztUE3qT6eiDDFYJWgwe4B68W6EvEgfR1RiTucHo97c2M5/D
ZUdx9pWVMquyB3OLalswJHAWxL3ng9fAHrzANUaG3LdyIDI8aqTpbo/4R0qGUTg8YI1aovqdr1Z5
FBvPJEG7lhWeOcYnb71gUptFP5IMZLj0HdLLn/e70OconLi5qFEkdHCtqp7QB/2Je9Lpd10ETjQW
jIzVjB/lX0314M1lvzU9C50orqogkwF0+HktBPsJ9D5ukMIRhq+YfLa3sej/fk9RORrBiIdUclb1
x5Whn73gPh81QpHJMFUeSyGx7s24smKsEPUs4yuhR1BADLufOnm997uH2UwDkpP8xY4wmw2FoEg4
kVgIIB4B26YyZWSi5/snzGcox+BDgp/nTPB6fvZLcyGOz9la2Wr0YH2Kqh575OpLmwT19VYBqMkS
IJmWsE6tL4TtZUVox83nSfCbICfeFA9VqFx+XlWcBVQCNgcICm0h/57iWeqer6//kPkuUmfhMvEp
+3xZe+99vEBnd3YGelm2P7M/aHK69EUGwCg00x+/+BNc3kmWr/2u5cDzp10/QOsamTfc10sRLQlk
s3UidNIaC2H+HLzudz2DYH1yXLy8gQ2S2mltKhGdP7ntkOz9rONqp7dZvPgTWArCUcFJC6/siqlr
padAqLaMiZF1timBPQIF+rJ93owC5PyQuvOQrmXBC9cwAHxLzOXfVNi+ZKFNISmBr26AwxVTibrU
4KNBkhGG/7Ey7JGLDHFq9FsoE60z18Hea/mvuQO56YCh9+7+M/tot9Cv7eg3S3E0NPA00ZlhovTJ
VLMM4c9oW3QK+dKZB5nUHLJKskcRZE9rrNxSyS/VydRUPMHdnDnO+jpufui/9Y+tMeU6sktPZ7ZI
FZFogaGhTznWdBTfAZLEPF1QpxJL0FaRxG/uup6N5Fs/iUzYQIr7grJ4MXlCUwuKempxk9oZs6Bu
QAfFY17a1Y/VPlUQIpR5eVPZ0xX1uyqEFSPLIoZOIEUnZyb2ACSKqlbagn5UzWdkIOCVKKoBamOg
cM43X0K5EvNUfT92ILdB5hZKyhX4AWE3TVif+F36iTSSODMzR5ZyEv3QIpChiLbpPxnpT4oflOI8
XOHYdLyFEQ2Y2pKsStjlASqdGGmep8iPUwzW2xnrHbqQ0lYtfVwYxqLNKJlaJ8AjoBwJXYXuCn+c
5PWsHnwuOzfXX3MSG82MIBoQfqx99celEocAZibYD0goe98iDdVGERayt1KqD0xRDmPQ+1bQrLUu
Grb3VqCIkWUOO/iXFlqGNo0bP+jYlb8SJrIzGzZYXgNzHc/6dW6//O3ROoCuXMnC5R13lGe775dG
zJnY1spb6Yp4V3tLrUSmb3f8qscVlnGsS8UkrbRzQH6qWzwwG/OQVCFZ2lY1gWBkvfyeXnYYvtMo
m16LuXcVjljI7gyMYvrXXOu1No3c6sISExDzSN9cOCwbUsuPxk7irV4+uEupBFk99/oaAAPK/dqi
THEBbSTrrnsO764yh6FN5fnKEhO6ijZaR0++Uhyq7c17dFY44qeUVY4hafxcdj/qMCIFH5cNzMxX
LrC1SWh8NARCiN+nLWeU5pPs0H8uxlwMXf+MbkVeNK0DJT4fO4MRzHcB3jZHs82KTSY9CTtcwRiF
Rz93UJmRhrCfqjOpe4ZQvjUzvzCF/mdtymtvXju8rB1MPa650F93UOHomf3bOfHntDJA4SKTZC/1
butjQeVBGcYLA0SnEEZ8bQnZHw6yaNzSDpFsMe42Z6X9bprG8SB8PeZlpyIENFTS+TT8pYn9k9Hl
vgybqr2lXdaDPHU2zKuywXW0rg2mjjFDO+mOjY2yyqyO3r1ee+i3eMOVJ8XsGZnKPVAOi4jd2qDt
f7T+i27nke/Pn/zQYCuoJ+814z73wFZ/9Y2APYwuJgpfugXVjNmxt6n/UTtgk4mCM2SK152TtsVB
rmR8walwpwN75geC3gt/9MhUsqgsSHqGr3Ek/9jlfO85qgkmUTvMK2bCIa5i5et+HTHuxClEZJFr
clqyTc8T/uB1IH7q4kgXexdVdizxrMbs7c/VDCK0ttF5YrJywD1pLnYmPck3FC5x6rN9vIqcWvyB
iYj6Y38x5aDM8GhOcdmlac2/rbDThv7udDmtwIFkVwG9lzGfhrp9jURt3tNr12+B0Kc8FRwWQXdJ
h3wtTF0JFtH29huYzDkR4hCcjM2wkaZkZiplAIlTZsMv0NiATzlyYzsZAKJ2fdmwTwDhmJnbofml
oPvfyNetf5OOG/8Yj8jW1lt/hxTqpkMlpQq9zhS2pAv6oDWxnwgBpe3Cfkf8CyGBgVAg1TkT/VWF
FuSWo459w4g1Zbk1dfN9RTrCAYNZn6C4PA4pLDNogpWOI9XjZTVvS0ok9CNGc6+zUR/L3QLPrh9M
O9O//V/TV04YZc6MNg/j6FzP+5pw9VthG7ZlFxczwNdeQc39EXPAMHYipCw1YfOLNC5M/KvcKPLA
fhodU3oGw1RsHUUtRYzpdfcCYQ7MF4QhmvnT9C+Lr99JEfyx9V7jl0y/117uMxUzD+8w+fcRQ92V
41F0jZweS1X1kyQzD9j0OidmHCeCEnOd83YoQ6DT5REix2ro/4Nh4TxNhL/xbQh8hvrzDChndlQd
TmcfdV9iPjWY2k8/Dui3pF1HJjBABBwyM+BKnM20xq/IITc2f2mhpezBT733G4x7f1XjlD76Sz6q
m+5n/MpXsMjTifPa4jJtdYJkcPP6doMEMV+Tadx1fxYYhEDTIR6U8QofgpThl7JfpVc+9RFh9P9X
5uvZgY1xRuhbzwE+jb6k03ybHvSoX5VFiQAmumyInk5PS3JEQzcbGszMA2XhZRGYE3IUvwIyNzcM
n8s3/epodnWzUe/hc2lPRHEeKYUhtpbcUjExGhPrpvMwHh84v929F5xkghsWl9DuQ9XoPtnH6clJ
5spst8taQgxOfJgv0yFdaQ2/JaiZ8oygm3SWlfJxOEXU8HznObPj7LN7dEYVyrUcYNBMFVvSMTTi
5caHAKBZa+h+bRjoU/0QE1h+kELFY8V8lzJRUpeAPeyeygTV/bI2wbUPHpfhcyX7UgHAp/ua3P2Q
foEsFEp2/oo8qlKeUVrBB24edCexeiCSMz21XMe3dxNkdO2z7Bn+Rra6z1ATzFfQG09hBVmVnvYO
dPAskH0n5CNlpCpTUwbpBxRr4VFEYXfNX3dqjZenDuUTeJaw/TVd1wI/Esz3JmLG4QZucMPZ6eLD
4KboiDLTUAUVORtgBwp5eszK2bzSJfc5aC/dazowTgW5kyp69JfigGS+KV8DqzhlKUfaqrg8BOAD
MwvyUWSWGfLOF8+7+B2S3DmuLb5uLd7ES8TlzggXWb9sJxI5R90et90G/lQO+CuyHBIb4OGojMm5
TN72gXrbUm8eE4jgnE1t/VU8WYiyU+j+tg505IO6Xs8F/X7e1Urd13JLpho+M4Kb2cRdW70ZoqT9
Fo+9UmEGQ/D6LVP22vXpstZkpM0zC2t/+9G1PS+7w6a+kPfz0F9YNnnHGw1eA/Gwk6kAftmD0UjP
YMH36v9Cv8LuFc3mUXZCVnQO/zwQvh1LbTYVz0z+/INZAcbKINn5d22oJIGbpPo8OeGtjhH3TJ/s
vfPlgLmyaj893oy1aDz1wEW6YBBObmeEo+ZBqRLyl5kclfdkvTHnKnZx2BP/YMC6GTFz0tVg0aey
jtwm7P3v/jVhALPVLNoHgtqlBiAA+9d8crvdfS9/nEgOIC436gId+WrKTNpHeU3Lo7QlD9BzJFOL
FyjMOgq0k+IaKyhVpZrmO//vCY9tlna/g/lsAKs42B+ygd8zJFnCHN7lTF1sHKTJgvi8RfGnJbH9
7aPq3AbfJaIWgt2a1Ae5eaETf6m2hLF2XG/5uYrCUouxwhIHRR/KqEEzKX2sdZZstuAmfNA7Rc6p
rc3d3tFnqLqH2ybW+COOMUIdtvLwxU8uDjcp12suYbXkwkEi7CsUFmvJMNYEf2sm+EwuRx1dfviA
EmPJn0ihqH9CjC1Cb07myVLStJu5+3l+KancqC+lXCHX5n+OzeygX0ndf2QtyETHxYayePgzUmUY
ujPCzLnYWV//JpqxhVq1LjZu6fK1GU18SVok+QCtDD2+cx0i6To1DcrnBrAMB0QE1uYeciaxmg5Y
j5IyBMdj48pxUnkypi3y4w8XXbRN8Gf6sPA4uRkGWZIdNwz4DnkBFgEJhw8jPmiHP6FVctRdULNf
johpJKC/Mk+6RkBveI1iG4o0SS3IWBy523G0QlSzAsAc/7jZyY49CAk4oV+7NfM9r96I5w+2XGdT
nJhL6QD5KsnFLqCw7CBy0ZcK09UzZrsxdxNAgcm45GWJUyxTjk7n1U2vGt6/o1hDF/n+PrQXDvzv
n5QUP/xtFjCgcjqPiX6dH+cd6L0gVH2dxnHZb4m9hx6AzY1J3gtwzP0VQK5Z92Ht1s1dFhC9JFbF
NmgIVOJrVxFvw5o3mgtAGAxcmwH+snhOMEZyovtpDhDT2nXdIBCbqBRO4MHPEvzrN8m8gaNxk5wR
8+TKcZGQGCISJgSbK72oFBVM7QeS61w8fSrEV5MMR8yTVc51Wzu/ON/tkMQxg4pwxfUXYba6r43N
ramxz6Hcm2opiXV+bLI1KLars3Id29NCHsg+RW15QFH3+oSxuHAz264P7kWfBVjFr0Z3cczqcQK/
fYfWhqqqYpHlqMEJJTtAowCmJf9gF43htgBXFvvCY/HGtmSSNUghA8XMIYrFootNmlfI4ZqBhFT3
L+znH++f47ErtriKFnSQgIImjhhpP5iRCsns/DLHLSjObRTYfXiEagXs6lk3hg5u2EnbhQ5SuuR5
VAWeNBtkorc6iaDbON0SFcXY9BhalDGHsHoLWltywed9UkRpXkn9fKENXls//+rhBhaJty3AC995
0gRkOLflvpdB7xaYQGutParTJ0BlKvN3H94FLIavThJom1Nv6b16RVQL5W0oHebcSeAzJWshIZIn
5NzkOQqOExvmGHhKIxnaFETAcKdBpZFb09slamqkLCXREiWu26RVyUMztKPUEQ8XXjriaXNxi8zM
TmvpYtoinZC1WRC2fzDyD38V7OD+Fd1F4qH0L8nCBy0BdXSzXw1vRk7nJMeo0Vy71len7GZuwU8R
ihjBVsr0mmykpDrsu1pL+LXK8wsRgAxM4xNDu5lISUbY7jstGiuTfKX2OeZc4tzc1mAS9Q3t49+B
NY941rhHAFVKIWiPWYuKjPfYn06PFoF+8HDBixZRGJID89pGJGJhOk++0Y7PeDWJQ9zUhFib19ls
doLzoXH9Z0QygoCuV5UV892A1Z7+sDzET1/rjty3TN+EJ4CSNI0TEU7RnBgbvaNOGyxcDeAw63qz
n7OEQmvd43TSbTx+cLsBxyN0kwF0SFm8P72qjpsn2D/1e9SEOZgue5uMPsrASYXZW/Pb/zYQj6gF
60DehO4GaQpWOwTQhKYrlUXFyXPPySQzAT1lIUqZbIA7xiyTgk/bDs39Oeqq/CoKusV5xnk5fZzq
SoAOQqY+osuWeHoKDT2JVB1C2rFk+zP3Niif8AJsLNAM6epDOMUevilHbo3fqNUBkD+GGTq59VuP
mqoCLHlT4EqbiPEfbpfPrOwn19FSQAK6epq2kMmk9/phUFpFYgY0N2h24G/lewbmbizQ2FCT2Tpe
qhOfv52/dwLMuNMF7FLrZldV+IhwntdPnlx5o9S1vIbSK2gWiV2OTkjT/WDJw0PmiGHwsk6cnJ50
4dihQwkTH79Jw6Cs7Iu9Ac4oCDGCU9EeXZhxVPz47Z5ffTSY/jVNth+uKbF00Ikcp1th7cJH3hlR
jnTz7Q6otr4qtk8UCUsrSOTSRG/kU3W5hlDlWWu8lWHzVya5gD/Qm07Sw2H0u4cxu0h9jutFk4ya
6AUEjZ9gLdaFDwyevH19Px43St+NO/1y/NAuXYub2dmbX9dzJqVn+mfnSrIvm6aXvxmEHq36Y2ow
I21OVXeRz4G3dxNH5jeUKhoQFrmZvVPH0Nq2bWdIzyDeSsSC5+pkCBVPBqno2T1eMWoYE1lovdMd
GClmTPm8FmJh44pSvgKkU5mDkHlNOoOWx49wSQbJUQavAjsPP5vYVjfJzGHF3u0oyJFfO5bCHol2
g4s5XTbzK9dNDW274m5vSMZZnpaKGoVuyQHolJWq9ORtSBA0pYcYOwzxSzAYJcX5clTdllbeVte3
+KeVA6vtA0ucWmO/6RrkoeDvZoCPMyBK1X+Zdb2qieH549jqHeOEoR3nd5WAGN6hWn2xuesXruzt
OtuMOV0H8aTHd7NHPmDNYN/0hOgK0iyNIVMkXqDjw+lTuhnpF44d8ZDRREsHRQ+bCoi9ilFSTlQt
XtFyEY6a7Ru28FEmIsZZEsIyHRYEbs6bVS7qUeJ/QR2gQy69idmnmtz04juiYGRCbi+jdnJC5qQt
N17DAK/E6An+FUUBtO53FIx/Rno+fd9zTynrMWgdQi6naz2hZMEy5iRzKKmcK4d+n9K3JEdWgRR0
63IkEcoYNHMLPQ1geSgFz2S+N/5jyjXIDkFEcQ0H3UcLdKDRydUiKkR1sCbNGEgMlteLq2IDjVEW
EB94Eb589oiSCWU50X7XRc2DNjxUvEQCeDdMVJTXlbzamT7iqJ4bf/Ss0ctqQMWt7YeO5BurILTR
BQ5E9M1cm41MCDsrGCwZkXDn7vENGoM7y0vQY9qHsHSWnrum4TMaXLLjJUICpEBnvCawTqi514jF
Fr5jvBxuFhmowAVmtgU/atE6NKjimLR1VBoX5+FMZayPgnib/sGmKE4vvDuKrsuERn1g5OQbX5Ig
ICYCMYi2wu1bQyN3HvdsC/fe9LP9puuGAyUP5lOaY3azi2gT94UwesYqTr7Hs3Phetvqhg7Kk6/U
jT0id219HrT3pX3h0EB8bvVyHLCwUyX3A1y87DroxNvt8ngEMJqkRmlZXT8ka5Yc5DAved38irTW
Q9uIqTgBi5DxKdXakkx72iim5kxbwc0won1Yo4gT6o5k0KxcgSEGuhiwQ8RjRsqZCNwFSmeGr5YF
kdy1MhEFGAyh+EVNUvwJfdne4ygv4RzvI7LZBnWZuuKrQ1uwhfJNiwti9+xIQSP77X7AbmbRXL1i
T5zR1H91Ohf/WxnDufONRfMgIDScEq74BmjKFCsWVQ5xKr8eAh/30km7z12H8LAo7leBbNeNmSnh
UHKGilwhXhqPgyY1ah12hEEV+A7zbJvABPHJZCYk9EwJ4od7RyVpfOK+QeugR5TCyXzHGdGW19w9
NoU4L+/03cxv75L8UTgmFt3KmGqjLOI6Bh8HAz5XW6RUA1UuqLCgULO1MEpTX6QoCFZvcRK2TB6Y
adUsLLYIjRTLxZxzVwwGxylIL2WAl2muexpFBo9uAKNyX7bnoF8dMxU8hSAaZ4tupcXY/RDwyJxg
HEILeaFJFEFqgR9I1emgY3dhqoORAHOrmpHd4rEBhZUOlmFOXPF6aMjIfn9+E53pQ3kkavZ9Rfv0
yZQrViDXk+f7fXz9X83t+S7KjbzSSMKL8QusWcFn/L7MyXpNqiA3xsIJ/hqueuZppDnDxxspQ+39
n5avRcGaakh1v6FD0GE1W4orUxcJANzX8c8RKOtHBGCQ0k6QYA29UMvphTIIdY7lYsLPPAgQ5GV2
gxiYjuInCEn9RjsgdKfXHQ80vow7byFwN4BGowf45R2cjwQEMHt3m8WSiyI6XKimTW9E1xTsyqOt
lO+e5JAEkCR2Dd8kZdngI7yjLKffDxlpqEid/wolXZQJh/pVvZNYb8612JTo7q0YXfmhJd6DR9S8
XERXm9YkBis09ndUm//HpKfD3rR403Dqb+AGH3js18sQcolNb9H4L9nt9q6oDNJH5Aj4WNA0Zfhp
v8poHwQdbY3rRYad2RS5qcrCyt7QOWocTZMIuy1yo45MEs1r63fXYwq1/3dW8IF95x5YGJoL2V9N
iOZTyIXBmtg2s3D7QHNl5on/Fu654lo6LDcO/CTHA75MpN84UMr5Sm8MfzbXJwb0J6clFPUXpnh2
md66tEzj4ojz2114/RPizLmIHyPqg1jB6YHbqmSaesCOST09i9ZYJFN6a0iiPrO17KjRo3fbSvx6
Zz+uUcifIaGCEzyx5EBLEVi5rDkHHxHg7Vm1FumAPmwZr1rPKy9IrFXiNg4M+bkj/wUhvk3EZlnc
VbU49tJpcioE0p73eBYg7ilTB7G8lkO0XoEtlJs3iw05OYbxl1VRe+wXVZSNtnoGtvSdv3lmWQSd
/rpS4MBeTt3xDpY/UPiIKo+8MsFcQRmLf2uYP6CEg3YX/Jjdh2q1BwzzdXnOBIeT7wmIODP/d6ja
T293iQvSK9L0mrQitM7PIVBEOwZvL6zPMBv2zped+J3BMR3LbvshOJgqJpLnM6vOnqYzKorJ7j4+
sshAAg4w2FzIrtx0m6R0UdoQNwamPHSD+XHWyeMmM3i784hD+Gbh3damVu3c705oOavK6AAOzSxV
6kNQN4Q/cUQdODm+WC6iALx4QqOKzATojQM/mlXjGcQglq/eGQyjU+nf3JCqo+Tb7+QPzHg/ul3O
kiHjoYXsgLgIO8lDsBgjMxgDS/FpAHYBMhJCE9EJkG8OFpy2lawBsePRxmUY3b8V9xB3M9ABWZRv
R5IHBhhOpmJI9Hlfi9rOo+plXyvlMnmDYdrPLrc1Z0VI6Y59XA6a2fZGlAxRe0APsaYonHlcp31Y
vpGSVrmBV7fFMmlGEQu3BX73jJ48yO3n260yLX2bz64LiTV6Ifq793LSpi81/7kTVLeEN94+cV9O
BVNBU3AqAbYfYOZngCO/sr+bQBXsFkMCmta+77XyX/rNnUgUNrkJayoIo30lDglf1eTPdqqr4Use
rm9yVL0dP7+jQ/ogokN7OgGkfsp+KuGDM5kxg+LwvUScXy0laKcLSpCKk5+6bEcMz975G3fYBDpa
wLT/a1fG7Rkc+kBRXbo5fKh6v0UfxeRRg1RZMXAQItjCQbfzVgzjWfHJzZRlDEL4oG5FpY1eII6I
DolDmFDVrvgWYkxEo8mrUC8vOOmnwpSjpQdtlv5pIGWv/foi7BZapNAozar0Ot2r13fDatU3/GAp
Xv0Quecnd4PDqqiV/7EpSpALpO0yVhGYwAFjvXzQG8BoPCqgBR/1LGqEcOcOuu+iZ659LDILNMN1
aTLgP6NLwY4SwhsFK2srWcyD+xeJSus1Vk6nJn3AtFgLBmPs580t0RLVK2PR9AqGQETiEWq/rXNl
j5LzdnNl9pQ38V7klBAAXC6UGnW70LqAFJi/1fVtnCJthGRWe2JFPiuyQEpYDqTtjUhLmqxg41OG
foTXc3yI+S/eBMf+VG9OicaWa8LvC8eEf6Gz+CRRV5OUwXCd66FH8sLWgqpQQT24HUs+0sz1v3HU
eURj/FZWinZy+4Up7yu9cfGIH6PKJBQcP/bJ8ZdJ4d431L4qfnPo0hGDsaBUhjkRe3Cpo05rk6x3
AFZkci3yrbUidb6HqS/T+nuV3gf845XyM+3p4K1e/iSMYDXDPYDtktb0woD4UvQ7ieor0j4q4yBS
jkG9kam/b6hYrbDmI+bV4Bo20eeT8FNS/kegLE+TNl+nZyC35Y9HkHumRmeMVqBGJIhJnRK38kKv
1VfoWBzeBl6IhsOAKrtLMyGSOd18CzRDEsGOBlWMLhPLRVQ7A0LtlQ9zy3yBhc1zqO+eFK4VOiGt
LL2C22OxlFh6WBx8LB1VE5tf6tjh/bjJm3yzEtj1L+8/R/vWgjOyfyV6KewQboZpWke4FF+Vut0W
GGI/xYxdFO5PcK3T5b7qRvopWndnavXhRRV28T+c7j/GXHsR00AuER9a3XShv16goezXB4iBnt8d
5vW/QQuOk+TWRviOYgqj71Wp+QRcPhIoBZLyGVxS4HBs4idVK9wFDbbhwgsrTJzR1qzs1xpw6Edd
EA2ZiRkVRJPsPYbQoEHw5YtyeqzsR3SBZP/yHHOKr3Gs5PpqLMFNbMe60I5kEXiFuYM8UpNk/W4g
mPSyR8TRhSQB4aP0X6KAUFBEHbUNZ2vAT2TWBZqoe/LnOeAiDONryAtr0IfOPvfgUQuNIO0wIfJj
qNXckIL+T8KG9Dpf2+wmiiByx0r8obyr0bzpBf6uG9VjEdcwAHfKEsziHg7y+OR9M1RsEzw0zQ5A
wUCFFtGA6bmE13JL4BcJb3sgjlPze+0Uqe2k5dZWwD/b8F654Kilnv3uc49BDgovOXvBUzl41i3W
fzZds1Wx7Uin3XKc2LO2H3cVuTvr/rp9H1ftPsVM+eEg4VLyxihsXLpZmucZqWKPWE1JwAXkEuxr
8TImQLpcPYGik8i7d6ulhkszqgDgIQcyYCn0IJ2CsBj61Sf68gwvdiQDec2851NSCWvaz6CNtUMr
OQkELCQosKT2R1WIr7zQ35BsvhLjZp/Q51VPOYQsUD0KZ7enc41Q59HBV4GFY+WTFC+kPqXtTPLB
MA98XHnRC2ro/BHfN3+1nqZffG3J6sS35VEuhoqNnIxAdNdhbROD5PzCWhBoHQipEeHrsyuCMPVM
hBXqTTcau/M9l4CEa6ZrcgkfORXHpEQOZffBGV78H16Z5VWMdMgmt1W9Zd+xCfg8B4VmnW6sMH3O
nLM2/R0eGeRFLJ48LoRR3GOt1PJ6fpkj/oQ4FuMvD1rTQQ85RiCvqs/oAEatfxhnfEBJ9+4/bigw
+jLRg/nY2AKglUt0NbSvpcL9uptmS0yaVd72DuICRo09CrI7aI3EtIth1FrdkCVEAHSqOyJ+qSaT
6cV1qns7p+msG524knbPXzw131X2eACiT9cXdYeZtKwmjTobj0mf7HM4a4wmAOO/Ts2kfERyx9o8
WHwX46JzgskhVhh32U6AV85mdTF2N9BQ1YBVp/qb5WfA8Hq2VV1N/8EixTaRfFS3cXjUEsXyPj9L
OQ/xmDJmsjJ8+VvFSxCbflD/hNImz2mOxtppVtjgiNA9e1ZOw/T8RInhL6Ahw5fHN/3bCxlJv1UB
+2u/lcMlroUiq2fgzkxE+o7OLab/MFNsz32IFwdchiDYC3TSUbF9H3zMa+kbV0tiDIzWZji6tjmy
FziZhPkB+Zp+CC1E85huTry66Fm0c0tfOwPlmaidnxIH04+EEgwWkIxU/L//KJ4TmngtrdSh3XPP
pyN4N4tPZYnyFlh10l1675LqMxzdPsu/ytGX3o8wypNUvTyA8aWcPUTlmvHyVAMO/ud/1kdYSegG
qWNBGb/6OBlM/fQIb9Dl/A34lSZn8g60B6/KZN5VmUWdfV6VXfRci8s7sZdfAozNR9kPzTJnaEhj
dQGkZB0/A1MOcIGsRuy7f6MM7pEVuWTGM59vaN0OmA0tSf5FVCxZXhF3QTbqTwYhCY+zQacqtvdM
glvMgOdozWOxralPROWOp6mD4MzAgX0XoaU2nATUTSQc2pXvKEJj1wwdjlsRHNzsIwjlibUjffkB
UT1PimzH1n88hW+RARuVDpQ8mGKzkdz6qyoDTYvSz/OCISvDWMuh6KvFR64BI7M/mPgKGXoqpEXx
CPk4CIjGTglDUqA41FV6+fPWxr4gvmlasq0NO7zFYxJUGr2GaFWEUaePBdaEHN3NDgNncDlmBgpV
sGa04vvgOUEbIN5YRecAEbOri6P2MLtk2hNYDTVk4nWM03GqhFPHbn9apGFM4ynJQ98jpHjf1rdm
bE9NHo6SnSl/VQbmkyTLkCx2wYYeTU6mJC6ECUwF0oRdtQr7n6YOl17E5KqwbS4vpMVnsJkkSxDD
5NfGju8fc7BB9BjWi/rR29i3y3z43U4M6SVjKWcsBZe4NMnVNplgdjOVxI7fN4QXtbzH5IJpfV0k
xmHS+EF6h2iYiKlsT9xIh8jpZipCohVhT7fXV0wb0ttaLVdnWyd37Yq935PS/s5FHRTKd+yO0zr1
r23SizJDqHu/AEA8TonRi1btrVrPO/Q/HSCVPcucJYLQkd1UK1Rx7NP+chBl46EdctaHkQIbCQ1c
ubvuxR3hMejQcYvC74s1aRj0pB5abNJVOWj/hwZYyz9dENTwByNz9DkcwtkCGmHxF/INCfqBnoqt
WCp3eziQb9/66Trk0njjCb+2WLTJx4ht+CBM41GuwvD74S7osn8zp8DLMWQrBmBLstWCRs/gdCZE
Qb2wkeDEgwq21S5p6sZ4GjxRDKg3toGIDIGtCYXezSfXZ5IkVnZLpooSBqowFLePYZpT4MavlVl4
NA5pWurakrfHaI1qre64pgS6ZXbkSbZzH/8m2P2nna5Ymu8K6VUF6ChsnZYDdbHUpRy8CU7OMMii
jXHh/hj2mkMz4XEW9zR241QQnF8Yx5qLZycvJgLcbZWH/wTmZBqTh2WXfz5BscYDVsu+Epg+o2ak
fdEEAJUFefmE/dfcMYr2mMYse4QnpyjWKnbDgkAS0v//khAd/ogZ9l58b8Iif0dbruj4A7klwbO7
QkpdSPtUF0w6kpLzgKGtWyIuGat+AY/j25NIXsNVFhs9Sub6UlkDhUkTGqPcmLi+l8Tj1itzbbBM
5BXwNw88QD8kiqIkZbk+VrisftAy2+8Hkdq7nLS+e/FpZpag4vETM/Idx5wvnGtGdw735NyVlbWH
C+KzK+Ff0p13YhgnVRN1gIvNQScl7NdpxszC5s9dwM1SZ5/7FsmIgvCz8vIZsjsQhskCIWTJytyV
Yk2rA0UHcJY5pFf0tYOdAjfYXXifozDOWidJ4CtztFADluVYY+Od64+44DDUlPeyvEKBk7+iTmXs
xiA0f4ORtQQ191SUSHdeqW1NIs/I3qhbG0u4i0YZTbDPNMle3aP3sjnYyiX1EN5nnttZblSlyId6
FbF7ui66G5xVfEwneh9lZag+my3Jyfsx1JH25wGDyuxKl37ASQBquobeCYTPHHV68Ofra78mawY7
Dr9Ixt2DjA5OrxVcxrn6Iu1N5KMKbR44Nexj1XcWJQ/DhfnASkjedzbevwER7zw91tq9Sq6aGZfl
xHfdkDBE3Nj+tgjrftG8ExeVaZ/lT3Z7Ve6Pd3LmihOIUfxcLMQGNsMsJsxKna7kznLeNgp5peLw
87migtbzIp9ryL367II1Q75ImWV8DGGe8ijKCm48Wm6ORq4+aL+tvFTEELfq6fJGRmHNd788+41P
YTk6t6RD/ssk4Hjxoq1dHxulssS2WlxDD75j3pPfvYa4kExgiEWQa8JdvrjtLW+r0Tz23dBHuqn1
hH1gZ46OhKoCcwwigSVwPrvgMyusZFAFav2vKcbPrYlnyGuz0Jk55bYxd4IG9Uyb+e0Hgf1Uw1NQ
Rbx4zTLwH8bDgx60hnPeAogeb9zMB6x9xKZQES2WSXTiYFJIWIXqv8dRsWS7x0EyIPWbu+RZ7E6Z
NgrcLstS4kXGOQYqYe8xBHitJBhfRixn8Pq3Jee7DgzbaBh15m+Ru9IN62Mu26cRz5vnrvKrBcz6
r1PJCyAbwptdJtawc8eIrH0egoYNmzU5D4tag4STzBqMstGc5F9IobzCtZXKc4GgcffsYIo/jiGc
Zlgq5yiQDBKRx86rqzYEPCqv45KmoII7t7pK9inKpLNz/OzzushL9KM6bDL7WqbiVp4GtanVVtIe
AUSQEn+PvyS0PkBrC0gw7ya9p2TO4Aaz4P69HQDTUw8RpUhRwD6AkDViPo6g0A6ZPjKUIMXczfCj
IsaNctQOd6e5Zu9nECOQAmosptNaQKXps2ylMjCO7Vpoet50HpMEk09ZZB55yHFJi2+/kweWGJSw
6ZQGEluBxt5evtNGNLZ5Nkal2wqTJjUyPWcAlnj45eKKrjLXmZmq8/G8g9ePCezmLMH4k18lzGJg
tmgbixU3/+luyFwfVm01O4ZkQb8mb+KL8M1xGh/5ixm3TpqDKNHdMRKfVsa2Gfn8FN8g53ZvJD67
aUwMHfKLs02RMXuqqKqvqtmL6+PHAeuEPWefaRX3iCSCj1i2uYpsHA3Qf17og9QcgDgz2MzFh1Nq
/alcSDuMM9alqdrPhP8/vVnPs5/+HJiTfG/0E1+b0SzE+5N4qXhkHQuuIJIpRk+6otxsi++1nGfp
SUBZd2Hf/dt2rwfQHTDhnQdmCHUpMFLnEfKwyP5WT/tjRc8eTEuvs1y8iIpH8kLS8hPkV4ItxmaF
fhnvReqbgw0UW0AAJtG1FXuN9nPbhVjFZH4ZR0pMRtjDJOSo0lblQOhIzmJf/g6bXNYIbmDjVT3k
TCdNU+BTOCeONafm+OMGhneR15G+ifD8zPsvnryghSm9VbEofrkrG6zaSGjN5wW/q9LvFoiNL82i
Xdvmc9l/uNPnl7z6g3XpF+neqpF7qxv6UtwZ726Vw1mJzUGwwNqj4Jit4oM4cq1QCu0O6Luv+5LD
1Bfm7wY5UOlruoYopOUCp2oUfzMhwUFPYnFiPrnI8z28ZLfaaTYqQUtb+kFr2mnbpEOHbrKRbklw
76E13CgwCSSKFUc4DgQLrUb8Z1XauH24Cq3c63DKnOFoGUZybnFEX4vftkcBE9ffr+jDIoEYPw+f
G6oUsKbnB/mUgejv8Hv2erBPUNHVLeS6xbsrkiPyw5U67hSKIiTfOPFwPo9WCBaG/rslw8EzdpNu
jV4dZEpyFQPnZzbjZ1895hYLK3ylqkrNv0tRS4I7/vQ5FtCoFme3deLxF71wAl0Umhi2J/Q+etFm
lTYXo4Vr5VEfH1kEBWJwhSsImi/7vBLGUjCfoJcg2HWr19fhBfpOtMJPtXzueESUUucBi4tzX+JU
Ocm7SSNMNxvHvUZQbx5AGp6+Q9ffvXkmEhRbZjmx6ego9OW4Ltp5nUIQWT0tPOdx1c7bg2+82ewZ
oEhIiyuf6dJvWPbQBu1RXnTztzoRuyW1OlAdkrho1kBZrDKBD7tQXxGmZsUAAL5BFAjHxo6R6adx
asSpXVq0bC3JtZpgpq0nZ4WaFx3xNEPFmifIYRarf99rq4n33GxOn4lw73TFhd3w0Rr8YCGybF4U
3ANdsJMHmpIB0Ht6phSE5xCcE+h+CWQaPgDkK/hLde4T7kccVUieeyplpJ+s5nFrJR12VbuZvEvC
SgmnesjmjTInZ9qAyhhuVfelS2TKeijvtHvJ9VjjfmvQpZmRjznjFCXYQ5/U0LaLZGMJ8f40uOoE
t7ots9IrOcG7F2o9SFIc0tYEGgjmcyKeMnVjq1zaTyiXQyYNqu08n4Iou6eIbnYghqliS3soc4NP
pS0B6aUxZiHPThwHluj3CLhCjOvDhRVESOjnNxNhI9mrweugsxfj/hqvX7KPLuRcpA5/C7Y72z8+
KnjcWA0zGxkC1PHPH2WG6gymgIAIetPERDXS5SpPORfR2yoOwCAIlNzzSMQzIMmP0ZpPWRxDfRrJ
p64EpRfxumMlQb8s6Rb9kzxmUEv5X8/Gag/Mn78mg+043FEjvSE5OHphmv6uzoroJlLP8MDXDPQu
mkWogWe9AbusrZEfC1K/F0hIAdJexW2HRecFSyhM7/mWyg0xAzvpz2EApFigYB8TeZ1xeuYw7H3l
JMLdQBPodPcwxmfxjylmZ7kLdVKHBsBJFPdKsFUE3tanV3uPJi/tj+5j2dxXjtCYN4APowTDvo+r
RZdntaAdrr8rm2whmmQuWuBmNoAzqCECCceEKp/q2eEIuvx4ertCSSDo8Lb1BvpX+Wat8mt1MWNY
/YuL/HXinq+1GweDaKpGtC8iWoTd3VFM4wmg1j3oeuRYlLA/C79dgemRH+UOqYg0YqGkim4UJ2dg
jiHkunXd34s5O49MK5M2sRx75VORlpNCFn0dTDD7meSAIwxw80u1OtF4a508Z4RV9jNVk7Z9GANg
sxC3Oi5uga8BErnNkJMrZYhVCoJgZH872mt44X+aBk6cTd4PZi9vMmFpDk1iTsP4NnMkZQY4+Xi8
xLBBzV/LqUfrZ3cmsQlODSUFdVwiXRHR90k/X+FGxET7EhGoT+i8k8eWdcmjeHLEjPhCySt9uaNu
Ki1qcSq6koRUec8wyRCeO47wVznmv/wrTUxAAFnyfe218emvSPkXdEHY4FYETgPX/ypxMQOjsTkZ
iZUqHY3tS4N/coJktW4dFl5MTbGWTzufAzjesG+Uf/NoDyhKzyfISDyZ0U7slSV8CmrOxc7ixO2n
BXidMd+7tfTp9ClBlqGH5m6N6DLx8Ov5I6NBeOZRBYujtEXQ86P47SvGgZdFGIh0qcDqRwJNz7N7
WaMXOvkyGvHCyXFt9QJvU6+a8tWWX69ke0StX83jAQUhK0b76yCe6QjX3gJAwkNA+nUhS5xcjszJ
hm/N7nbBUOiL0FcdxSkIvQityVco1AMkiALPLdLWV+eA5/j+b0qWvKxWrSuhwXXhEs4kcuSOdfmT
FcubvVi/VTvvmkg8UWxRKFfxntii8n1pK+QeNEtbNPmX2zIKMaM+3A6mYTSNlxaQIrIrraK+ILyu
UxJs+AeT+yFI0uiRbUoovmMGozo9EpE3QqWAmlie2Saw7/hTlI5KtF55qIigvLMCpy7FiHg4ubEf
QjpjKM5Pk+NAJq5YVEFF4gpkP9U45UZvx9XMKtIIpBNwjay8IfmI6drLjewcjj8PPP+EUbFgHrsO
UyPMTEJpKeQD+VVow/nOkMp1qNwHC1/wn3FK/57XL8sEer44VNRU1UH2rZtCvPkqdVnTV6n7D1dq
KCnYicpZvPOz8z4BXW8WLhKV2AVEsrVxjezIG3momuklWIcDQHOa8ucDztQLrpqggHZ8tF4ZV8IE
P1g2hYN2kx7oHqEKc/4B4iE5Z/L2m6GxgNn6L3HdbDbSwPfTyApm4hFDWK/0LHTHdlMK5yXfoYT9
zlUab7kqfsgDplmEGCWp8wcodi8V56wKremgQ976xzcdNM0h+ICyhD85qaVicF6hTIG3Cu11wxYW
zxsi9YuOkfWAQhDeU9mfQqIF/QOrKKYhCybB8GXw4BspUJj/Kf1tQl6nXtaanbzhLVpzx5Mo6rHp
I834tsKJyHdkg0ORGtOJ9+71RpPrZ7leA7b6DLRG0DfGmo0kCkl82zUgqlBamYawtZprOAzKVXNM
BTUbXgimwULc401Lo0IHA1ilrZ0BdQilvkanFuvI/AKRNINMGryzA7j2Ibg7VzpJFZqtKSQ1SBav
ld6JEn5M/xqnHARORB6prp6gsvRmX8RtQcBm2ZfebnKhgCLeEk4Z7Xus7yN8SSDiYdzbPA73GyMT
8dwZLZ317mHCTknXci/iRzLPYAET9AZ0MGnj6+h0jbccPfQKytlZqtpyHp7QCmPh/ZMWJ7PWyuQR
1uBgCBadAVBqyzWEugkx2GnCq6IisbA69hi9HdwT6PLpaCbsgV9ygAiZ8DkbNTbCAtZgjNz6hx5b
P/BmdRLz20lYUs2yCyK7f8ueQW1ffX2tZpyP3R/v0UeVT+HE5PNjFCKT1WtZOMrwleJl2noUucJl
g5cv/WghCWbtNhagC06R4/SD6kJxG9lVittkoEMmWivGanP6SWwcMpeV7A/nPUyEhUHVEj6+M+hY
YV8kPQe7hEjHFMpqUyk4dAcuMl0it8/PlXtN/F8T7GoGiHpXyNaSBkW+Uq0MduNLlnpaH67sz6CI
UPMuaErkFOQh1sde2XSU0gRjnG/d4IOzwpvtGbR0vLPJ/KHAaskDkLmN5QBeJiauDIJ62q6LKtiw
BFpo1qEyBxEgNOQqfjPQLTaCbrOGVo9051gbvyxPzp1mY1r7cw1E/iixUbDbsHP3wz5OGt+nmsm8
YXnlrg2MusxiHPsYDb35AOtw/8SHX3HBJKkqHnM74ZFq/Alnln3z4v5izm+bEPFfCNDJJgicspW7
18pZ95v9sn6dE/MNC43A3PmkmIJnsn+r3h5aAXHNFOlhGqV+MUSEm77V2qecD67g/R2/Pg4ngmb2
viTiog1TDARs8iDhb7sb3Tdq8jqjjlDs7sh7mbraZ2016Ex9h6gPRbuHtPorz3Agy/lcS+jvMLTa
aajpuAkdQ278LtPwLLY3QragxkVKFjjM3fEYjSF3t3H1iItb93j5LWqJdH04kSkI2nn6wByu0tY+
h9fiCvW6AgE5TCVMUOMFsF7Gq5Fg1K01J50GQX8Uf8a8onEU02QuS6N/shThF1CXtoLcSi4tFubD
cIKnVpsflivzGUpNiUGa7OwTZf3eUwPWNTOwbf0+YsFwlBUTzzhHOKmxMqYc/ajdXoYfA9MQJfVo
1KzMzNVR54pUtZxYp5kNRM2ZodsV3PtEkoJZsn7o4Pb5OGFcDSc/jUawEQMnQLioMZRJUaI2itFj
+6LV05pZJCqt33FNxCCsxcp2RZpp/BB/msBL1j0ZgTg9gOH9W8aqSdMBDbgO1CgA0GoMtlPRe6wL
qUkUqrJgtRbWLMrcNCpgdpAoynwX7hUsbpOFska7aBlRlkx+Ct/M1xOJhebh4T1XLcZf8PDRcvHg
m6xNoaBHXEbPfsuvHMX/THf+4/fYOoCnUlT9tpP1sao/fLk1Wj2VMJOreq7/GY4urTqHwlQbalGa
P8x3Pr///X8bzJkU3FF6hnyhQ5mLIyJ8TPC1irA3faxJmYLaQCACh5jF9wI8ZZyBL7OqmD4rqRyc
DastQJCj65q9QHCbrMVKn2m8FdboMum0qbxVPuLB+tlz5UXfmCt6rLaJX2Mx4eoUSBSXYmzusJUo
YqfCUIkYnheVe2eztUg6XTdbDeQrpem+tfGFGZt/wKM3AdpHbdwoPgLQRZSJfOrs07XKcsA7J9ww
8sD4SkmsOBlmsse/gpkdprD7H5Q3bkqq86cVg7FTWBWXzAKV+f7sTNlzBmQVJJpE6h+3KpKpqNzo
DZsDaJKBHSxjrUpX9OfHNyg0c9L9QLlR4tvUngAFlCJhmPz5hZtzw2UI+Buv3Vol6xOjrVhWcyz9
x3rwUWyegd/Ef1qVKdQVvA5Lk9+q4G6zfpEmlEIFsXdkWWrKG7GNp0HKFR0phrjyZfGZsKqC3kui
DQLj+p4NKgqcjv2gI3980rw3n/PxD3BFzm1yurtXJ2rA9wr3wnFEjdeKmZ3wDzOJFq5odQj6i/j9
gY47ilCZpvVzb7SqJ7be4iXX7Kp1K0vTM1ZrdDoKjZ9EabFFbaLBAc5e5GyH3iSmM65/4r1sihXM
cI2RQsVFpbJ74Cy3EGjxb+BO8qVuxQTdurugSZm3RwVrpCw9x3SFVJqZiXJSq3OYFXJTNWNv6KGv
tke6Y1Jx+zFapkMvm3Qw+eN+zMS7l7ob4cLQX75LukH2MN9QGY0kpayl+IlW68qAVOPYV0QqCAd3
wUXKLUZ0vhW4GOVoKjVSbxWOh1R66U5YAZLlsBqNpIOqNSnno69chDpCxOfnEs+dXbaWzhZMXC+7
28dQXbnn8RCTF3OKRmQiIkVT5lF+5YnhE/OmbtqIvv62psmkihsAyspQh/SNezRGXVVjmb5ZYajg
KpH1SYGwl0zbYDNNVoQ8M6UtWviO7aHy/OiHnUCNYZsdrGkF/0U0Ha43qOSCURfVPLUrb+JYpKyA
ROycPuk/AuouTccJw/f2Fv16H0DUTeNADJx6mwlq4HVfBAsYinayEZ6J+giacuHaqPBzyGqSMKoU
OYBV8jCEe2mWuBDK0h5DDWO9m8diyNyL70lpHo342fZ1xTO3WGeWL5oQOTyHFDKF2Dqig8QDc0NM
ZHaf0X3Jtlnk8yZarhUqDwpkvyNEv1KMbUooWqo1OoofFTcWK6yuYfw31fEDnrHQ1PoUTYaYVcQ2
mpoeo24TV8DS/sZZtaDMX4Xm4pDlaLcSka33McfX0X3nuPDzZwnhGzmYlanWlQFJ2UNlM5WRApv3
xNSxzvC2XCeYtp3wOyJDNIfLAqAunsfuYUgHZsuwUn11aQdldFdHllA05YXrjjMOxjtG3Ige5DuQ
mLMBHJhaCAisM8f+vuSJHVj44F3c4pWb3GSuYBgFcTWachrQGtVa0RHlJmkmjGVJ/mI2yjhCbPcG
dz0rJv9WX8BNN8GKHe7ZIht7WjkTfvFx/6sWnCSfm0CsF+d9143bQdJ0TabABqstbi/tfjWT0RMT
QGUiZzPD+kIao2KEH4VQh8/d2DQx4Utjnj5wrh0gyoEhlyCs+aeBBMvKWepke5osX4cJ9fX9y5YL
8GHUl1iA6qyqxgGvsTy20QNRgq81n9rPVZYlGinA9vFQDtUucBQlPcijUtWQ5GeSu37HNFBVwGmu
Fc6degUuw3Uqm8mFkziJfFsivu2hDX400CyAZ3/RkaswoDdTKXR8UAb3WWPYltcuNi+tPIBP3XZU
XWQ5i0WLBv/He11CpSI0v8X4nzffo+M2J5iiywsLD6aIa+H0SHQsQzbuBhhCgXU0PtsJsKY4wV9O
sVlYRi1zrvlbgpCwTHjiJu+Hst3wsjDqOaZdvYtYtHF6nMASaAIbpUhBfA1Te2brTKWLWaz0Qua1
aDoCz1KKDU8h+i4XoNKzKt0WkrZZIvwHgYDtmYeWcX+esLzZb8r43nmdnrWYVp9ZNwcglMFOOyyT
+KONiF0DSBcXFj9ttqdHcN4oFf//yLYB9XjK/rllRwyMFfkGFrX/V4oqgvQdj5f0y4/SBgznDroO
t6IXn+qUvmdKc0u1MqHwob7pGmE/Fp061upW8Xc9ali8s8nmOZJbZjOiZUh4mK/vYqOaWBgFR7a0
Rj3kQqPhZH1C+/jldpH7B6Q/koR1+qqu4gDwp+uFwE++U+oh1JwlSMm+L1N+VcgwEMou/7kCnrmE
wwDM45DPGSFtKWxuPOrUsyWHoBwv1+meffVG8lyoK/fMhP1UhezFrKz0cfUlssGQClyCpLq2gjZO
nacYtsSKioz3HcubH7BBagH5FrcTqQlvbbvibalQ80kgbYGzReNc+v5UaRLnTo5s5Q6/Xlg9oDBU
BL2GkMs+USakgRbyhcBD805T2jd61tTjpweFx/6y7gOcClweHYD+In27bPD+PkJoOqmTfA3AQfO7
BcaJV56FrM321l+UAFkXuTBXgo4IrNtj6isMeddqmp+njMsAHupAGdR06CTZ8noFWWdmmGhqNVLC
i0PUh32VTEGTdg5Poh5zWDpV/6NZg6euP6UDjArzKIijmQmG5Gze0pXBhV340DJ9CagKpi+KDT1q
iI9bVA+/FKJxJVIkh25yxx0m5UyDPDOplzRt9qVpmbFBL9hfk3dehcLt5rJgsvoXSLZuT3DmEZCt
iRLLjQhC0XnBa4L2IvLZrJjNooMjxF68nQ8f4Ueu+tPiK0IwG0gcnn4ncpo4g5sQhoTH/EYMWwAE
y+Jl3Lo5djkSFjIrbt3YGq/7t4PVV2XGHwFiuAqedvgFQDYUNZ+TMXIhStkr0is1dn0lk/bWVVYF
pgC96B/BNT/RuUrZFCwG0lJgs1iylL3ZdgGGgU01xIw1ORJvi36yQRxMnZEi0EOovnfDd5rz8Uqs
8t3AEFesRwu2eTysgVW7JtTeWBcOKlMo3jsFEDR2NYmMnF7rFzepJnAdw6Ysc/iCICiCxvzJNpCG
3hayNpP/hOGfrqHWiYt0hqNkFzzwzpqWEly3rnc70NI1P4K34vD4Wc0ZOxO2w48cEu0r02r88S4S
yZsYK/CoffexFXn41iOu4ziXjzwTI2qFaTGS8C8y8ucRVF4ma7miMYUPsde5A7gSp3tlNnscgv0C
/xlgNHC4Zfx6vzsC2oZlxykA6hYz+IZZpTCsV3KeOqp2PcCMeJ/SUxyg4YwgerVZ2M0Omhs5rsS4
m5xBa6ly/P9Yswv7GrOKcTIFUa0OrDADJKXSYCZcHM6rimxrKAMhTms7SPZeIO0HuxveGUX6eIvd
iz4Kn5HE9xcJ+169sc1bRh4UcmgsgOcnAMGDn58kTJCpkkWAAos1vc3Oayo+pCF9zL7VjvKyPmZ0
9bARfXc44uKbcO4OGNiQCXDUzAB0eWySzKyLd7QjcpWlf+rne1nYFL2L1nbOg4YDygBTh307rgKn
ickWFfJN/ZbwuEEDwYrSuJ3HKGgwUsJ7oHpzGJAqndW/1UNhp3+1NKa84vZk4pWbY9rf9asfarJQ
N2Nk8ZBlMul5GnG6C5U7c3y6rNzD0kpQDmFp99F5uhSo9CzaPpvsitjsJih4PQeEZUxAEW2Z4sqs
y3NHgg92IARqDxycTPLXLPn7MEaZlqWwTYsSTkShCnMPp2c8mb6fU+7/FweqWQA1C5qYytVV9Ckh
4tnJOUbKmid7ZyNHSrwALcnRA3kel9rLAFs7F1NNEw9B4LPEmMmIftoz1WUC/g+hbbUBNLVEGLpu
p+EM9UZocHfceyFrlyE0kf4UbqC/xf2C8JJnDzXyHyMti1rGHbigbMIT1TZvsNaChMW6Wbz+06xU
x9F8DGm90LGaAB/qRJbE6lqQB0vFKVXxnrZok3IpWkj8zk2GYleBiQOh22sksjm4IT5+2A2YkQrc
CINzzvAuupLQ/z2U+kaR8Q1/1egGs/Jx5nwKKgqBH2MFUCwm3otOTYmkcbA+S5KBpB5OE7v8GxJk
s2uNQoZhXivKsDvFzNsThJVukX4aC97rjizzMMMB7eD9PkGD3bxKguiXEduIzmIYNdp8jDdt7OPj
p6jA5/8GmFLjNaLprOeQNGHV0iKkwd5GtW86rUiaBFedZv6MBee4EPOB7ZjPaymabVSr91+oI2gQ
xamJSThVdtU1X2gJpcYB0mNYopOGx39hnagftgmVMIiHozu0kFSSQSsoWpAIi4RuYvxz8iRDijVc
sGDKlSfdvUIWmyO/84t89toSqwIeHpfpPOx17XV30V91bsRwnEywJqQGI2yQqoyqJ36LcEoUXKyH
lj1n3ggOocH0QfgkFk3dga59YONM816tfDyRlE1HJNanrGGtVqd51TkwnM2rzbUtqk87fKXEOODR
h9tHws7Dad4+o4L+Gel/mAbVCJk8xMtUhdkuKDLqS2waxJri2O7ykRt5PAYUS7dZ1xS12WbjUmd9
650E2Ld8MEcFly8R6Wk3whoWVOTpPX0pAkAJpyuhSPgkrEqJWQ04fnhCnu0G6hsj1Z2ilCrT5P0W
1dk3D83SxV2Q1xOQ30xfbCSlO+KDLHKMfFo1HjuMi/HjFelbIN5t3+9gweo6sEZugIWTHBOn7/Bn
qzoVe86C5faZ8SfSV8UvsdsIj7T4gJPCBZAf86gH+FPnrcKUi5YS+7/dk1h/hUG9NUmxqfUsL+XC
GPhi629XyxF88bEAuH2w71h0aNiL/mBgT8L9JX9z3atoNXVYVFkIakI5jPAKcksHqsKyGNk7Uyg2
b5qwV8qCdSRfnuItLiWkB5WFP22CrfxaBf5H1Fh42ueBx4ZKwyACD29BZ+cFXzaRVLWCB4nb5tEY
Hix08VkF6DBGFMYzhlUunSSRXJSoOmb1BHKOgsEpxchH2shOD/DP8iR1l6ezUWAFL0r2y5O7S4AQ
4IwBVJ/F9vXqXO0L9lZDYPZhod2cWbcCPregQ/mUOW2/hqzjP9rTtPIbuzY7wl0U1yoSGvUhh1xT
2UnwXA4wuyDzqcyQujz9JQrTQ07j9O5XNKGv0uTBLgMTf8sKk+gu8B7qSZLxGA3z5FM47LWR1S90
nxSJ5kw1ScGvYZe+GtKDQN/x8I+uc73BN0kCVndgriV744XSTA/n0wRmub40foYSQXXKffrY/LYL
nGc0Xoq+PqftAXpt7f1yp1bUhSm+Ob4iC2qXCcD0O52zNfWITzWVprRjfRgo1NZG2VB5jP4TfGFE
2TuXLTq6Wmswef9gdpCUOalw4tYID0m3tSSEZ9SpOrYwFRYX6V+A4g7M28iDIDV4WSRp0V70AfoA
/9f18y2KhAi3BMGh4xAWDgJ1xxtgTy93XeMOSTjMjyFLnwZ6VPugTLS+/RTqyEDfHOdzXSwnskES
J6LhXCQOyeFIeEZ9AS4P408WaUN1wAANRowazuw5cv/dwyuXK91SeCY+sqxr7jhzxSjhKdqK31Uz
583kkl+57UcgAQYxgi20/ywyxtkmZ+PGjD/XJkRT9R6R5RC6WDsIY4ytI0wdInku2KYd+iMdc2MT
oFSZz7GRB+58LiVaWTeDQlqp5C2IEcJv/uYE8jms7rWZ5MNRm8bn4jvPmM0LQJI4foBo4DIKX0vh
N3DKFImB7WO51kZCa/xA1ZRMrBwQOVFCdRxNBtgrzRolQi1smptDEUACIufbP7DzaehQnl3Hiwol
ZXPwgTTUVFeg/UpDmM00P94743eiHchz/Vktn98QmotrUpz7p2aziUu4IpEnGAhkzY3UquNR9nuT
chDHAHgq3/0aSXTtPTPDQhrQb3+3yfYAnn0/nNKNR8rgYa2zxcYh2F18pihMeT5UYxECApITi0ST
hrQbVdzGpoT2Cqi/pdUYMhPCb6BVrnfuk7eOgNYW4pvxfxBkMYZrUK5xyZD6MIVsX1hpg78nGzab
uwLUugev7rCChPpbBCuBfwpAdeTrVI0h3uyiKW/Nlywu8M5TjBxamAR/+XrL5PfW1oCK0pz3yE37
hTudzHz0AbD+DoPaBmV7iwgS7CkgNnQoBuNubzlVyPLYMa3JJxk+IXQqxHy77IoOZq3l52R35Q5p
+L6HF3VXVZdzgSMjFqPLLSIgKms2LORvBnGyw68dRQcc5YRaeUhfi5eo1Za0EUNC8X/gVALhHZSy
u8tAa+wpMXusstm31016VlQ/mwV68HGZ8yyLpLE6X6e9PpLonQtoIUGEC9tyO6F4An/WS6pqYue6
yeDVBKLepOCJGMED5dVJASO5AkIy1G1w0OKa1owzQsFnVpCRt/w+BRqNu9gJ94xYt2wxSF7znff2
jAcAmByHZGTYhM6QRqExfCXdyL5qPj88xTn0ALnkx9mBNWMjiWqqyX3a22xAP2uMN5+T/NDr3foH
ewr+Q/KFat7hW1ZESFpocHaJzuG1+LUAX2E72jysqwi2UIydlKXl13MThaCI5/Hg1QeayKht80kS
YKB+qGYBpzUXs4nArDFDza7Hr1zQeq8Vge2zw5CuN4ln4QP2HRz3EhJo2IOZyVVsE/W4k0OunD9h
6QW5hywGbRUR87RnbEhyPXyN/ubJcnCuBqJkF1qTh/HJB8nhzc5kqVpmBcPYcDuQ7KXNUhCPexdx
G5rII1TX1YT1md+yY/3NVaUYgytnuUlDEENlTfQZXT2kr9+n6+Q0PA19n3YOQ3PB2A4jlu7wFfrS
N2FZNOInLIaW19Ddf7I3cF4X9XGbtIjDHsoVswaOXGRO+ST+vHw++qycCVZlD9/vBlUIk6IYsPFc
bpj9JijAeT8scToBJWU5iofjaMdYSXS3gDz2n/rYQyZe+t6yzcru8AVloFOjU38vcTGIRFZjz4Vg
zhGf8+vY/JL/sQUV5pLC82eSdoSY5n21xyOZhw7UBnVhXV59weq9qnOf5NYeZ5neiX4ZAdzT3y+6
WH2EnEguASCmwVdnj3feHpdzunlaJYuwBN7s/Z2mZJUAq8L6rcRH8MMNZ93NoRAOpWTyGUax60ye
J3o+w4lpALVicPNAZrmPtcRqAzpkufW0xGKQB7FH0hxsWxvmMAz3MAwgXJV08+dyBqkdDGjVioTb
0HE811pkQ1VYwTrXQaTWugY8g0S4TwpLXZD1ExxEwj3485xBkskxNBS6Rwy1XAsserxGY1uSVtSm
o4FTwUh5rM35mlKkZKr7ddZApmOzoeUrYDdFUsgYRvqJXMx8M591mZR0NWDbjBUQjGghThCYuz2i
iL+xsaRNXbIgY4xLFjDJJI6l5+7QTcPdccq+bzwP86ocSt6YC47/hED3lEWicx46Eoj8AWjhl5d5
kxdz69QSKB2PLkbEsuVSBVC+8mRDMHwoEDZm2APQSpOR+amkeCUI9Hr3ncUt3K/oz2Kivj6U2RZh
IJvMa+e8+sCPTUju5WjXdmIeejceeu/iCcckr4KXbHwWWoM/Ow3smzJbP54CligyQF9cbqI68NeW
i4RdWsrdtjeTKqa4MCVplJiaa2Jvcne40b08zo9+6kPC1sW/YyX6MbdvGq3TOWsxhJg+CV9mOwpT
idHxOmToDxFh4hSCDKIr85DaY9pSGPGl71prXBbR6vkLuBazgy1FI/w55BOmd1xAwpcJEaqfb2O/
RMpVzGXwk6qbOiqYWe3miHlOrbEvW4kvV4sfCtwqetrQ6VTKkcrdHH7Ta6wR+cMBn/2el91qP6jM
m5ZleJFia6ByVYrMQqQXmrjE0ySIDzxWuB6yk10L8baZAndgYq4EQrx/1ORYce9uQ6BFM7wCyItR
nuOd3i1yZ4tLuhi27Ef/TMC1hwtWXvBos/bUqJUxICBeQhItCuP7pcyYFG5um7/0/M359FM+InMV
i3geCftjk/cX8VGo8RU55WXZ/VXYx0PKOoOEsERwjwAAZJ3cJPLtjnxbNvkx2CFbgQKvo6DBkU5f
pePLHQfzPtZl0QzH4vxF1MlWFcZqsCX1YNSVqHP7USXCV4e2jOAKvC/oicL8mTZGE5LTFh9yOTwl
G9y3otmxvQlnsE2hGaFjL1RouOAaUGRKzIs6A5VhqqTf4J8t/VkDUJIBmDfkaa0kRa+yky3fBa/e
gI2ZR81G1beNnSns8g1XcjXz/OP+0cUjPqMHezuin0Dmmi1HzvoDaeAEgvSX6mNdf+iAfpcJNsqc
b1IsRXRDViLWDP0eil3A+N9jFnX67bcOBThhYNv5MNoEKpkVwYHEJJ+6JxiCmUBnbGpve0BN/Do1
QlbojQQ60RJza10+dNXcIVOPbXfRrCXUYYO3Rc0BiLg/0yJx1rjugOn9ZwPOHz3TQPY9pVkoSmFW
KxKjgEvnuekbdz3fZny6du5wDfxxq8UyUH3n64eDSJ7yE4A+AiPJ533brQjZrHFwvh/+Qdu8oYlg
RfvBdssN3DJm11wYfAXQro2Vg51IYhQxSjgtA/woJLherSRhw6pX2ut7uSN3uvoMaAk7cMuiPKHS
oAEyw2VeIKvG5AmO7+CgY4zfqFMWWsqzS6yhhacMBkBBIzLmODxdktdyl/5XFz6Oo6QooGUZsv1R
PXFqEwVDJYZYJElnaIsAMJ4/s2kNi6jL0k+BVCRh4S8qpfiidqe/50jgu3kcdFfKli/qoe9Y4ppa
ElZIgvKLyfQ/G1BvKpVMCuf/Pgy8Y0LImhoC4HPNVTRJS9/lX/HJbQ3t2lSnyPad2dMq37iVtouN
qLBcNK+Z4hqT5qwuPKwQdZ1eh7Hq2zX7JM19N2+6T5epplf97Ni7gBp42bKBkRlAHU5GoV1J9tmW
bAPUI/9GAW+8gN+0eHFVO0v2Xn22ww1NmiGJFBxu9fmvsYsWU1h3nP/861LQARbsZdP4m6GZ7iyD
pdFs8pzwR17pnzZHmrYXpbTtWMCDYklnr76ftW+2xSQkh0Mu42xGyg/2gTkrrPIQKXXsq6oR7S8G
t+NdlaeToMApdX976HfDohwxer5xL0HmejpGYDBNOnerD/1Pn24IezcHfXzBa0XkZOYgs6qPsADQ
/1BqAgPPIkckipgbhXPiLtwSH+mRDyeIcmlpJ0Yc23I2GEiGH3kQr1clQ1I6OgsmVbQRLkUbhJCJ
Y+GJcYdAXtmwDPfdCjvmPIDdt9PWbE8i+qsUm6JacYV56A8o7TkZGOZKjFzVlCJ6vWHPdBQnt4Le
PFYadIncNV2hAoMWBfKdMqhr091LYrdE6seFUYFrp4MjoKPbpCb4NvKX+Hrjj3DnVfKY99G6PW+l
Z9m/j3lmFVdK+xOfmVOzWg/J2QktiO2xR9NYXulqgAQg2KuxGDzo2Ic1iPZLoD2e6X83pvd+YVDa
QZKDFklgAm07RUlvySmx5oWv+wcmgpezNWmjP5irx3bkfVDPhtLwmqsuqHTdZYXEg0XAmWLXg55J
x9Jf2e2YEKJ3omPjNAPfGvfz9wXkC5FEqx7M26DxDMfhcxvinJfnHTt63tiYi5BnVrKa15DHZLP5
R6a6BDjlXF+JlyWN4eTlk69yRhDVUu3wccT2FUkPJoYN2vRnjvxcM53ldDmZIUDfXUw2C6dWk5EK
q8tUZWtqtaAbxtMA3NbfYprU+ikcRO5kp9ORK6qz6ZWJ/W2thPKB+RLjdV/WMU38sf0DT38bHmJ0
ugq8XaEwyhhdmI4iVauiexiSm8wjsm6HOPnKv0dy0u0Ys92lt2XMf2FhVXGzU+yfikD8qn71ol6P
IBfV7TppU6lv9QzOJV2ije9ubxf4NZlMMeWVkZkir+fv3rAPtfNlqVEfMMssVjug0AKWlKka1Nj4
3fdk+UMx1P9vNgKjBjfFXxfp/6Lyv6k8ZuZ+48/vYFDTH6Wk+HN3aV7yf6GJwxbi4bVvLYxWUKlG
41Vb8PEWxi0yRW5QQ+D27xXmkQazJsqX9AI+o3Ky5dOxOGQYIcNrkw/4gwZSM0/MUSyBJ+E2BWCs
/N1th7+liA10wbwzHzOETZ+8DkjSoKVWT1BPIhiDA4XGsE7NJQrv+ggA6yPWnGmk4dJPsXvllHoR
zwHCuC/axY5A03lm8mpEJf8bV8SQ+9Zr3f7a9BHdU2j5KQvXsbr3Bi/KXG/c34cZrtCr3aVqW4QH
oJJMzlGZClQdnaxMEDQyxf7XIj5l1MOwHumhBJ7SVpAZQIiNLCv2aRCuVbvC5ws5kVbM9PW75amm
LgyagPcY78uLeH85hTGk5GgzXKmSi8/d/lSi78F6rBzydgSUAFr/uDXWAV4GhBmIesBWmp3NWSJx
Pwziq968Ol34GQ8mA9mFClLHOd9Vum6dwhDnz3isO28NblRJ59I/He+eFPo5iNrDp41KEbZljh8N
LLSpYHnHrAoCn2c5wXZ3ZWqHuhx93Q2yxsR5QZvFJeSFnb187TlvwEPExsBvXlS0rUqBI1PKb8qn
fsTvg8R7GZv9QQFrjSUBKbbKAYHba2GCqBZcNaGjl48K/yKTvbpNcAxTWNkMyWVCDH8jgUAIeOSh
4QqFErTicU3ihKTA0l+SpEFjnMG1lOg5C0t2CO6wfB9TsxBhuPr/bDYB4AmeyYkv4quk3sKTVt5L
gpHEOx+/7qT/2AJj7CKzX8vM+jM+kyR54/1hUz0eJIF10sx/jG3gFtiTpnG5yH2myfFLqS7+VUyA
0xKb5JahAu6b9/ncu9W/z/U1ygu+TwH2qxq219uLSRsyBfJMhg+S2b/2+HyYlCa9+baMAoi4XtKU
6ow36hdBaL6TL10FExataPxO19YZm6iaekuuanAmUtcXxBmQN4W0HmVt2juYC8oe58/Yf7kyfEas
5KT5o7/jTEwK5ju8Mgo10mO8LbE8mlkZrcnJwpj02ozpUl5Suy3CNdbeI62NnrwptxwZzdPW/pu0
4GwG8a7vGzjplDdyBmY0oC08CKH4dnlZxroyNcJKfcrQqTDN2CXK2iUfpC9pNXh1WRHPcTRnacAM
g3f5FfCn7qBjRqsdglcnG+0amm4V/dK+PdNKsHpmyBsWRzFkQXCTffHwkhC+uouM6gyqg+/A7TkW
a6AUNR+qqcAPGm/uLKeigaTv87yOapWaVQziQX2XUdYF1M9wgZifyo8EZ7ALcEGO1zkB/ecmT1vH
Vb8xDINsBMDXAQgru+wb0yTH5KM7S1FrEGWNoX4ppBgBL0M4JgN9hyBexPRIYH3fYlrzmzlc90xO
qamdRBw289h80ELVAOAFnN05o8b7sx5Nw554s/jVbcXanH0PyxHXAxVHXPp/c1ntVFOhpyoDgwQC
cnDK5wBNnfZZqQDmCBMLRTJ7lAoHzAzrtkU3JVB2oQ0S734ORGuI1TVyLmDTb11ZtzT1VitQBGM6
JKiRX/rFDCpdSoj/3LFqRhpBNwS9uQgMN5NFr1Hn53HTEfpSsTq1qhXniJSNCKHimoLwdUguOSzl
J/daYnxW9D81/awG4L1cZEzWaMDS02W2XBJzNIAkwD9iFgw4QjzvqFuOG9YYPeOjqzEyKF4perSa
Y2TVqhsg+LJLOrjwQtxO4f9EsMVjuVKIHG1n+ONYmeU2WQvBIB1V6Te2C/enuCfXCL6OPSDytVAy
vzeJkiVlkaOpNCzeVl2D+HsXHMJU5co/oMsH1gJ/428DgPl6EPM+sxgIzn9TkPpPwcf7tT/pKuUP
w+qASaQO9f4L7r0r1R0fsNo5b7QqcZK+tjI3v20aoaMle9rjfmca8T2xIhA5qC7jyIVEHaZ19D2L
R7LiUW9xPeaZGkjPlvoihsMkm01Ixip/pktCK1wZv7OSmT/k8BpAY7ERXkUdoTEUDwFyIuABK7xR
dBW0Zpb2qldA7n+LBfjr7GhKhMft/wJtwOKXLYc/WRM0mX3nQjqYygjXMTdoeRcJNFq8UAYhV+NN
i8lfNe6VYed+RInXsJAF+Apc6lKGD4IEfndW9J/wSs2Xla1JudViNLYXLfRe8VfRc3qn3XCSOdyY
Yp30Iu1RBMgc8y6yAMubFi/oI/LcWqY/3UoQkUIMOm66MDk8JeLeV/GWDoTX/u7AilGg9cfgkIZ3
GO8Tt4QNam3WMBx6RevMg3puRGk8dZ3wmr0SjsLbxOS6oxJU5q5/OHT0FwPi5ZOVZZR3ZOhpssSO
njyVH/hWgdQtPpfFnSGTA5fe8LPx7G+1XYhvNPlrqRm3kNS0c4ieZWW6G4kvVSwcCERpjDIV2x/K
yy0Z+1QVo6HxR75vIHUs8/smOE0YhFT+XfOHqbc3miWShaJQUh3oxGRtQubfxON9u4zTF6vgcbb+
85HZE5R/LUNnxfyxleqxT9gt/8HfgskAmW4qEe8k/PJy0oI6klNiYR8otkLTkNGFHt/0g7wtL9q8
V8ZMNF1f8Xnxs4RnMfpU1H5Cy+/CpPFz9RbRjRZdomR9jlUa2dRmfxDbeX+zphz7EdzjuCNht1lB
9q/V+czuJNM+H2cDUNRdntOM/+uuOYjwJyjzo2Y44pb5JlS7a57bFPpwslUbBwkoS3IA3xXhBq9v
qagZvxP1MGSt4O5HB57LTOSEt78cxj8IMMpWNkhbDe+kB6rVDrJpMU8nX9ChMpjfYTwFMEKBuW1d
giN+nR9OQpOtyOJDMQdSs1+VnMXAcx3KmkCM1p+9m4myAXeF/ctIUfgpuyv1ixgR81OXEWRN/T7E
NYrBJaNmQbgiZmB8polzMk19YXoTeT2gy1vQUEC7kSisDbQhRvsvkJUEZXhsxDRn859OEAQFytG+
yiufzqUdTyyK/5+dBJnlU40NDXnJHMzAj5cqfCIA0NMj/8PKOY94srh4VutBGyGvs7KenfoOwkIV
Ef9ztxGy1nyrwrYhq25jgmnHwyOBHlU2HG7d2aTz5AuxdK0bCHlBP6S+JqAIq9/XD923yoOuTcVe
YBI/P1K4sOOOiTcJGymn2bPkSUWOiu7ot/zUZk4/X2YPwdf8H7PwpzqEHjHBpogS4rbPYmk7jEQL
e2+kkGXjbXPZNorCjPeRF9v9qsqWH7k7LTeTPLwn3hx562EXFmsaxyuSYhrGfTUy2h9wVvhDTTcO
yZ/xtkYO/Qn65E7e7Za2cc+zDEFGTzLaqNtvPpEEL84vrlAJcHwbnKbvSFR9jvQfNuYNk3JIV8xb
qJ3fxuX+RDtIYXCfnFG7GSvIiPvKkA2It159NKQTOqkR7VgxAz66OteLTonrCQ3vQ+Bt3kFuA9R2
SHJlC59YMnZUNxEzJ1h1BZJt9bz+VbrLuQXmUO9hlzmJ9ltf51xnvVCevKosntuBXx8o4FCS/PY/
0ZWQxEvXQSA+ryeMPKLDWGFhI+DchiujN4amJtC8KMxNUs8PA8UHU+VKmndca7tV6rzVZupW1rro
+LWNN37MZoz48wgXUvoDsTD+qplErqvih2vgkuwN9CC3t8YcBLLHedj9MBLlMWqtN/r12ShPFXqT
IDs8tixRJiBud0pPSlR45zfALBytRK3IiBjJHA4dOmT1Li0220RHEYVzefevoSqHyW0RKXE4MJTv
500BU88pMrLHuVFHYRx2KG3L4ZBB+C+ZtYSy50dRr+H2zlVw9oXgRhfs8OCHVkwI8lR+HtBUWRGH
ZhXtb5+0Abt24Pf36h+pa1t09xCC3CYEZTncX+1G7p7ub8EL7EGBqErQoVEYbA7GV8e26v3NAzHs
OG01b49qMh1XEQAzbjyNyg22669miAqbLhtBmA0tjJnigBpt+1PuWYp4sypFeXpmt52B6qvRcRHw
CS6nK7enucA0V+LnlmuW27sHUjD/V7kGNburXWEXnOcw1RPdpF+wJG097lTeW/x7Pyi+9v2KDAsM
81XqEoF6DrKE7Ysxh8wOp5o4v7tD9DDPsAloQHKqYs9KWV3WKLtgRdpLmweZ0nu3TrAUUlORocFR
lS2LMmcGZyHDKn3h7LJPlXx94FRsANd7Z2EeZ/80OQa2C4TAdOARa/Goo/zofiVHLIMpMcfBa8D9
pRcoGibQY+ahgtk7ze7rSD1kfLc0NoANyXjkuzcHju9+xwA0xniBdE2U/E+jeW+xqzvnz8a25bZZ
vEFatujZw9vDKCbC5CvRqA9CKXpIOPAx3Y/TdsjXBesawKh4t7Fc5FFDHDN1p4BBHfAiGv7uDejT
Lpx9mFipDo/HRlWzfhmfGNW4j9GOqcTtCgTXru0ZkRJNylJswxiFp8fzQUKx+5yHJ7CY1ZBsJkxC
Kfj6MVkk4lBiOpHRjuS+QD1eB+DO0PPyE/VkH5lCjvVGCuWB0sX09NnK7lnJohKdb0Sjye5+LsZU
PhanAdR2yDzbRmsl6oAIlS5k+ZGgO1ZtoxtSBkMyWCXUARJ6m83X7D+6+8Dqg3BTatnORe6BwTn8
Was7H4X0GBY2SoolTCHzpx4AVV9WENGwzF57KoCZ1VFCdThqEs6ZwBHD4gvXAEML3qM3hfg3lvyv
iNcuJHPVtv6NatOXM083EAnCTsjhtVyC4AepXNJaOo748wWkvvK/NTS6vM+nWIOEdk5jPEf1sjed
e+u2d6fK3xCMSQn1PuRRbCx9cJRzms3So4qxjYk7z8FzarK8Yg4Zd2N4PzmtHzze9IcC14tGZA/C
G50oc+0gG7jrcZFNpHVPGsCbPMzKi7m4OBdVHOtwC3ogA8F68DHZuiZD5EGAfqjh0IfpQg6LLaU6
6xw0bnygRRbKGMOCve6BQS5tF1w3xgRMlrukOihOhnZoczTqZzoNMfBg8eyOmbFD6w+Dy/2vAcc4
PY+d/OElB+/KlqfpcjmjqZU7TU6u4qlnRWvfBWNnPIetL2wtM3cX2ObMCNlvVylFmkt2lGbqNLJY
GHemEvgmAAoUToOwSSbh0iEgca3AuhZ1svFzrabwtOIvt8DgclaVEpfdxH8pB4vpnX+7Vyo7ffWe
a3IOnwVFFdXKEVILxmpqkVRYUOQzAnT2aydbnNaz1jkcEe6n7kIQqS10ThZQvn2zb/1m/iEvPDzV
JhVxf68Px7jae7BwlyU9FO9TYLYY4McXwuC2VD0EXOYIh5JkRnCT3CaTIvYk5Via1l6z2wazDp+I
pnNjFQtebhHrCy7PaWyRSTDtZznOUYQSoUxYlnEWY+thsnnNlDO4/W1xmFD7vHQTV4dPQ9a2O/Md
9U1DT6XHjT0sCDkbnrNq+BUh7pKG6Z5t+aVFyJOk5+ZcNw9kakeBYBdK55YNMJ/YFa4snSJ3V/T4
xhHrCNdpkOvkPQiL2RRNSaLjR0ZGjDX7dd5nJ5EXtfvfyxHPNlKCS0ZZlaOXBAY/4JoWBQpj83X+
FXMtKvdnV92gMeYsp8HWXs+agckf5fsaNiOTkaO/X1TQrR5FCGiizAXnaUpLkatZKXfQ2k7oXT9F
hO13I8a6HbRHePX+QihA5rlh9wY0PyEfNcLomj2wS+2K31m1Xoj1pxIdehPoqi9/5fFfU2+bq1Bl
RHIbkOzCBa6tqQsD4k5wX2/+TTUm2cMOoF1TVRA5Tc7isNQblXeQsN7MH30utktA7y8MBJmyevCv
33Fv4cLt2sGeFm+0n6b46ePPQ0e9OWEcVqcd7n9gtDXefD8QVIqVtj65H8NBhj2wSiT1uGtwYfbN
wLZJshgv0CX0Y6c8qjmDyYR9IBcPreE9vuTO/vXAmJJKK1D6ukUR5RWLMUqX6tiz/0zjN0Hba1WI
aRJbyZ9DFiffP6Dq4q61EQWGrCrKVyp632Rg6dkXgJK358LJrTiEl0XSI2S5iOdCvRHyAoLxY9XB
b2CM6TCLuSuKTkQk1yFZk2/6K4jjO9Cz+DhRmhD/AXwvv+CzVDvWKIPHHmCEOQIcB0+vjLZ70zKa
FOMP8Z+zh1A4vPSXQv0x4ecqX84E2wIUJzN/f0PTJ1zy0RJXBX5jwp66ImSa/meagLRnURC6qKj1
/bF/7HAKtYNKinczAGWDqmq8B9ZAZZj/3KYGJd9qnbcLQgEfp/MCqchmjrCUz/yy4TZP2S7qw+VP
Y2y+OO30sD/jKQEbZoFWDJrK4ciANwkcZBd8DcyMqZOrvuQ5gfHO8yg5NGBbz9UOkIG0QMlq3iyx
l0Pisd5uyopSRiM9bzsYrQvVIPjLPjUlDFpGJcYNOm2+1Zh4H6OplY/7B7NZFy2Q8klGNFPBGDmZ
WY8dU7c1XIyVj/rXlhtK0xtgwmELWqCx61Sz/LV0QKU5MlxBnQOBkFhSx/InLDPNHIaRjovVJr60
iSQtkMLYqAX0Y0dZRoF8BKLKlExhSRbIiPH6Q02sgtXbHf8K14BAM7ks/bwuSlVPSnJpCaUSHb0E
x/b869hD/VOHO2HWpVvQY28JTj1efcpMBogrpcqE6epvpj6/2grz+gLrKjjIXyQnG59AoSkEQLC1
QHZW57f31xNEPjmP/GvJ5hLwXbp0UmOkZ05hCWeN3cxz3MmgHCN9Bdsj4/c1ECBgs2XxelBboL7z
CPkgyWwAz81k82lSYtFYBlH0S5fEaKXndgskn2cbuogOvN0TmvCgHzMoD0WGyHAEq/kWF1SmVieY
nMY02+qndddzfXeMbzZxh3nD1IU2LpiGe6fPXOAxtshqx0F2r6HFi1nvFBf5SzYLOxJ7pst+Xj3m
WpkRGL85WyOdHvI3YbRryfLz0kfIeA8wW7OvVAdGi+jRBX0nCUShL+u8uYobnE5j9NAxYbMp8PRV
aM3ST8cwox7C9da3Uw2KQoNCZhjU+CBbhjuQvGy3VTvTmW4Pcznmfg9zfxK9IkMyzo2MJWJly+H6
9ZH03gkJSWIeQhxyXINC5dDZ5ewPbWE6BHpOy6eebyYd6oGlUQTH8AJzfgu/buRehgEbC43TE60C
+GoQX+5fQZ0iyKoOZVgfwmopUxjpNGcsA3Gg6CIo2BFBzwQW+HnQAVmp/usc45HZQ27vm7RHZwot
xL7EW+v1vcwRW1+fT556GeVz/j3V7gTiW3nCkPQwjzxoTAayn3MIkvw41Qk371AMM3hS56AOusPf
ftyG5eHqS5jvZ3I19SEOQcvuyCAXm0yYiCgD8P8kvT+sl8Jv5w/PBdrHgmr0gcrA6rZfo6pFX8UY
pPfYx1vIWtNB3MjW4C3a50bsiMBtn4XknuD+mF3P/y2ukAJ9BBAOvLOLm4xoAeQKRXv1XJ4V6c30
1a4Lekh3ALcqE9ZDTBLPPuRZKcLw6N6xqJEUIfUcD5Q+6fUuOQZuHiOZyqOMgj8xv9YvF3OP/g5a
/KlssWgKXKH/Z069G2jbjvX/jvNLEz5bhpR8KRefRMG3UIYgt6ns/7WJP9ZW7DQwYObKaduMnoRQ
Fs9fSUe/8tv6pqMXruvWxWydWnkJ01n4lRAKpSY404qt1eD46tqEd4AksKO7+uYT9hhCSpeML9AS
RkwS2hVqTrUyjL3etEt+2uaKkS7KUKuTfqDbkJYfIpp8owmyRit/tVlpogGmN5fhZfhDmgctvL5I
xLkyop54cNWipr0gXhIeJ1SbykTmugB8Nh1/rcbBchb8G3U0BlepTtFeOsImMfpMM7Q/fXtITBfH
edF6RNCxfXT9mIR9BkJaV+ZIaSIVjm60iuI1MTlrN0IWM1lftqu0i5Qv1LmA+miuqrO4eF6XrccL
lVdpGXHIaEVyeVySJnE6GkkZWVAHfZclltnAC+5HXfQwIvrUymDBCfqAYgkXnnUhSsVQifNu6per
JNBkmK90cFomme7mMt83zWRh0Ppvt8SuvKGDq2twCJvtyv8eYyOqZBASfVOyvji8G7+QnAfni4yC
/IusgaWQ1O36XB+kZHuCgS8ahSg6+cATevCCDgGz0xISS5NK+zpucp4VD0Uw0lPLPIhMSoURu3MQ
Lu5Z3a1AgIKgdbJCqFq37DaTprh29S7ICY7lx09GZbVm1WTujOvNC6Jew89XwnUeSeFHj4YKwIaX
PptBcWZ+WCyVhaaR0XNAZ23LvWrRHm4/KAv5SODKkXEYnmh5lO4Nhtfxi/r6w7nUCe7Cmz+HP526
c3L9yH7882cg2hUu+CxVdDAhZqVLZr9ulOKNlhjAbWiqCyZFdxzXcaEcqJCxVcQgaLQiTS7H6mCM
K+DUqollxq6GpGDcn+P5pp+2lLz7154JBKrx+Yi2CHXI+zbMIl96EzHqe+1v8bCVzDlMxMOJFAMw
RDt2/xJyH5C63n0It+6Vh7D7O1RMehqmgN1IFEJ9Drq3K8zel+JMhG0szLmCCfoTcPIra8GL+9N3
7j8siXGRBo9m47IMp0wM25Wuxluneamg5rlkkCP/86qtgStshfqFBXqmTsIpHBzAWJj/7SV/IBE5
ynhv94ycWq36mVKwh+uo2AuNusR0IdDMpm0ETBMMQdMRfG/Tk9n8mMFe/aLWmlU6BS/ckN4qxUkn
b6LgnihbZm5I0YGPoTk0iI60s5oUVbx12zIb84DUc/MgO2MttaNMRqdXcBxFO5WRVCOW/3A8/Jjr
0J2ldFHiBlb5YwfmEzxmRp1N7iNkv8+X6DBdcysOr+C5AEhDY1wf5JzS9gBrkbUKJa/inYacU9TU
KWxUXtmGzOqWh2V896JdDCgMFBzHOPgCo/DaPZcxSpvNyFyVy3vMXjyzy9/W4VtwP0nMGpTo5NWb
aGu6U40SGBdYGGby92LXVacM46xnE1WWWvTrT5wSuPgqBQsLBnqVHCgnu7uNKhicUvPYZ+C8di8q
Hj1s4QiquHXqIQNsVWIidtCsKUsT80aeC0pU2YX2eIEhGkHYiTj38IzjIHOB6LQw862+C7QCOjJg
Pn4Oljg/UV10u21ExToDPsRiKIpOVl4jr/eCz8ZR5wU/o2v6PwlmrhsFHp0wxz5ZYY/OM7Nai0q9
5zwB7OfMGA4HNPw8DdGdoyP4Yuuh0waEB4n0rejJGtzw+FaVFCo3i04Pdf9uQ4qp3xaLUllhBIiH
PBA0zB40FxsCdR6C4kEsgZHRpUAds99DTBMoRhz6SzKMmXCcTZxpvpBq4X0XpUPqzanOpqdngYnd
ChdJkyFxvdNBCXxvJym1vE6Jx5dJqNGS+Ck/D3v2y5haUCMQRUPs7M6NcbPthnJBRXJuE0iIJAWA
lTQKlGP3H26uxn/Bmrt45P1B0DTVZT+Mb5QZM0ZOYV4z2wNF4Kt6OlySWXbyPX3WfC1HRfa7zNVR
qJayvzw4KUcEp/vFS2+ve6HTBO8UDB1BfcdxmDdFNJwJJOl5BktlirZcX9p20NFDni04FNKJ2++s
1Owz6il+8UPoZxnqKuVe4DSGM1tVlUxYdDuO1xza8Gw21mqEtJmxzRmqYbOi6+Bes98c6RVjcjxV
19Xlvljwp8hOwUlFwhiquFZFg5CsQtgZPsIJ2nbj/k9aUilsBVqm9kH2im1xMZ29SghO6h4RzjS1
sbg6XhwQXd90PTRUkKVCGMgsNqgvuUvHij8PLd/Y0uS8cU3k3MdFCocQoNMvUyVHsyQF1fASYtX4
mtycicJZWoeiJwWIQU2fXMveNcQ5l5tpXjpT8nSEMDY6wgm6g40W4Gc1sC2OoCSyVAC/I2LUvxF0
Xezp43iSlolzoRSPsKYgrg6X7ykQsQE9yaSq4vYe8UqfjWbY30C0kfhl2avAoRc6phUGMaSx9z40
NOSV0YuYPREthLu3ut3SSYTWSpM5VhL2KD/ipxsesmbVnxiVtC2diIBPGWO0ZnkU5elId6TST3pb
7Uv7FKFxbBjy58isZX22UQ5yI17ib4h+bF3YpCMfzXZ7pjqn1XSDNxtSDkJXJe4G2Pj1YxELI6NN
aNxAmQ4I+sL4aAufdBBRgejQ4V848a0BkEaQBg5g7wacUKTQbjj9ysVhXGPGDpjcxwWEq0+inxbJ
UwZyJag31ubgOatHwLefjqa2syNv564/PzYg1O+c4OZrsuz69m//ioXbvHnMXD3SfjADZQViubgv
PszpU8qQp1vOIz1BfGWPMOPaiKU3fUrbi7lzH6aYyOhOBVRifjohWcgfhHqWZO4e1MUqxVIk/28z
Gi1SaQcsY0wk255FvgfZukgElYJclngwXhS9PgYl3V0ZJFsU1+HztYDakFiEPzdZTe74BoyIqY7V
rw1B2wUOhY4k4LZ6M4PFb5srM9hb7SKwYv/P7eOePXMfgNDuLofVOg/Vk3FUvr/sgQdv6SemfAgA
FrRgcTVUSo459xb7JgMmU1qCnVWBqdx/KYZDkRArFZG0XgFgksIkBCW5Radij5qko4SLfJNX2pNs
W1DA2MB/gniSkbsJ4OC9h7E52VkGcEPivmUxmjoUnSXlzZsN/6luWZf5ILDEHu+eE2DuR4Lp4Dex
KtM5fokJeHu2hcCs3q5Woytf4FxMTWT4OA15bNPk9WGd8s6aBbb02S1zO6yCq8xyOxd7IXRpDGEn
tJw4KT5j1/OJ1gDADSkDqsRRYLy3Vrq/FpKxOYoKduGS+gxZowkTrDge6tEa9U32vopoCLkj8TMl
TX5SK9WBU8wLec0zdRKK2hb1QOZhWTbKwEUosIsE/gFjCNGo8QP2gptOudSwQqlJA1W6BWslB6rL
QO4VnBozm8zeP3YKj4z1n6HSj72qiLh4TaI229OZXJP8D5V8scphqhgqKNeqvBWr85VdbBw1aEiX
zwzr2JwCXbunF+dUiyc2krRRrq0vwZFzR4VNU2hVgxL3hBNy1nBsFM3QgNjW7OK4x9FveixwTL+U
5NiRgkUY6t9u3HK+MIU7FrT49GXuexLOQoNo164hZTSxt5Zl+3qhBaXyQIcEm45HzxQ6A8oAIDH9
dqpsHieQs9BPCSdvw4y39TCFm029JN2K0EFSOCLOpzjhoEx+bOjs2xAnsDHbRerAvK28U281uiK9
M69vavki1/XSzSC2Ne239PAVb/FSHmWk1HRlkE4JaDz6wBzZxPOkmtHXauo3oO9Dyo8Ar6FWj4iT
Rz51XK/JRly+XGp3SsSqEf1TJJhaaW3sgByEZPZSE3VVRGgOv9Ji6FKuwwvQAClKA0wyIRASiNHt
FdCXyOZkHqms3dWyMbygqe+tJtS1E0Qz80hTP2S0hBwK+8ni+On5xOInrkV/tNu6dw9ySr/S08Kp
tC0eqjhR++gtAmV2MKW20ZxY2i9lcS+mNNYSV/yPLH47dGvNxSYaKuakjF97UuNI5H+pvl7jwNG+
IEzHIr1+9tjVBe5Ea614J6usSioLXvPIBg/hFIlSPn69Acr7JJDO4zCu+z2eVw70wKRMJ2HNzDEi
plo2X9rs+7JeM+Zo27gL1A2Axe4Cdyndj8W/V0o3pdDQxlKSipBO2FghuqoAEsOPX3qcBfMPCdXd
0VGaSqh6Uh0FGGKriTPsFm7VMA4VZJZydcm57H03SNOzfdXwxf9F2CTVB+Kd7mBCJOlDDAbNgkcB
IvI4aIqIEJQKtzBXqOr19Nu7ddEBg+70e+ooRA/2aRTWrwSD1lAViJhstSprGgP43qub3tp5H7MW
8OoxiKRPtvZ0kzmHo+rVrONlSgPO6Mo/wyhyLq9+xt/7bBuRRBVqOtGNTdTnxEIIc8qetlFA2sKA
kOZ9c2K9XB5ymBgJI/2zG8kzSkX4oTd8GQYONhrlIu9MPOfJnC6SFSxNHdw88lgfXA2aVMxmLNRw
bw+Alvs54KXl5gBtFDJMfLw1ShooiYKCOE7fvdUfen5SBqMdL5PUgNTuCfQoGkvZQgp1fcTOpbUC
RB2mW+S9Num2JJNxeBEUrx4HWSCHE5DvsI8kYlAUNCYsRY4/ssVH0NAE0RADP6VilEAcOrGDsRK5
Vtgzh/kWuaqZ3XWdbTd4BMAFIVUeH50IkaznGl2tY6lyFbsBZVhMvTqtbKbD2CHSHmsMk+iqAfu0
IcHbeldWS7oea6YfmTjbr8te+GRm/mB8JFRx/uowMt6F6QZjFLW7VUU0zUCl+hseQdvFbTd0xTJ+
u3qaK6bUJyOGY4Sv6y/hIrY0xI7Afa60zj/rynXCUVL2FCtw5YNk3XaP7vT4h69E63xOyrAOA2HN
T1Huqi+g5j9WJ+cv9y6hffRBZX4K8hbz85G+eo4oyuT8GsEgziOSeTN48BuNpWNi/MIFVAU1zXbO
9eNey8s8RsyiNts6D29Hd+9AWAZED2SHJ62f+9E0t6+ZzSQbH5hNGzQSm9udUzd5wEvC+3SAOz4S
FwAMQyfMSmk8zLJWy18rs6wwBTYArFW907QA+vnhOTchpLO07dCzfY3VHrAMHtYKdPP5u51wpFKt
jVb3Ofw/wj6EaGQzxbvhpTPQZ5GQuVdE1HyHUXiOcQQ4nZZWL3NuGHWVT1IPP5Ktr5SPeOtEFqU8
3DGEG3S6JgKKaewdGTGbETqV7pTYiQAMfLMjOhzaxJqYirT4MTYuasJhmio3F9xbBGispH1RrOsc
6XumRfCWewCOBE8HVvisEJmGajTb93vfvT3Fbo1APmlz37AW7k6P6W1Fopq0AKDiDWc/T2LGhoMj
YMfT3BSaLYw+7diwGJqT5VVMnCsX9xoYnM87dslSf1Y+kGoETIZqy/n27W7DPtxnhIBcOopYiu/K
ZlrzB2jENnOEuOqZxqIB0eSmbWztJrtorWbYKRNc9IziqHzicaD8UU4QnO475Vj3Gjrc6NmMG9tz
MKuCPjqfwTdY/7127gXkDQ77CWoXYJ2dZelxYFzoa0ebsZXq4w5li28neUGninYOYr0y3b6JRgDS
5OaHvp2u2kVUWeLY6TrYiH0yb1MR/KqbhwbmrBC4m/fUCIHyVqoWXhlEE5ivbCbpbXs5SQ+akNTV
v6iGgaFnqfYIDGDtQ4LB1d2lFObH8snULsc0HjqT32hhjUDusdoB/Y72pWdKBn4dt2AZM+watYez
l1w1WrsVxPLOukSvbfIwNDW/nZFm+XyTulmzh3HMT0VM9ZMjejCDcxOQQ1EU9sZpOuN3k1h9Mqa+
Jc/2/mZZxu5RlOMA8QfPpecws/f3S4417T2fSenL2FdiAdC6ckj1v0G+QS3hz6p05UAelMDmpn2Q
oyePfDdlMxJ5sBjR1Nl+TGUrdB1JedFmOA5Kc9Kv4zcbbqXDU7s0X/Z3MuU/YTHWgT5vnsGb3iBZ
Ah7mKrcx56/cZADlVTA8Iv/14+pszfTmrzrkQAce43p8zQsTNL60xpBi76OiW2n63QNd0wqKv1fQ
1GKMPhxK7DnBY3I8olMr0bokD/TF6KOmFz9ah5nnowxjKK4D42U8lqrSVigY7taxOOoNC1sPUaM0
fP7eoE2p7Rs2HLcxnAeQIBEzCdnWZZKf+GNqgtql9oSoyVKv4EJtlMsYoibA4DxMOAMgRkfnmNcg
4u0u4DqLeGhNgyqJgn/1CrbIXi44IMOCTaqBlSor1aphUMwTSH+EjV7oX+o7sMP3DWVATu+aqa6d
/KlbVkUhf8qvX8P9ZJJ4NvX+XXd6JOX7Vf+WAvQKvAtgu/+j+xsbYp2TowwnWbQqKMjRV4gR8irA
JkmkCjuQgQcJJeGON0hcxBs7Djth6geCthBTLxpIXWae1+EzU3Gj99Bv63NCeHKZQoEfEoxNdrpn
hOXejyrnMsNavO1Qqc43QXSbqhddyvRH80DvNidVG5RLwFtSsl0EVZZ5/b0U8cLQqJJzdC9rB7jP
jDa69p7duvEg/Yu2JU77Iojrk02ipPemms5p0SKueo0YkyVUUUzJBwTDaMgMa3RiSt8oVbb3Q/BZ
Cjm498e6IGPpbnVmzLi5Vh72VRMZHSKB5gP7gmfEIsQgCC2oaPA3jIp4oDDXSSLj45tgeg4peZXG
rQzURxOcgCppqSqvRNVdf8st4zN5U2A0huA7V120MgruEcJyjHQCr4r/PxD5amT4sjkBqDIVwonU
RLzXCVOgU+rrGxxTtm+qer/RBLOQ9FMiRYZjEOlnZ8M8XOpXRup/DRWINRmrpdVltFSWq3Bb4wQ3
4wqlyKDh4SRNzVBYHKnjAqBZq97oJwgL0Hzck7lhlyaoHbOnu4Bype4iuJkbqjMb0ltpNgrb9V1L
9CsCH8zNVlNg2wEjqqIPhUnit00QgP1kgVO7IqUwpOYq1xgI3w3+6ix9IJTdbOviNyf5j/+5U1w2
WDMmfwyxHvzTmYGeJHIlfru5Dr0AD11/f1u5+9tKTaa+/Wbg/tjSLJSMKacVcG6F4SVt3A0gGSxs
8fhmrAYhuBaOs8KyM+BVI4A6gT/aiwjGKYMAcSR5ESSyyX6SFiMk9WJdzLVAhexCLi7h794dnHG5
x67mgkGENHJtHYuYNFHU2etMIqOdJ9wPq2XjSb+enPv+a/fcdFzTMpx8Koo3PCKAnaxwTkZgpgHs
3KxtoSt+BUxTaLr0Lcbsd2fap/eDdJbNYl3hnfLd86hbht3J1tniDwVOGpN/GvKtz8937LZDIyGc
y4NurCGz+gvbzFKgY1hjezOObeCQubXjs7oDvS063Vuxd4cEAJsGE7p+pN20BQmXntKiXA+maN57
mjjyEcYqYzBmFyBZ8ChkH63BDixpxdhspZpWin5agKSqPYaEEfju1kBbzuXHrZX6acmsEL1+dMgp
QlECb2QTuDfLaVxODs4aJ8uTJKyAwm+BZvvNQN6xSNAWkK63L0LC2BguNXmH6wVFfGTg9gLUpDTl
0BQZL8zaTrLX+pk/8/cHR6QYkTxPMvh8j49Jy/2F8em/55xgrLILZgcSR6IP4Ns251vCi8RFchAS
Y/YloVQQTz2JdpJZUJ035xzSS5LISAr6QzXIkorYzr3VbNJSzztQ6d2vT5rgNTwawBWDmCkdUfot
aUQb+AwxIu7D8c68A8YZXUxPmhFsjtPBg8GrYnkBHxIsC3qBfkxxtSk8FcUiw6hMbm986mgzUq0p
MtJMnvCdb/atrI3n5wboouC9tK+xtly9aFfbhWbuubsE3NQIQWCK9x9hmzJyl4lJDNrQwsPqpjEL
lFum+H2lGHGBZ9fQOH16YiK0WIqAXLRpuHVHNjV1NACcwKuRMCLmWI1b5CNu3/qAGc7gn4u4UvJK
CnS7Lcsc1Dk5yQi3nr83eg4SaZqX0j5d33mZZxlXfmlD8008N0nc+s/AVqJJxoPhEY0OgoxC8LFo
dE3PShZSwbaAZ3CqXKEB954fOMYIq2iaUiVwHGdmXrM93uYuJbuhZ6K5CfkegH0GDqznebno/+8V
tJa9KcE03fTHS8ZxP991xpJhKNyJFcXzKSapRge236GCPK0NhBRs9NttlcsOGT9smh3gPgK3f9sG
aPy657BAYbvaZgLt1W346/QZYv2qTfqWiqejvR8LGuMVLAxzAK++OrEmDT42156cK89hu77E7Bof
N6Ns4SxH8xBoRW8iLFEjwrBQoP6kyIMKbg3rll4GJZoxp9JbKAe1bqYIQOj1EYLctkK8SgLATLyU
uj7iQeoZs26C5wTsSn3ZDabRgRKz9Y3DgZlBuyiKwizcU4iQ8ykFrYoSeXCsiLIKYD9y3hedtVGj
snwPtGG5Fa9VXAStvrKSE/Ykhlg/ScxGNFogE3lyTAJ2U1fS/A7ppTl9Z3TICJOngcg8iMR7C3IM
PKgMGgU0fvAjnFvdvqh7J1tZ8LOeZZacu64MddLsciayuAxaYS6VsqSmf9NQzxWrEUgyouo9KbAG
O8oWET3ziTZ/Qi7LKWBBNSvQD9M6JrsUSa4npakvKvT3TLJioTB5kA9oIu0fOI4sQ8qHtp15V6hP
BlGETnXFcmtgpTO0qoGRqtXhB1sL6KdGM7x2yiuLoCWnhW5fteEjAhwJ/L8rm0GfqgeDhKOi4ACB
lkSbjyo8EBnciXs7rKhh+PzyMWbWS+uAPE3Tv1vSJ0Q3bqNYZJ3LLyPDNWHPxq6BEsEUK+OnFXk9
TtmCju/raOfFf+YEWH+cDTjyXiK/92RYYk4S1L3nIQ/s4AeTs13rM81rrqu2h5IlciGJbq1xJmo/
hOQkRA26GZlcOL7KFZpLnRE2LIi5B0U3dEyrdEv8WW8wRABmNyOTej9UqeUMOhUZiRIehZWm3LNm
lm0BYbMbkLF/ltwXkmN1N9HVqYOPFKd7VgEzf5rcbiolKN6wbLGxgFjVsJqx1oaVITyC1jFuv85c
Trl4r4nCN1KgSqW13l1qcpfsqhGb3yLauVMkl3tWRuQKi65Xmzr5n5chgw1XSGxL5vlymODOIX5e
x4W5aJzNuVefMX4RjKJgW1dYhmZTqMiHeGdihW5RnSqDaycM4kwfJ4bXfhpRvUTCITQayop/omgg
NYagZ/4O5+qe8WnHZplhSIz3Jn9qUGGWagNWyjFHFu6gqzrq0+OWHIAgfITDACWX6h3MNYS73O8O
cJpq0cvJZHlufbgnWrpNpFJiIvOTzZDJOqGQYCOidHsfBzafvmj0sbkPsqG9ORmPsUFhkx/0HPEf
afYB7lW5GNx/Nn6CJ0KcnlGe8E+YM0PPvg4dmp1detnA/KoVC7yJle0rqOUMPDjF4GHQ87/w+jnV
wG7h/CqG3vq3JIt5GK/ysdmSijIh3sEZTXtZgbUzosBASVgZWFxwCcta7gcHOjDC6MsesgnedNoV
GktjxQNLfP/T6aPvMdm6EKAy1POArsdNzHI3IkuaYoGlEuCkU82l06XgHvgXn8ZgnKOGvGGaXbpy
nhwIuISpIlKpFpJNdOz1K9O2SbbhXW/zUzALLq0VF5jeXUgwc8211ex8s9Jm/2DIigKXGBCMifkJ
VsbQz3PniHDK0QKe2WI7bj4mteeoQ8IouecDd6IyfBw0Kg6mKWnxZEwjD1F7dKvd5XvqHISDcOcZ
BrIgdXLtNdpk0v6SnoypKwYu6UTuNCmXv7QNTlXOzbv8S0Dizrz9xn+zjhhwzzPluwQlwPjGxaO2
ecZiN9dkecEsGAuFHzNe6HlQXlOD/jbVyUlvQTrxqI/hgvvrB8NEfZApEwTRHZiHPVYz921F4AbF
S82vrl/CN3OSAt8mP/cwI7UHt5aWHqsPzOLVgEv3K2xQsRf1IceYG59HIxtrmLiP6qIFoCWdfjwx
EQMG2fJXKSwTHDAvcIhc1T1L497HrFL98O5mfUnCNlJklBDqwbEtxyY0MtLyycyr+2UIpec3lHCM
2No9LvGhUuf8OZZ/5YDWb7qmxuS+XtG4+jC8MXt2oOq1PPXdqSPN72qXjaMS5CcgVLfaau8xd+LQ
B/s1JvnUepv1iaOCGy+YHjQwuhcUtS0E1FNbI3le5Us8bO2m7iCsAZLM8zYkS+8gJaFMF6Zr6Lub
DRmPKcqFvrKK2aUz4gyLAgBtlGkVFaP91ccOcXS+1jxc6OlQkXb2fd/1/SNvZAnD2cToC57pXet4
DeRgNxt7A/V29OjKXe/NNIrYHHyAMKwpnYrExmFpAx9a4bXXpZ/FGsgYTag9Os0tw98QSmpqkHiw
rtDl361zbQaOnq8QkenXYvQr4U5/9JN9bGdeGJ3SpuUZahnEUyLFhdwdmlwptr+X0otDFcH7fWFA
lNuy25u1ithLUIZ11GniUknvbB5d0H+MEgSajqLW5m1J4p9tk/CxIQdhh84CNZda2o99P4/lRdNF
pjN9Ge3VW+R2iwOD2P/bbuG1GmqQ2KULjZrRxUi8EdMOwhNxDqrRUdXnOIlCHaIiGZckTUD4UC4R
8TUzUe26Cgr9sSUA9Nk28cYUAT4rgElkemdTIqNZL4KZVS09+wazfVHav62blVRl4xdYtgzOsep2
JQShB2+RM1o/RkDfazAhyeOoK6FBQ4kR9e+c82TVfPIRrtEuAsPrpdO3M8E1mgnRE3c81Uk/A6Iy
1WqRVnOX1/92sCVkAGChGuteoXANMBtHXNzuuC76yyN+CDVRooVmuHi0bSE7ArsSjldqzn4imh3x
LgWnJn7vhSqyv69RXp56e9FRu9FMIv+RtwDja0oscYVUzAxllK28oZjjfY41dT4l/SmEqDDUNLLK
Mmhu5+IfAdeqHSGUb3Au0W1fVTjZgk98lvI9RdfvJ3lNl2gDM/GQsqF1EyGYsjGgkw258Z2HQvlQ
cqNxDies0Eznp8ItrLn4aRhz9kmKqKuCSlmQbOVZ6sKljtY1GD8RJqAm7odGrL9yPt13fwmqH8wd
Vm4TRgUfKgfpV673V9y1f0bltiaBvr+a8Q/hhRxRg9vzJvJ1esGa/wVi2IzsEGz/9rnE0lrUcXij
ixzJXcvS55t4KZXMlaQ840l8Zy/uqya7Y98xO1RO1ZJqqAvDlcVZu7PW4Erz2UTTQ6vbXQCnR312
Cn+34qH/PU3/uhzGdMZZ4v1BoXxXZcc04muDELPpkbvHGsXfbYhIUR12op6oG3roNvc9DjmfQydR
CxvwPKnDVeCxnSufg7VCuiANcZnFbKeIwe+Dw0B5T6dS08DIMTH90/j1pbeae4H2Wn4sb5LYnI9G
ELnTBXrwVoQANsOF96afOxuYghKzFwL3wYHX6FOShxd+8o14leodvUDaJtih9cWwTcoYdPgHXZCY
kpQS3YvpB4NbjgdHieHHwHIdyJFVAGdujAJoc71ZkXLj+tOGeksfUUxag5mayaMrLRpoep8KXtY3
qZ+fKdYksAuFswGauHq9/YYP4UsMLfLpqIaPFZnDPbkfzCbAAVrAOJObeJzvJtSb/+LW7XDMh4zg
NNU+0wOVn5fZOkBwSxR00jGqjc3AffJar+8B9DLZyWgfC1ZlYH02ty06II8kasXB7gJ98AACTlzn
AB1c84dzYYjc1DnV/OWLh68otakUe90X/d7STHZZoxJab6hB8ervHPUN/SXQVdNpg5Dp2pTpfKVn
6ipvtBbPJRG8YUn9jMdRQYNRYkGHTuVZAHfgaIcHd3KPOhLkoARK7SNyY3g4BqqKr6zIQ/GcsjVx
pWQE6TaPVyNXEDu1EPv2odHuO3bqak0N6jcv3C5JaU8lZu1RdQNQR4iPQhL34YavC+vA6j+rhMq2
8MVEKuPKgRIo8INnnaOgEyntO9cLfwSoonbcLlZUSfe0sMIqg8rYeJllt9fa4qJRxPwzY3Eg6yos
MHtgvhizyK5cEzkAzgVGKOn+cdMwTYtLRbxTO+WnEPSiMdO9u/L7S1epSoCVd7Hro0WRG/2U++M/
IFAlgUUfOMLSvvtyhpVAXe5TEX3vvDohfgxAiIeBNA3AoyAnS539reQxuCGWZQ/1V7jk40KHxzQE
8aZriOdOMm09Xynybjb9cwC8sOsmk9A0UQcDgx46GWzSssM4VzSd25JOoybvzSpmOuIh8ldcnxbI
auvejamkZEzjq+4mAVUmy61jfTZH4KDNN+f3yKZcID9HSy+gdzWC9e+mVs9k8aER8QyFufA7qSwh
S/PQKLw2911mqb3JwG4TR8t7FY0Fa214h7yaycWVccK9qjZnYEshLb7mDCMkvKKw8pH7HKSYk1Q4
mly+3rw4c25ZNlmj8ifY0bgMsb7lKudARI+NY4R21WXCee4Pz/dPPVzjFEuIkF6rzZHGyj/npmh/
YKCcT8L3/Hd4BO7HZLCEXoaqnp9+a+nnHp1+zIQUdvlYOyRrMz21GQ2wfIFuvfnKe1Rjim6iskRQ
SOTz5YuehnzxlTg13DZ0qPj+E3EmaLDr6DLctILnZU9hLVhTIzddVXx7KDExhKLOh5WM2lLxPHlE
FlPmUJ67QD/i9RJaA6FOBC+M7kQri91twZY5rp+6QEKR7qzsRtttDZaEg3e62e5lC0okIYc+p2N/
eBCAYdRGndiuTu7qm7as3/4+AtFCyzGUcbf/Y1iXMNNXQeR2PsS8bXsssyDDNWEVNQHeKR9zWTLJ
QHpm7ljSJnCzgsVgPjaND3t4u0WhJI9GhmtxiulH8jxxFp6+9uPfK1tAHu+TdDYrp1QU9bK/10Vz
gItAjsW3j+Sv7iwObFlWgw37+twBTKak9xxxVBMIPU/ExaC5gJ8iOQQHRrbNMvSQ6FwF4L7euRKe
4aNxCLN8HqIekhpKKd+W22TVJFVpmycwEmlvKU0A9GMpJ8BaHDxtE4uRLYOxk314iM9AO6J+dQDv
F4QeiOtZKmTN0QqkMLGU1Tcm5C4FS18MEk2Dn2eUSSfbZq40q0NJ8Qu/F3zYjsSlke9o3dO8mcWE
W+OC1qrpq4bYgIRWRJKVydVAG2Fym2E1jDVgYQzrTXgH5A6kcxVoBTghjMecwbRbbeKYJ1oHVc8D
aUK5hae/ojyNbzE00MeP0kEmzDqex2ksC+Zqwy5KvzC7R8hemszpXG9sIoBnDJwQFWXfYKSVcGfk
lhjC8cSQUfjgIU7k4YU3TgBnieYN2Uk8AIfIK+yZ/ZzYDlOCT+2OA3OGrUsl6qPsP3hukThv1Rdg
kXHLRrF9h8EkXpn2S/lCerFcO1NA82FYuk9wAXqa8Ex6qU+jV0AxVLkkjsOXE4cDG+gsMbdA3Qpq
qMyFACJriLzG/CKfnpG1oytd8555EGOIXhRTUdpxuBTB/mgkYmFJ5cVAz3pVFCa63K8fJ0OVDZvV
m6dI776yT3cj1M43f9UycHKgeof0HV8tbBK3Zgqjx96/W446F2miOQ7Xuc7NqaM7nUYJgNGDgXDa
elpyH6H6ZiQhszjHk1n7CtxJUXgNxF4oa78oMDkmlUQ3UtID6gBlkyd6XuuvSKbe2n53CdAO43mf
mqur0MJSjr5FvpipjK9+BacWPdnc4nhi/gOwM/gJHGW7BH8FxlcZ0a/2A8A3rYO3RDcFrtwbxl++
qscQieN1RiCC9TljGs7rm7/f84EcvkPrB+WTJAoov8vpiVdYRGoOKUu9Z1t0WFSx7SrcPJAJwplS
7bP9bcs+LYAu/POphJH0kmQhCpYouzreiEDxss3vu37g4u0aORMkEpCeHW2+n6/Q8OqmK8RN1gRR
H6KQnTL68i+NvkKki/V1qe87561FELvXo2FFY16JwmFyXHVbNSuEkxVL8UinMk8FYXmzv7Op2P4r
hHldqcj2TDPoR0eOSLAx397UAaCOVhVdZ02I16MS9up02J7cfxcdLpi0656Ot2dd7miyXdNz89Ql
6+leTv4WgzEuGqUwezN8rtmuAldxgPQGaZdsdjZi7X6s0Cbwl0EEOzA3kubQnK6ypWIhoxzuW7Io
CAC3YC8BeSTU3YhX2DivzTCfRNqMQFlvrfoI91oYtefZ+8kmJWmuv43MG4CQnvdnzHZ8gNeffl4B
CuXJuVp6XYD5sJjp11L8hpcG76KjIIx/aOkEEDKKTslvxqXPVBEGAoh/gAurSMau+DQ7uuEN14so
fFS7Hsl2Zt32p+icNcKDN+XM6LoO84WSHU6ercO+VSoTrTN6Wgd0zHP+ysH38YNuoHZQLZ9v0GPl
HCiSoYScbg6NIiFWFKSIuHSx7Up9InV3olb/iQeDpna1SLTi99dxIEt9hcFIOC7f1d637ObNSzLp
2jYQOEvP0PFYenkMfp8lt8UqoaGOAtWTFB325LJ3uMUxyv4HlIBAmoCZnEAVwlWP9SIv9y7LqIjY
Hb/AsJVVzIFqlTpYJa+y7tEGkhkK3jiAVQ0peXnhSMS4yZqIJ8uSVftfK2cYS0V+BMupdIUOnOpT
IuTrFD+ajWHErmGUTyuNF5bDDpuw2bmHCuuRDy51db/23SKqsSFJHELuUWPKliHAEwMrh8H/M4/C
nMsAaKg95EI2+aMYTG6O2NosWGpUs8xUnMfRvzHKKpWLs0few61VPWEylLRTfexyeIXQi62ay7oT
HiQ388sMP+Mdz6HM3ZdvKIhZrRc3DB6M6xq32xwZGjObw/JMZtoZOJSdRyzOo5XelmgMyR8T8cQN
bnGpFmyIC+FQDi2Ypn0K18nvbODV7vDV/t3guTkYAT2qc8L4dAzL3HJ1lmqgUfFG8TEk1gDNEd8H
K/fVMHRZbpHzwbjK3rrQ2IWQ+nnBqC6OSOcFf2hN3TwsCw3V4OUuA1kLW5OVHslFB0cRWoxZTikB
BtbpQuCuij7aAhAl0/yB/qUBEsfwKhNIhULL9MWefmRiu0uhBASlIzt0tKD73bGr5nvbG8BSjP0F
4jQJhpCkxPves4dra8M4gMjwJR+erShtfIEc4Bu/55YlncZIJk2BsIn9EpnuJrrplqajudMEHR3R
qWYGq7scCfKhjDXdmgCrEwu8YdtmUtDG/p7B13nWpD4KlVWOhDUhjcpb/NXCA+bBg9cAu31B3/+p
p4GaWEK61lv8Se/UWnsu7ABQZr72oyiwZHPuy7rDd7NPkh2b7zUb8h7SOmepZmyxrfqHbkY5DBOS
fQ2ENQ8bnGV8mvDSoL8hxmgr63SUz4BqcyCqfJ9aU5IYOwEP2VzNBCERGBVZBySij3/fGgABtUyg
dbo0+HS7pkXWJF2jdFc2x8sIw5kBsWjXTA1PFHYULksCvSG4Akb5z5FwH5S8G0CnrifDGKD8rEoR
3YMAZ9OSbZ0J3km7lsO8qg+gYHWja9tlxu8iSqG4ZEp04aoIh3gReivdEIRANRnoOyhOqiZg0/dt
crCATX0ROkFw74iiI9S9vzrD7WsaBO3dkxOdR6zJ/OnoX50oyAu2q9DUQ5kL8A6rq5kEZ19a/ELd
JUUd3IQTdHQjcKtmiuAXMbGXv+IvPj734qJAia6ZGPAnzJ3iyB4PLO7nGMQLY4GL0y/OX3bLFX+9
4uGSPFxMp8WKS2Lo0WQHghYGAhQd4nVdblXrytzwWA1KEYo5l8Nd0+yCwm4vvVL4ssgNEnPMESFE
TyONGapA7EwKJtdovUZnsYdyABIAMrMTG1FsJj32guWW8fsbxyZGkhrSvhg2n2IdqJ01SemPkaYz
nh9OIFkLDe+vcflRCNIjJ3zD/l7NZDqGRgO4f+eL3rJgBxyOCKuveBnYW4/2leKMHkUqOmWq2mem
78NRn+WMWPNnuhUcPTVFj3Ih33qPIHgFkDMb1j1aNIW2Vf5UWTNgtcxyBjxLtXDr3JGdk6uefIs4
RHm078KiUYOeAEU7oBM4j1i4HH2ulzh6itbXZbgGc/V2XsiK4Rm2DG7hka7LGGkXj1UiXCycpD/E
4K91z9ri0B2/euAAmLdDx4wuC2Po1OCgCMlAXhifR8syeOsyi3Ozoyq22/JkCoIEaOlxQQVstVvI
bYdZNo5yg0C7RchuJEFqMvpL1JugazrCNluNkw3Di16iu9r38GGjfX8GbLjQ7rvgJtlg6IaxihFN
5fQvrmw+WCd4fHdijIa0XO0W8i6qFBRsMtNwP/2a39OkLXXHZkWRn5t+XDynSQURy77bMXm+9xC6
E+JR58sAAqQ1pxXFsdZo3VWXXgIFG0539CRb9uvpuzfdhFsgmjavKVp71jO/oKPzs+OLtBXIlHyi
W8H/61clG0H2r5G6lCQEE+Xz0p02gvdZmag+WzKHg1eiv+VXYhQNU1v52o9HAqqDy5vB6LK5e6SU
NX33pstqPtkKT6eZG3uce1R+NsQ6xLUKqGvtnjioAu//QNyjnzkufB/ihH8OsxIyv/6Fg1B3bgo6
KVJcCFphpBflnVmcK68otep7T/MpydBXSLMO2EGPrOkrw+v+7N7P2ygPkiX4NetpgRlm/jQ+NNhZ
5Lt+K3/KVQp4Ay+hH4fSmRbhCp20QKc0nNDcmzpDVMUBQyz8DHqL5m/eIkyya1emvYTJ1ILm4ure
7zYeMrfX+Td/G50RA3+Y5ZKOgOCbh1S4ISXnBB+IacgBQW+wHhr9YS254KDwswsbcTugVMUvbbbz
YxXSr++LuumsPL6jXXBWhamNJ56zD0Y7a8tNfV6wlCJPK8xJzThRtOi21/yUTr42wvvuG79QImbb
UXRiM04g3t7x4qwIQzWX3DGaFouwj9W2GtOgHzcNtDT33AvrmCm7Kn38HL8KLeXjvRm2ZGAMJ9ph
gxIi1hiwRbJK3GLuIEfQw7BQz+2a2gUGFhkLw3pV4218tFk+RIalibW78bRn2X9OC7shhEcwoLAY
8Znp2nwE1v93Bx+cyvoIytksA9THOBTV61GpagagJZIAU2H705peX+g+jk11/LY3A+6zjOE34AJo
3d9dCCf14tHkhWlq+v4/iJLD1KGNdX464GyTi/btihp7GrqityhB4Plv8UkgxkXx2Ti+1CHyxG6n
hFIw2JAXkR2OPlUpfm5W8IiZSzzhllYUMp57ztcKnmnlyYI6nqyZkWfHC0CF1X94tz6rWjJexfx6
8nY+Z61YygC51CS4CA16GuAWNjDs5i1tJPL4OP71WIL867bSgxHgAHGF+EwKV72O5lDi7wLM7P/r
H+1Rt0DRUfXdLPcXe4HsdmO1fknulT7Sysw5kACOy8cskl8mtWIylVY7mf+xNZIlltMXPyrF59pd
fbk40k9ijIPj4T1mEdsSCecYREqbRCa2/dEoyfBxlka1kJIienaDR8+mfUC0QlSMUDu4mX0xOFNx
z8Ggfh5Bk8OQ3nOJyP1aSDpNL7w3+1FGJk5TY6KkA2kBXZEo+aF11Gd9TT2XyejSeip6gt1CZLaw
tFuz9mrqj8hsgsM9IW0FbS1dX4BCGD/frqqZ3HMCigtmEWghxwMqf09kTh4FNRSGCYqFHHmoLxkV
hkFG+xS+reT2qC3/2ihU6TaALqmKg7eZgEfQjTVX1ORg7kOpBMET/Sz9fGnSA+zdNzcgz7YEm69v
08nu5iuRZDQ6ouPgc7KROuR9iSoQ4ybMEN8fv0OFVNErwenLAh7MIMLnmfy7pHnsGa7h9T5RobzG
hgmJNdQQGppNeohNQ2K6SwCCn1cg7FbTdWqJ5Npnpm2MsVCX62Jtj+Idon3R++NE65es4AxM/VcE
6Nv2j/1VHeRlFArUo9IlaIP0F+9+8Dt8c19qR19RPJu8/W7bUKTe5DAMfkyM9LtJB0e/3Pb5I8gJ
VEMg7EZEdf2OIM51UYvJJpsyCrXv1XIUMgp4aUS5+1vou0Psz3kjoiJ0aEMkzqZpL0sBUrpxWq58
V08UdqjgUeYaR5/TMJNhQRTapQgBAxcbsrx/ExQbgSUIniyLpsasiIHU5/XlSJs3UsgkCAhW6IxR
dDcJcNdM5uMsZhBkWaAdiZm9I+Pb4gXlxjO2NArmnk1pHNqvdSod1Z4c1JTpP7F1h9HnnWxw1KTd
+wQjr7rq45GX7Sw10Yp5rFE7tmF765GW5w8a4c2UC4SArjAlB6jQ7CWC0W1C95IG93DkWZIA8nLD
DXYPr5xGGTNpQwv/y01/5xJRg5VhAoAOj2FT4miI69K9j3jHFCpEiDM7QvBarPVBi4jJIqjMPdJB
Buuy9xi8SzawxrHQ59MIKxHAAADgoObispmN7lDZZI2DowRbtSSX1BAnur0/0dRjSNvT9VU8eMGT
EOppZYm0PWqevUWetEGTx8FrbCbzjGF/5WpRD+WWzk7X+nNbu78gR815B3Je6yOocF5jagc+idLs
VvO0D7qRQ0KQvGXNxfcKQHM7LhFpS/rakMkFWZ7wzPRae/YUgQJrkctjAzKY9OPcGfoHGK0iFqA/
r0Ee3BiA3IbhgYo6OP//hC2RDUqokLjn+9OZMmPRrHoxfLzn44i4xDl4Yxj5nnVK9YPIXEGE2OKh
x87jdLu6R3fmVsBW7MPq9qPCP5Mz0tKKrcLjBiXIidWLJuE0018GyJmzPZ0FEaEwehCl/Edgh0YA
AE6Gv05Tyr1dwWeKOwOvkj474bDuWGhjJe6iZRjsb9rCzbMa96MfGiIR2urc9L+NBVudpf1Uohhg
DqxPX4VB99dmu6PKwWmSKAZifiQzjl9ZWuDKWdHmDITcpwZuR3Nu3Fyy5jWzoX9CB38h5Ort51g+
ohtg3RDEUFdVG+j74CJrzsosgqGA4xl8DbJynARzVeb7tN3ulok0Vxc4RtcC5dtyA9HF1EfGxbp7
aq2h0n9cXnUK9XR7ybD/Fh7NU8pxuIt5lCPWo0O5wArIJBclPhIMfoUGZCehzq8xKxPZ+BuAZXYK
7NasHl11d+HUsJsFb7JNKtx9qawGMWfwMPcdZfE5yWjZmc9vArU0e6UBZ6AOk/mw4qlQyPPxy2qs
hksiI/ekOX8TlblkmczDIgJHRu9DTMNCr7NszMTUJZYli9TmP3OU6x4iKnDl5TpOo+1tZxw0imYt
qRSS51kibW4KVxMtweQrMS9rCQiNtVF25NP9S17NpIBASaD5cA302UoLpIFift2YF+l+IO1NQgIh
Wk9a7KujWh2w9d+icYY33mpw+DfxJSVVT5g1O2ZX6t6z4t+BmGyGBP8vgXUTF9Ldiafyf/stHQXw
FGFZ2nfrxs7IVgj5bNEK8qL/UTtb5jzsNAbCsVRe+hQ2faPQR75g3b+t6NzQwGqBANPQ9rvXh1Rh
OSaHkU/4HK+3yt97mHZV8vc9zgMDTvJn7PC9dN4A09mWkEldH4DWBZLsNatVe1MoWrtvbge8765h
xyycTm6hfFePY83vYa+msF8idoJAnHtMZjT2C/zrNoIsrKc5ffVFjl3Iklc0dI8kZuICd+xte9Fo
LP+yf6sq4yY25qCykX5FseU3tJyiGKPlSL5PHftfUKP3JlNZ4QGDhEOmj8xnDSTqd5Yza1wpvsV3
99GPuW1RbNdwLlIvVAMe9F8FK2KmK2kBbO9sQMcACo55NHLxFH9m/hyi09HNxB5+ko1c0Rn1XIr+
ex0SSCImtqUaRQnvk+dZ3y0f/7/HEEazMs8xeE5CmELnxYSdbN61QaVEXdmDgORv4OjIc7M2JB99
AnA0YRcqbo1R4IPO6oFSAZzOjg5ZFJyCBLnPGujSAT/7+ig24X12KDSyON+/LtN74mTodfjYTSCg
imAUXwxzrvPHb5xDmW6pKxbhsxHPSx4/CTWfOmAsbI0mmmn9wlQ7tk5NewcK1fRQKNiGe6ODvfnV
CR7bwpDg2qZLZZU7uNCWaVgoqQMTvyB7NmT6pcJ9qcf6+QX2/hYPe2E3p6l1gyGHu4nGnZAVDxWJ
0mH79BG+v/Mf81zfd5DULopgbxi1LKp6kOf4YqCMwzoRWGa2LMN2BFtArvwmei8y92jUuE5eFytT
RI84txXII/g3J0eAyrHSYxwLpQFz/YWAB2bHRxi3uH8KnLUUp5lg1jWEmze6fLxvsVwvmxfidxh9
g0BF19/unTLKw48qt60lhTOZnDrTTCD8+NVofQlRrODo53sWF8eEU1UubtE4GBtZvA7crVB0Ct/u
MQjliiQu8ddsubtRxwJXCgaK0WloeKU1Y8xlKNLbuYu02QlnfkutQFRDUO5SBDZAzODzye+toEYO
MZDb8N9FqJoIQbPngY3YJV8bctCBEl21SSkOpT1ruCpDDHdva4yhx/sdC/LKUB5EsozNQlL+GDS9
vwJe53eZHCMpG6c+XB3hBKRTdZ6T6CGRb1guZWSxnCwNfRdqr41FPL0d/PWgonLovpQCAXseJpfy
U+MbyDyF+5/Dij8Eucg2HrZVUQ9V79a0knZO0li4UllINv2wN7U2HGm+GomNW0IahasTHQF2WL5O
Zxu25ussFjv+hx3khaVxzRSqW4R+SLNIKkwT1W1qU+R5liEnV/Jf1QJAQtIdpLcoZQUmCS7TZHcp
NaaXFaginHmAaONMz4rdpiAsw9qUbSWTqUuZlVlnGoV8Yv5VgCNzPRBsiUtxkNMT8VbdOuXpMIMq
zlKEgZk2LX2kJQWg9QDAqYkOJHomnk07Vfe334ETV+ST6/ZzsS26cSKiptucI+rmEA0WvF63MYNE
ca0jk/QsOc+zapuXNyQr3UHMLoZ0GGgVaUnNmOuweu/x2fQhWrRYxT1qa1mlgGICdsCiS9G/GUgm
vu3rgYOAI1/zi8mdRprIEvcSLWcbTmdOJb0ELZvlCoK16HyUljkPi2B2VXb2bCyulmTdFTWtzzxK
OXVqVkPHT7vTf7hyv8Q8d0u1BB/J1EePM7YlPC0DNZLv8vY08qdbbNqLPskFxsdHDOvo1V5bG6xc
MVa9Aa/OeFpef44phEeMYADWtDVyUq/ni/G675ebw0iZJR1tzNSHHmN0xMj9eGxpsgT3j4PeJExZ
mECqZazSLgeLXHdx0O27qBxVUr/m9uX5s0FormWHkIyNoD5uWpE7UiZq+qxPZ5Dd/YzdRPNcFWK7
PxDs6zy2+rqRxEi4cJtr31oMCt7OXW0hX+3I6QAixV82XiEsrCgdzMfTRMN7/wv8LLJyGwVxqRTj
AyuGjNXKHaSoDVaGsOHKF2J5fqvRilGR0jK8ldJ5hM/swsAX84OjIG6jdC8aPfkGGOLyhsH1MWMv
1feZEyZMuEmkNJp0qVrz9KcH11d8U0xryPZeapGQIuKZe+5O/P3oJ9hhSYsykBmpzLk2d7torf7n
WjdFGp84exJnEkYe/yOCIWf3ncpNtYna5xPlGGqVRTp49miSwKghV8GEgUm1ZpDnp4qmfqbCW3ZC
2p6a97gIyERKCbxsu8TdVDrUKu0SkIXeJWMRWwq+/dxh645RGfIjjM5GjH0t0n4UIuHJeyOECSZa
qSVsigwqlN330mTROYOc2F3+eIvU1w3ETz2Q///MUuPsDneMckSk4QJWfczVrmkLEzGHeVOgBcnV
9GJpjCRU92JzXdn4DcVC8rYAmhp8TzaLJZQ53dqmsIKX8OoeyL/uBvxk3prSWLGvj2Mnbt8xGygS
/xAF5ZKpcnMgthcl2voYAl/xIVMx5OuVCJmJ83xGZTO/uzDTQsjMS/n20m3fG7UjBCIGoKLW3KBg
TKlvFfHA+Dejo2TaROJSBv6RSpvXwjU85YpUvZ19KRuyu7b9c9yvRzhmTkBSHoeIWdUzzL5pGY05
CaD7kED/TVmxNCmY/rYqGf8MucYLYTMJWC1S1nw85b+WDrzgsTJSiM0ZiNMV32h1TtM7Ob1pKPHf
HxUqR1YgrsatpqyNQXahol5K1R2AC4MrwHjGOgZRkSnG4HPXQCzn/sCpriadU4044y0yzC/07oso
tHdKTOLIezgvDlPRejNZeSrSn2YuW1JZ0jLCuublXgXnHGQ1dK1cZVSJ3MbFGIf4yjKLaFDTguAU
SnZtdJVvJ4AiZGu8wqSjZ7hHuPwbE4B8dk2fpdBgHiT6owLDmWrBuGCgBJMPXCPsHZyrEOGdCXwd
/aLJju01+5e9oHVNW3+/AU1AGHGIBRxNgeR5/orl7xv3tpAocEmzdJeVrFMEtGJYjRbZo9hXzays
TNvcRg6FgiEINoaewvCMbWTnCWIeKHPTxMNj77XcXubirG1z6KNybVXoETcskfDPG8dIQcpIkJNN
BN4wF9sWY1aluEAHbllMHTJswLMsgUkYVV3WtVj20zFL+h1UED4oLghzYLtalflFItkM59n6bybN
jb/y94fYbaCgGQcyNPuu8K6ZctK/mQDVACUi1PeWQY+KTsWko5NXgOD1WdKVWFX1Tee6bE3s/XDI
EO4Ua6B5IcigDf6j1fiGTAFttOvfS2bvJ+CVM7uu3DxWD731B6QyiPaVMZiiXkCTZSDiO5boIjxw
Dc7HyakJ/3BKaUb2hWHZ1hv8rH3DiMsMlkbDdxX879S4YWG8IsDcRSXfpHEhIoXjJvKVQCcd+XR3
9M0WF26OCs/Ph5Hy/o8HlAZOX/l5qxL61TAqLQuohVxWFI3Th5Y5l7JL43vYwaKMJ6giIp46OIIG
by1HFCEBMOAGNjRefcI1+GTqibW1VrpNt6L28XQ53pYRHhXEpOIyzjLQGIpmXKv3m1NFmGCt4j6C
OGXUYHrAiLWIy/IjCFJA/diTu2YQQ3vGiSq8+ylT5udtaOZ2xKpyWzc26/4fvJzT142m95ccScQa
3I+URD9Ku5QC6NmVn1MppD4zn01AyEnYi0mFnCzC0ypvWHqUDqsU29XRwjLbaasqy5YoaujELWON
P8mnELPF7lG1/VrzVcFMGHL9wWlPslmOEl0dz1F1fyoVjvuA1AwXdRtaJF5Pap88vqPlwmpfXXvd
Apo1Y7hkk6eSyGlo4Dlsyu78ZzwNSyzePChNkqpTtEicIXIfAyLm7Rt7J96DylsnhOiaaH7pN/dy
iDjR+o22r3d175ZqTwZCJxV7M6/uNJMllNOmqPq8zdRiaZLbi03uT0/E39kifYH5LO6tMbeKjSYD
rN+dGZUPcfyG6rr//39IJu6t6j4C9+I0LvOg+/v0t823Tco79NjxZoxNgYjSPSRxNtxgT6zvo7Y8
D2Ty9uy+BZ35p/PlCcWmq7Bs02keq10Ae4tOOWD1Dhk1da97WbP4O2ECOuRG1OtTmXY8Te/GVprH
Po6ncA0IIV63rTMjdacfxOZPDTOqlHVcDRpJXq+W7ltUPd6rY8++CG1m3eQPaN4eDQYCnIT4pptW
O66LXa3xMREQGJSNm7WN8lpf9sjHM+2DnzzcX04s1kv9AE8j0dOb/Z3WPq+kooV5LAXYxNGNR1yr
O0/loG7q4WPh5/BlPGt7vgcLAzXMqRfMKPpLa5oyu5LVoi4Z/ttsJikfnaoGrGnHfOy7rMYYausb
i1N8LeMMf6S7vJZHd7lj81kvhuQ0SnORKDpQB6LHkuj265512x2jdRI6nL/jPkp87CmF4qXqzKg5
S3EoAeC8VHTlt+CrZ6ViQl/1+Kn63OrOhhGJlEwqw1JScz161z2D1KpS0hu+dNwz0Fn1H3GnpDb2
OktMgHT1n5NDS/8jdF21I43uSm/Lxcjm/XfMFug81gxjMmxTEbgBweit3JFqddfRhVL2lQ3IJkoS
zveQYUTLet7CeOn+qAO+R0lLEzRfFcCSksBmZVsctViVRX7YKYXweaxE5bZBu72FVzz1nVo2ekbA
boky/7tsfFV6Jb9nligHQLbNeiIsLvn+OEvxAMO3g+3Kc5fZnhDwBlphXdzOMlA9hS+b2gE0VW8G
HkBFWPGPDHXsPWDAEUr1dpNlE+ugLPCiOI8Mb1CRUa+Khd0BgsnD8kD1y9Qmc5Fiuf8e+DWdngh8
8NF8Has9cFoGFGsx70LojTtsXX1FteSB4tuBErconSQfLt1G4sVZVZkXSHIfZ1z9l+b7SjqPoCBD
mL5xnWc6KHq9Eh0m1cNy8APe9Es2QP0nybBvhcrJYy8q1kh8eryFC1kLR+9O77kQW719h92uLTt2
Jvqpwv/VQ79iyo3hM/NscI3wQ+AmXke+Ns1hCzKo5lX/z7FeRMFzYkXi614KFreBmJh2YakNwJqR
M92KcoEltRvgVzpXMdrP2Wx1W6vwkogilTFQZ8q2aOTLvqzXdwBESt9AiX8qBNdpM7lJjbTNE3Fz
PxNWV7OANLRcqiNFI1ABLsh2XFKBx2ohY67/2S3OZrhNCHfKc3pCRwzwHqKUufxclproHaPaxcrP
Jp/PjTAENFTA3e5ZXJ0dgnYI5mJu2Py4W1GvgNMED3owHiwHqqVqIU4JeCUAQEpOwVuWvkh2dr/A
2miBAXaj73H9AXr8LKbO/apiI9n6r9pt6bX45qUryM/W86c3I31DoUTENoKgjcLa98jZsBTEFDdF
1INkt+foD6mOTZysvj8TaGQtIki68DQVk06Gdd7eorDyblDdMioPexTelCEmoUBU07ZPzzUoAPBU
mUMpzSfwECBTslTVCq7fwIeqaLVPB2lb8T70nawM0Zto9fALL9boNo4JUqMWZW3V0X7EA5aJfK3E
mPwQKEg7dkb1IV+Pa1dXGRFwj1Gyp9zlHCQ47rjMYaHu04AWwZgESEJvC0c1sUmmQlhQf4vNBuaI
ew2zU3734vzkRnV2+Y0E2r5RBf12/iFDDwiVXmwcpm6Nc+2U5YcOjQobPbSnyBSAb5+32jtfo3zX
z9nNM9afDLBHePSOktLb4SToQ6KrGwvA7i//E0wv5hjpDqcojUeqy/CgqfRLzhiq3DyM/pX7TJH0
1r67wZZNR6JJOxlidFJHYbDtj6ilu2pKUzq6PMmLKAFkzVlnw0DCv11HDiv0X2xT1CSWmQJTFPyi
W7pIpUHXPXSSFD5iGfZIQOXK+POveb1zuaAYJSDKgPbggu5CmTsFlWolvVpKpg6axHl1BgcgnOTN
2MnqU4hbFfKDHhE+F38Fayx64CcyPFUYJu7G0TY0ID14XjcrEWb7X/rBppMt3o/PVy6gohGUnlUH
IKupMyR2PIykI8L5IS9GLp/1mWgXJhJzDI4+cHgOvZN3sLFCdoa6ZEAL8uoDm4Sw17cujq69BaLg
RZrtAgRcQ+FZuJe5RL6Od9roF7ttTLBmqNKvtVVwH6JpzalArduCoJiQ/wVlDyQDoqDbt9w97cNJ
IkQVdApiI2kc9qjXPkO9FgXwtmJtdHQukdVaxfXq4EFsfN3wh+g9Kjw6Jq7LaUHc7hmZfRybcE7g
ksO+UQQmFpns6z8WrfMzPC7bnIp9dAsVdkUgOi10KyrHDEBq1dJWimGok4xf/Dfl+P266TzYVEC3
QDbmEEYgn5zbFp0Wme8N8n36DpihWWfEVXLkOdPffUFNSyl2/2IT/vCufA6cJsEazgyDg6bUB8wP
lMYXUuUo9cPKaEfzOwC1Wm5afIjxz5CrTm71y9LMwN1JUiQzafbFfS5/iZ02YPXg4L66YBV8GhiT
0755VjfeoLD9karvWOJ5bAkc4g7jD482R9cmyzVNH1Bs10jl58Gw2benkcJ3kCIXhYlHjHEBuKE+
KRKmyzr1Pp28GPw2yq/02b9PZAZDxNfLsPhadGLIoynRtWM1+oV6ZMQ+ewCinCSF8aEiDZPy56dS
t4IIjjjiN6ouTgbhVon9oat30gNeCW1uGRglg+qzDtEuJ5/U/GNeoy158gdgRK3pLblw6D94Hf/E
gu/F6ZirSAsPg901eM2Se//RY2HdcRghjn/uZJRjgo/NPPNQsDB6Apajbta5iU8PLp0Wnb572t+l
xEqZXMaPzFDe1PIf+xrKDANk//0hdBeiEnhkhHH4o9/NRQmvSu/c0MlPKArZ7waK8ksRs6c4CLcp
mJxAuazLkV24g8KHryNipKbLSWk/9HCBSGRNYIVM06TucDTWmpjuyIaxlIUGroF+7WhNMSsgSdYa
ZRf2pHlhvevZjAs4OYTfAf2R87jCiAUktrkCWKS+YLah2OpuN7vBt3uKdr8ok4qWt6ryXWNbUuPQ
FPvb+iBFAjWkO33+fXUQGnfdwmBZXqrKajq3+m4zj3aF5PTGV5Nu605feX6fc0F48VZiZR1RYN+X
UiZZOZXp6ZNthAneOHu/Zq0ospmdujFr92/aWkKmeS1FkRNaBUI6VB+WF8/zXwApQf1h2lWqbV1A
ep5Vlh8zmsCSvLuAbv9cOQVJ8wdYv648DgMJ0IU9pqEGjZ0MlODdRoD92Vzr+3JMdYImrZG1MwF4
Wjoe4PsPs9/hsxV2GXomD+ERibABBge/zXgt4W9b3Ln/VqHxZg2GBt3qeEGG4gFisFBA1yY2Rm6U
YY6A5cQywoUs5AG8O8a5U8+FVhjW+UTXOiUknXqGOuligO0anvP8V5543dPTW1v4fKDiqICViF61
T3UAERRQJBaFZ10F78YOnt3cQxDrNY6dY5qCyeD76jTTP5C8n/7dd5OVRXVTpYBFqcYr88scMUeq
YjPGfVbMQhgE/JU/gDxEl4GK9hO7PVZ+hec56zvSFT+lOi1aWEW9zaecSyb9TMFf4+ak44J8GDu0
/Tf8EYYz1tYBiniYROWDlbRUnoub71QxJ3owzOmVq6NrvBpCDDod2TaCSGmfomOJx42HGtkeMBSI
3WjeIPHnFwnLAnQKb0q5kjLsQhw81GcwHOIeXfMDuWzA5/LwK5ggoGsOR2SGAwOHG8VkLfYnFhTG
HaRd/EeVnvPNQ6RaIBXXGoYUwR0Rew+ZpuzmkpxX1ltTl3irbTOHAuzxBdghMtMT3R+tvKz+mUV9
uk0oxNikR5uc9lQRSZbd/HFG7x3fZJGha6N/8Q0oy+X8h3SbDjoUX+7uekjh4nyuj3cv6dhNrliV
FG41IHOTM3X4rZBhFveUAG6AiOYBhnwBOf4PM0qZS7XF2AudBHECxsjs2qba5lShInBvJRcQmDFU
jn6doCRfLoscqL51u/DvccLYbfTBsBRS26zyD4XM6KDNRtKqL71HQPix3FSJzYzoztA1x8/xkjTt
s1TVjDDQ0VGsnVHgxoc4+9QD0h9rb0jTNudXn3Cm88WbyaIFeTuwyIH0lrFjfZrzGnREbiXiV9y3
3S4EzREjlXZLxJMdQCQyVx+20DbuNC/OY/vmpCW2HBEZUYzvccmBGr+UC2sz+2pNc6lXXDZ9dtot
7xWbQUiG/CdSenoYOXQxSvnZ8Wo/l6ctA17ocZ4V/wpnVL/579/H7C1Az0z/3YOccIiE0h7mSvmK
T6CQikqZPtUGtaGStV7svQDzVXF4A92chIC8Xq3m8GhPFJdpbkF75KaJ7kABCqIY3kBlkeN1uYeP
fUQmhD191nfNtmOYwnEpcWCkXsWsW5YJQq6pLUR3XVjOaeyq0i6TOs68tmP78OUeaMm43WXw5Lp7
wEJ+O6b/tq5x6ef28b+se13XMFaTk8hrQCUbw7PtFLVhks15BCfkkgV033Irg48z5/c7KBGQoEI/
kt9KEL9Mf06rni6L6JiGRY43/h0lkKfx8yyRysrBEcYCyun6h1vLefLZa7od29VfZLd1oxIp0pzp
2GZOrRLVfCFESlsWbC/N56hy/P0qYFRXKeC0P3AKksJYU0k8KLWbCBGO3mCsmlWjMMBLZ1B94nFu
CmuOiYu6cg+b9dibj1U7LgwEa0zce6vjG5LpJ7K5Fa8z8PPWAqZKY67rSYU54EVmSx4OBcJDjh1F
FoMBTTNmyq7hg4zmSJdeijW9wKy/k0TyyGfPpEvDkh4ir08TOqgDnMZttainPcFLrqjRqfMc3qGE
OYrCfyuXLsJt1X4rHW3cdw4GcrxwzM/bWNbO1vRbswzcusqQCpPX3A44HQtRSvSOERyDSwSv1Mpg
6SD1VSkJRLgabDcalbYcADgYnS6hbpT9vxPe0tfLr8T0vE71e2oObUCgoMyfmVRSU/gxXKEv+T11
SaYNvhU51Nrm/XaOqP3WuaGoLOHvfT9vE1OV07hDwzncn0ZuAgG2EdeVRXn2Qom5xAOr4UUg2gLp
uvpc/VURgOXuwKtFxM3HRqJ1fPhXkKDchLXdmut516Jxh9aBUZYqKBWyuB+2pIjcgWvbfOjM9E9s
L8Su/fArdbMyk99PXHmh8ar2/P3uL+zDr8XHRiBsGEHdJSDHFNoAQIe9vBDo+Ihqv/uUVWZLAC54
Bgd6anXYde2JqjiWAERjOIItYRvtCWFNwIXWT1UtiZrB7BcAHp4wCIfGy7po33jyqh9eLr1pMD4d
Pls4pBQawgVjagKhN8jFvmjRJEVMbjtCIn7LxO0KZ9yPYGDkVbbh2Jgg509aDbIMu316qKjgnnZT
MsRI0vHkjGZIB3Pc2UTjRW7RUkOPfrKwEiUM9KcWZ7Dq/1ibZ7sAhGMOwc4RqzIGtkME9KdCPeNO
Cy+7zcxCuV6/SZQLg3eH2Y4EG3qcY1y189GkkJrgD6rS7ZOnPOL3y22kCgXW7OI7Y657QU80sAr0
lfrl2CKhpatU6f8Wj7LoArfILsw7uOieqgglWjnoHIOhRKHkZnTgr5sEu3c6+IRvkExiyTVUl7lq
7FBHgiQKNfXhDSMR9hhihn/1cM1cdtZssupscslN0HbDxNf+ZWyDCdqs2cHROdAxHs9iT+7Yu/uh
b9hG7Li5iw8Bg3KlG8P4jqPYvdrZDMg9CTwohEplVx5lTByM9LXHx+x6OltLuva2QD6YmzVlgIiO
3BBksLV4yE+3tipoklPWdaILT2sVtxh1hMVzLkeVpBhoymzK54H5qKDZT3h1S3TkHLU0JezhpO8H
dQ0jQOE70FkE+JMXv7L3fGoLf4atKANfqOMa13BlCD+OHxjXxwRbG5CX5ztqon0l/bUFztClyQ1c
thzXgoZRNbVGGoVQLRGs5qOoQO8zzmnECsVN+1NYO37SUtiuwsuF+vJoTDRS+CyYGkREbO1vY+p4
qzHrAUIoxAcuywF5BthhxuNJGPgnV5dQJ/LLY0xHHIsEpYMVHQTYnKL+tuZSU12wWm9GV5oYKPOI
isXtWpB+ahtg4xyJo/L4KkWCnIkHFoqoMUaXtKfQm6eAdhe44NpjI20y5uRYk8kjIiqHe5JJmz9p
R+sv9iO02sDOOySrm8qnJSVdF6vl/NIrnRoaz/6/v3IJXV2mZIVet3fK3/BM4yfEqeUvL9dJQud5
3aZYSlLWQmNqFN5Y4lTPxjUQsiewOCS0CaGKPPoj5ukz94F/MYoEtybMzTk/iEMjglmVombi+Krw
TYZhfs5LZd+lQlfjpLwvi01EZzpyecW5defXcEFOtaDCkPdpTc6sEbpsDcWlntBqPXbMY2D5jTwT
JSSw2i12T9yQcJJmXeDuQ6qDn0pJ8eyeoNJva4TIIdYifXmwyiMjeVBvguSKc/L/3YcpjsgYqS+n
AEQG3C4z0SlomA3VKLRU3DDbtiaZsxxlbBMAl8ECz6T7Ipjb0G7Y7WcSl6eq8ZRfuUdtSkrjk5L5
OSWG8Ay35E2MuzXudITseTzE3NCBJ1CnKQaR7FBMxt8QkNJa/4JeUnOHDpsPGLwMraep4oGu/dR8
0ICE2+PddL6Ks/wnW9pTS0wJlmcNfBtRFYynWxHP0IrNa2P9KLRx35mdKWBxe2UYuhPBNf7EkV9H
hZdLUwVf2QhQ57PA6CIYLhomkMM4b4WzSiZEfWEkQ+4HBuivX9VFy7SjV/cE+NKsnUZh3udC12KO
ej1YkMcY5CvDu2UZat1AwIzWnmcow5lAxfjSCRKhco8LsImS+cVk4ozXjgPd2y1WKcj/KrGl51Le
ZpU1wuSL6/tnVFqM/mmB2xbruLf4K7uf9OTV9rMLjjyI53Tqku4/JwyrlST8kONw7E/nRx3WI4LO
G1kG0W0s8ybh1aZPQgeHUAMPI+mpKDxpdLLvZgP3S2WzIYDuDN7a3ztPiIfeCxddsHouQdU/DU08
qOVMTpxQmC6s0n6a7/yvZSs9NWz7EMUoYTWkebCGWZ3owf62N7kdAlS/5zMee6JiJubhPcJgQpuT
M2qEbI7Aq0lya3ALtlX3qE/o+iKLLvs9qeDamKqIMBmfw9Ai3sMge7AKxcFPgfHYg63ioRSEKnLc
iix0n/noj9G1nKKQFC9DEm2kHGmn4dQxpzb4wmyQCUwLTESoKJB66ZbG3ReBw21isgJtz1K9IQY/
xeMT2jlq1x29xWoaTyDn54aPLeeCzD73uwa++N/sQ/3yrcJtfLXFLrW9e041QElVEX19CXiFgnKG
0GvbFQ8pVxVBCc6FPfoVLrtKX23HamweitU28fj0uy7/02YUiQG2s97OuVRkEM6MMhsGvk6e0QRO
kjV3Zht5LZOmoR/UB65QpEFkOqTk8RbVMNJF1OPTUMJCjXMFHmBDbQTHnPB8ZYlZBPRd7shJFfN/
r47mjKQLD3d4yJu/k7P9t3QE481JOiq4Bh74HYs4PszGgBn/t3CzF3/DSgYAwmLYPiJrPz7QtNVw
2ITxUjuQRoHFTKVwlY266tYpBLfx20+5uj+/eJtMzSuPROxVnwKnWSeJy6DvVG3JWJ93uQULOZnA
LwRcJS2y2LTpmEX8G7u1NuTkcaYzdWsYAKsUxKiG6ZTtfxPWgEFSNzP5xo7P9URt9dmYGFpmsoq6
xwQTygSRj6iaTfJ2AxeIqK6j50kt5S+SGFryZ8Bsg9HtIlH7EM4ZYhubig9ggTYrsMVik5UscRct
uOXccByE1P5stF2bYQCFQu7oGSCyjMsDHZFcRxf2FMLzO1vX5LCy6/q5nUZY3vEJZMxD7u79i5yl
IsBhoiyvvhT11mzhUsCqB/s6BeIewV3yK3D3Nx92/r4MfyWwiNvz9/wwTL/6S9O3nlpT7X5ExsDg
aI6oltOiTPqP6IqAQSDPNCh8ZM5PtgzlrSGwPQgmW/LeObaMyEsKyHAj8+iXzu9n8f34NwExvdno
EieRdTibNtlGqLcC2iXwiMNhWp+5Oe/dF0Ij0kJJ7yLAKTjMaqpAAx0ETDY6N+w4VgNlmGYertB9
rabiR2zBBKrqtBJaCRmSvIR3iIew7HtaTNAWXYo4LnbrCMnO56GMLRxvVDLpyKq0guAG3duJbFM6
IfoEvg6u1rpeEID7WzjvyWdzr3HqlL9oo1otvQvZ3KsuHDzOxH/03f2fkjk2i1bkp39WHNuTtbWM
b26Ponr1l1OUiJ6QnBCMQbdkHKuIhpb6MmYiprpdbCMhdTy13Q+c0+Yk/dZKkWe6Fh2vpPum+Evg
x69zXb9QuQUwSB7zaVAi4N/8NooW5Hn9RjUsp02zqp0EoD+7QxL3AgGySLVGnKtbkknsOvmCi03g
wz1BskmtUursC1Cgmg/W0ZtRipZeXOsjg+PoFX1pf/WeXVHbO2qNpuFpmrpSkEMnxykTfKEAzGPU
8395ZyY87MQUfD3ABCheEwgud2LCOAkLxhAQe+yfC+F4Ufzx4Ebz3HqauQLE472YgxDheCnIDTeu
JbaXQnGR0/Iubm8vwiR1rCdTV9MhbkqK90/YCiXvuuyiI0xm/JV6lcLU2g6mpRw/mqhHV2trURHB
XywuelK1u4aHCFSCLc19LEvOqj0y2qgt5a/P4zzG24AK+djJ5Urm4ICCfBNMwL9YwC2k2eCnplw5
A0UgPE3pMkjpmceqzpilba8KpJJVsFUbkEeCYQl9oEgU8h78IpdojtTfpeQ+09xeAtQhFBdEkTzX
kkmDgNVqb/Ifka43PSUdGi4MEkXJmUiKNxDJ1sZffYNoJM7cQWeWH3u6IvZbhznVyfT0iG56Hic1
otQoY87PrvJxS4YJT6ZAEhCHY73o7M3+Val2fRxilgUjhfHJfFQpUiEu6C2TlJh1ZwK4Z9m21w/d
yKYrY12WDD40F5Jcf6RhOs1SvVieXo1iv1PupB4jCS5S2FwYaBR2m6dKjyqczwk9MkG0F2YbhtVF
xnwryX8qXrBwd8EmAzKbwLwGHMK63RMfBvCQS95re6YvlW+boMkQ/OZ+7TPeehC+d0n0yWiDpEYs
0EDIYSsO5t/lld7YW7Ag73iCcp6IgwpFCftUfAO8wx01RQCVhEFikVPdl3ba1YLLvXYxJVNKyA84
HAn84SR0k2bZ8Oi+zn8biUOAgl5XK4QQPCFdUUEq9S2vcRIL10JMvo/GOR2X8DNjc0ahJlKnKI9Q
BSSLGSh55n+wZaMDy9EeOUKv0U8MS6nMR9auU6bRzI5jW+RWVVd6EUFctk5SmC4g+FQgSujXxhCm
IlquDZrpzuYNVXXECNeVg1JIMKMWlCWHBo/t9ZKYWJYgTkFMRtg9ZOadmHjYVq6hH4f3fMkwZnsf
NOQkLLkg7iRidDdJNpLyQnUq7jeGHgNQw+x6l1ZFfuZ41H0f1kInYcgBFoN/aoV/9a+y5ZURe8sL
pqRc+5ZOtplkizljSn936pcnWqk+Af9bNAsNmWJB7euV27QT1CwsZmmU6U7zgK36lew4gasaVKt3
mcKhQZfb9y7BsbWez3EjSdQflMU0uzDcb9d66SltnHoTPbnBbUWUl6mL8JksxqpIXY2zLt7wCnVJ
z8aLc0wKbCpgklRYKcrjKTahG6bzKvVKJzwYbGWQ+BmQnt7xf5ns6rn/TuJKU69kTjsaWU4z9OFB
uW1MsiFq3F1D7ZzIFngJbRMLxLhpRdIKVdTZRiY9YOWsIl3aFHY762bTapS8S0V+B97+GbDtwPLu
UNgdW341NmuO7mdQAFGYDr0k11BLjGZdFrrq9/eEDLWCOGC3l7DE0ITugX+7H6kMoiIJuQEgJFcS
PToUe7i0bc72Xe/hzhFq8E5H7uLdnN0pAWzq5DNENKCbODhDxjt2RNhEPg1nwudrgkTX4PLU6vYT
o9AJ3cak9oS7YBW99FyE4THt8DazEP8OE3fDZ4AJUKObSF2+gUazLr2wVRHQymfO/iBTdkfbWjlA
CDWGa2Fy0JfVLCelNf/ERJF7P/z2dn4ZSOoKKQ37P3jg7ZRaeT8NY4OM8mfL0b0UvcDSB/UljE5B
GMIprtE3vYuZZiYm+V/nfeyULHLvxdjEncCTxelaWZU8Gl8fFds56sGHQbxgibkmJiqcDrY22whY
VndSaQVQpt0MhbxqyNgG6gG9Mv9OxyZIkCs3j601ZBDFDpHV4ztuGG9ZvpTLjLTtfmB9jtNhIL5v
Z3uID/qZh8p0PeqDVcp/x+7P0KOcDFG8MvjEdPeGS6yftGjMnRQQqQtJAh1zTk5Ie6zHgcPoyfWc
PyH35Kk1VWlD7E3WQ9ZAP8DwbDj4DtRKJ/Yq3DfqZouOPL5MRXQG0Ge0rkWn1nCBM7XyfYPbpEVv
1X0PIqffO8kal03nqa10/qv41GwwddHbjmytOKDDHGyUk8IGU+Me1+C9bjsOFuLX7Vms1H8CpK0U
BafE5mQ3YRbD5czgxt2Y8btL7oYSH4EfixWUWXJL+cIp406YNL+fAzdITxcPXTinrFPLza5cJb6k
Jx09mIYiSlO75I+zB33cQcSXmZoRpxltlo2Zi/SWfkk86QIsKkh0WmKGDhC2Q+uZg9QALr2lt85K
oVZX55RODWNhneTzBbFLxtwQtBQY5HZYJ0shBWVZxAK65y8usHxeP2F5ZJwwHpunlUgv8NBQZvwO
YxQGJxfoBzRrdJmeSRhaqbyWQfwEZO6fVuaPtVMQ0zDH3cASKiq+lfJYm14lwNz4ORqX9GM0NQFv
eeXy251g+5iGFwcAILQvKiKEzqpSrkGjfwUTCQOpGWbCGZYvDyASw3iaXHcBIc/bhTxyLUpzs1iu
3lwGTFDJMUo8RkXbiM9bu/I7iwR+F4sY8OfzEqlznS2r0iFsoN1DugU6QnDFL5HQ6qtzGEYQXsnB
UkDwrchQeGYqVN0g5C61ByBW8XDwEDCd3UstGu/pdDeSXy4jmeqCC+xvyDxl8Fk0Qrs5//V584a8
hziB7FH9uTPnUsW4RtkHeKGv3V2jeT3QUR1RAv8RGug2Y3Acf69SFyGUxF+lnKk1M+a1e80DQl3T
Weyf8OkfXfUeVE9aUD6TWhMbXBFeTd1GSHqAk0oCofFT2QxRPE76WJSVPUdBbScDqY8DGONGuqGs
AZ3g41Lw11z2t6keQs80brXAwI2+o71IIbzc3cXE3uA+yVYjRnOFYw+Lo8EaCw7OI1cqSLrIDEUr
LJB+bqErKo+bMll9gWcMN9yvwTWd9RyY5KPHMLFJU5rUhoPm5IOWXx90u6qW8nk0AHhI5evOSiBL
oXDOe7sJaeIi737YkdM3HaXM4+7cWOuW0LYOeXF1rQpdsAtIrYkDhCEHkByB1r9zTDfWwXcpNWgL
SKcoT/7O6JxOgw8agQ3fiQrx6kdWrq3rKtaDA67ic7K2w4CbMFKuNF2YUBYi6dG/8osp2/RYoHT0
4SdgG2jGtT0hnb7Hs1qKhH02Ci2dHLQN/tLJk8KsxmXh/pvZuYo1WvK7naV4Y+pCf2CffhOmGYgH
Wt0RJ+iOg1mDDA+KeVAxcN2/vhSwe+vlkJYOBnG3L2SRROZ4s/JMDRFaN6ISymnr31gn173bKYsM
jGJ9EFw8HWpBZNUJMmvQpvM5F1FNrnFaxSrn++LLm4eD1LtLgkCxCDV98i3fYfhumxgMQW6T/i8v
0FeGRtUSfyWkh+woocHfnpnzGYTZ9mvSkMfRgn5eGBSA1Iz4ICaw1BjXk7utcAtIKQkNcO/nJKou
xHKXJ+LRLD8EX1f46IdMIEjaq/2kNVTMAx+jVHcGBYqTvBZuZ/4nAC5qcZU0k0R/qNDGg5MmKcRp
7MG55/HnlUXTk+IapHlxVxQQ91GpwEjYfEgGh/Co89hooy5dZ3ty1jWwsvP2+KCqjpBZApPYw7uE
IlzdbVhf3U978lFXzXA3hDZPAiJ9xJdzGzLGggnAeDzwkzLXWHO4gf1OHyOfRVw9iWm3X1ykCaNX
hMCijiUGnvePDqY93cvm2rzqkwEbbm9w++4Qt6sbdcT7cs6qAwV4QWvCjhyZ8LLHUpaPJ0YzCueE
eQ4O0ZLhj+4Rz4lDrBCazqfnUBjtpN2v+HjZ2t1L/fHLw5PC15UVCGt0p2vfo9gzqIPrmnyd0KWB
XecR6yg9PjoE8RI0XApM4cblnLb/NHmusYYVwCzi8/3S2Bk+hNaAeV7Xf0cT/1h6cKr9yHElB5AK
gUn+e3S4ERWlDqtavRuttpWyTr9rpDaacffeQ+dCX2o2AMeadgzL7h+hEOhT/iDwhpx+oaHc0sy4
wVW7rvIQHMyEynherkJ9b5uDYpe7no4Ek5GMw26xuX+ElCnKrdnQ8U7uwJ49BWayVv5XqVKLsWO0
MOqxthYG4l+0nMtn2lUIDBDjB9hgof+Jy8GxsDFn+S+12JlMBUHWUse+HfQJWwdCn+qM/mIbmd6+
eGY9GyHNxfpqxXMSrIxF3QhJZOpqrL/HsAXNeuvET/Cu8/Bvps8CmmZB+CpOOKlV9DAxDumnsw3r
r2EDiJEPUfCU2wV6jcDXM4giCcGGWqVeeu9r6ce3qcGtvDJ7Euefss5pUFvbPq13idpY0j7TwB0T
P0vN87Q39zEeoXo6e6H9QsLG5TbOoV6LKD0GveSdrM5ZjE+CXGICriRaPjDXF18aygjkQMk8/d1C
ayBz7KrKVaSK56uIEgJgr/i40njlzItnvK/M1MrYF+hYjzUvS9VoblYq4PkhSEV3dRCtrP7BaVfr
SpwC84mtWpIAEh0Ys0LGw1omToFBnsEAFfqkVPSIpmh8fd1AzmdzjLUGjJ/hbv653adwzG8uZFKo
1vHY/uUPdWY3ZQ3paKxeEwrs4qfK4GHfN/mrhBtnYy9Oi9+6mSrTO+8k6FWVw6+vNMeVue9H78fM
4QHOjjj7g5y5QZx6Wk9tThAQ84dT71mpp6u1jY6uxaJtWFSHxUdvGvCBoieEX70oit63Ylw3n/BA
PRgKk+jYz+SXPAy3kvg5tjsIix2zkDr2umEq05IjSI/rkRPxlXnoJAtXCCrHt72MOQRO25FsTAcU
N3jfJ1k+EH3FJUuClbJ3wepgY3KAx5mYR9QIuxdVDd63o+52li/gJTFz74hjOvBeWTPXyIa7VpE6
uYNxztkfSNUf4TYaN5AuDFestAE+8GvMpbAnurvC0Ro7ZVYgKHn2av8RyL4Y1LbgIrVXJlIRR2WZ
yXgyv4mzSgkMwio22XA5gQ+2NWQ0e5xYqxTM6t5NgGXJjULJWKfCQEGcheeCl/VX7Vezvj37vDVI
Sxra/ofc1i+q1l/tyNVvESA5vnEiQeS/niHEDjwYfSSyeuk5UePjSqiKHk3p4FU8b+5JlN57Y536
wBdSMxcqpv7s0t3vpmowYFhuWPLdQofiCY+Ti4DKd0ita6dpU4LYTl8fXWXKeLDQCR0/FsR8aom3
eUnLjd1e1GtKNtxhI28M/qQGn4HGy0LrW1KJ3Sl9fsp6UhyxAVZnnvbWuqiqDNq6rHgbfWfYf+QC
tlZrjM53jVqhspTvEzDFn9xI3AJtOpb70MwqrJTyWaVlx4y034XTLrPWfeeWCtaSOC61Q385p5w5
y8KBc+1d8UMt3eobny4dXgjalWquWb6XsFjt75zPM7GOltNTTwT0dzwls0Bxlr74NCiuWZKLrJXa
cW9ohgFxYvZxb+6gbktMm4GcTtNBn6312n/4bH3tojKD/m4H9xzvnfWmrXvUgdlDo2NirAwuclSn
1kLtwohvt8wCF2prBYRptLLG2t0DVF082DJG9Uv5qSaS9HD8jmpkQjRMiNY2YJ7DdARFfV1agrRy
awwSH8AiOmuQcfYzS7nXwH+4j/1uKSPVQXd3YoCy5yetBDiTZj5k9N1gUIUd0zvlx+2PN2Int+ge
G1tqQM36Cl7vnye4+DZ7PiR2OwLMsgCRqti59/7utVgaw8ND8wQjMsFt+LZCpeKQUuamoEwwc0Er
fXaLKVctvBTonkwmhqhfR0ZC/a0+1xL/QAc9mXKZR9EHnSKf6pkhLuwn//tZjca8YvikeTi+8Suo
OlC1nBOOPeJ+V3YD08NmrUENYmD2LjCIeKnNXXOAiQLYfTEhaRF2dHMAwd9ugoYT0PV8lMvGJxWC
7M2raZf7++lubEQCrtnFV52cnP7wKUbvikxLI/4foOmk/J7wpz8PxsPgrULo7/COo734sqHvoZMm
cYij/vlUfYK99ThKoLh3HHbyhe5K2cjb2UMp6NNOsStbzWgAN5UZydukvq+zpGuAbglKzq1DZuR1
RpbTreq9GAHXoluuAYBwnz9zbK6cfDyylwjhxq9f5LqXbq4HQokVeLxDwz7s1lBVDBMs1qpN+Lsw
quMNg1FrYbGzPUliKLbuh21bVbryrZAO5nGgVbE++Phb4iU3uaL/fQZkXNT3XwlncgY8r9TBdQoU
GYJlyAfjml7fkuUq7ykVLrKLjGrYViZjxArh3SqA/FLFhl1ISV5fFsIUNI/oNCsHKOofOvYagsv4
CShpfbc26NCw2M42LnsK5HkrbJce/1t4YUots3uPI/Uwm4P1vJfN/89xihFAuL5GU/McxYO5VQ76
aEV1fiCzV/m5BbCWOiojRpIkSFyMjMmhc8GgLEPE7TcjovQ8MVvKzNCxiUExOkK60Pey7ix6ijuN
131nn+bZZ5Q7wfoANUz/lxh5XSthsL1OFxK9Y/Fdj2SQMMn51PN2gXY4OBnTJ8v/M6j7BBJRkatP
xyIoy8UkAfI2Qr0MhAkg7VHk3hQrkzUDXuQGl7/nhTefR+REz2N6Ts/+XU0U/HmO2Rp7wyiwmggv
LeoYoakNUnk7yh/00xvfFYO53uaMyap2bhS8HFJQ0DkX1WkbstbwEOwe536m7W0D2BSM8Q34fMts
V8ZbaHUesOKVSYCWFWKg1mdj6ROYewP6upK+E4R0tuG7KzNA1mPcR2JW6k+nueKOWYlMqJVcMOkj
KIiF8hA3dXJ0e2jIS4wpeoExkb57dS+SnlQe1JjwH5+cMHLDAjsXbh9tykbb2JF6gOr7Rf5lbHvD
ppXVNA9Yt/kWUE4GZWSuGwsNi6z6lg/RgovRxwseFH/MWr64xwErBen7rUkGzMLwaLOO/MaICfMK
v9qXw6c5BL/y5BV6h//SALyOTUcFNw3Z0JUpa6O0FiVXnczDwB+GnCXKDsbpl5xFrF2X//Y6hoED
bwEVA89ufZfv+xTnpZ1naWp3dJsjLsxVNVr1b6HhclvOp5drwMS0nSg7e7ZjvI2lZrCRYJgrimro
Sn+0Yu9U3P0gnpBZNiaR/m0qA5C9pgBMewK0a2rCfVAtMbtApC7UfU0eH0WZkP60mlWC+g0BXByl
4y71MZgoHU0KgrBy3mJbfXfMCFQO32yvIuilWd/qyM0jlWpcOTKsnBdLncfE4IBtWuUz69bO4F3+
r9ZeLYw3JenhoM0lR5P1BURv4QxDiG5Cee7VWiVc32sC5F260DjVeVY4+yssOYRd1BYtu1ki71Sj
+vK/jnQPodQeq8wPSVeEgRTjRKfe4M6phDkf6E1fa0mFoKZLZpBke6fefJjepSubGg0lqObO39KS
SJU7PfiD4zGgupaoy06vG49DEFFZKcGFNuWEu1x8pSRwsJ8cmd7a0/Wunm8v0D9DtMM1S1PnlrTe
lo8UmHHROqI+24DlONNWTQh8nAWjbYXQXBwPC9yOcG2sxGSA7Dhz+ARLi0gaQiXlsPDf2+iuGULQ
c+rjVc4u09xAFancfGVYN77KmGOfnBvQc++Tne2KYzJztJVl2jqi41LkzTV7fdnm5IFWQNMSdjHS
3ovnfaJDaas+5KEr+oX4ZL3URMuDbxvO5eb45qDqpg1puuDn7uiZXB4Kn2VwEmFSOKD1GZLTEukz
aA0nBpgS2kI6OEwKYRlTwvkTynYwNntfFiy0BTOMyRJLzTmYIwxu9b1vQH6/YFBpexOPrWjpOYq7
0L4WjUZtM/roPJxJLWYftxXud9fk6rJ+a4v9d2k6HpuC40WpjVjUKm9ADxOCz0JufzEuuSH0p6ny
1vutjf0o7Y3uk+J/NEAA3BVWKVBPGwJur+IuCLcTFMGtjtw1sq1w6dYp+aLl8kQcJvywoCxQh5Hg
C9ghiaRyl7JF6O0h1k+TKIimt++xbiLyVSNL1ZSFethjpnN1bAMXuRAShDK2f6lSS8+tHmLG+IBp
KnAEi+huvax+F/na8CUqBvjsqnHK7lidoQci//cqBXV8HHjzbMcut4VOmECIUM1cObbDt9NMlHDA
tgzVMQRrF7FxRRgo4R+9lfB8KYcCUXMId4z/7l1MvGzU8oQ0ecZWCmSO7ZIyP9c2qijTesOOzErj
3tPcZqR/hY4Gt5VO40ER7kDacpCF+yWazp9B0ZaqILa05A+buNck3eu/o0/UOP1Cd4R0UxL57lBO
m3G790IBtB+zIt9dWgVsxoGcI/cFz/Z40NLoq8GyI2N1AJ8PGsFOkZ9BJtn3DQfRswB+BjKHVqzH
W8qKRAO88q/sApV3hospyNu1AnhYM45gQxvRoxq9k3517BNFSggR4MQG2RBKTGm6GomrDOgk0uOS
nsVaRTjtVA2V4XF7yGXb6Vji2nBr7xLdW33uIz28DiQX5YvRO7JnYPvZBc+uVu835j8Q7slgUd3E
qB4kNOP93HbkqKTm2SZSDdTMrFE+qWL98ltqMtOBlQjZifI+V62Vreleqzdg9LHDIpHJuJkyBK+K
9T9aCXQOtyjCZIkceX5TAqSCkerOfCx49d0zSQQInp/mjiKi1uzeX6UW3XSQdXDkisczmGfUDRx7
Z0KANxCxD9UfrU1e4NyBn6lbNhsj3yIen9ixFi3KidHVn/SyJPFGvfTOQTGEu2WN2Sg8GHDyJup6
oyAwZWaiGqgLU9xRFGAph0tVPONBuT1LZAgq8Um3PCW/sJbtvBN/ximdpRN6D6OuPh55raDpn+vU
KUK7p8vnIwVq0/9XhAastGLDvlJAz+jDVCcwskJYhSyypsonKXWB+kYCqu0FNYuOz+//zYcOt6du
g6OmN06mrORlWhRfyhCARy1RFcFsAxI4u1aSfiR++3mUB9hfYCAfY8fn2HEiBlephAkjHCpa2rx9
/Gzh9sBEN45H9sWePhdkHOzbtUhOxx6EfY0mDWKC52uWpQIrOdNtyNt14uq7T6cDqFAS5xU+uyP8
wbLsIw408lLGhf3fvpydQ1xsMyWa1Yv97gY3EsZV33PyM/a+TRQmo1ajfOPVuCthcn0Tps0L0PBK
ELI+jp001GqcrVp9IR6sH7UhNF1U8rBBqIyO/P1JYFb7aAiXiX83Pih8zxZS8ZCxaStJrRYUF61z
mi98EsrX1O8B5K4VBuaWbnWRKZl5JPI5FqQnHnpJUTEzAWFq0lYnb9cauHVf2OuAY4Hzw6OLFHPG
yPLcdYjtHVkeYOXJH1al8R3Sx2k8CjQO+zFIHpkbnfRfOg+FFinuuGYwDlJ94ZhlHgHIxI1Sb6c9
TpdhYHnr54/DQo2CfTxfA7xaDbot+4EeC0EiiItqXSoM/4K3aEBeEP5Lolkr499h88+RHSma3C5n
6rLQ5f9g5nmxHE4b+FnUfGkeVJrPlhpOZUve33fJdkbv4UkfBAIMJ6wj77ADWlTOgByEl4CrYSGf
vLIkzm3hgbDdHro/qpN5KQhw/DENB/NdQqwWM++cr/zHTA+ut/0OFQs+qFusZX4GG9Hx0Lmpn1+c
GhP/6Z/X7CyTPAQbX3uXk6EySzHwzEvmpyCZ14gwN2hsZlGm0J2dIW1fh+Bq8my0hDmmGhwvZuqG
VbPN7G8AH58ZAJ3s2BU506ffGd6594wWJfNoZGa/v6UhJ3sXbf6+/b4/rxwMZoHElDwSbVmbzQXx
ghBnkyEHLPyz+UBUbRH6hnsNCj6Lg3dUbls8BpI28MT3fUy6VVfa4Ipjh3EgEtAjrEX91CtIlA3y
Jp/9Hlj9yz3gMRE0er1oWoTdWC3RU49E82UyieJKdH3XxyMXpgvF+nc0w8CS/Vh+QM8IzZa2RgS3
2HAU6n0pSyZhNJkgmTQ9Szn1K2SrrL9Swos/6Ee7PA92MXf0cBhw30+K3iGwoUugNCmM1iuMVReP
t6X6RBFxyiXiTZ6LdXMMKO2tzpiHgBbgQn2OHZnCz5zh/InvP9dFYip34wsHiznND43+TjAsxm0G
f3sm7/vtanbzJRYGLXWRAbkvSJurvFeNaOcxvjTtomV40t9KAYqVVVVUhyuy9bIU1w9lFoEQCvHA
iitMJIkpzf63X5UsaYI8dPoluTZqoykjhvKIa6Mg7Rt2zBIL5Q2pmQuPwvGyMtJqqYD7w05xF63h
3AlzNH3UHN75OMu8httrEABhcrKJCIRj4l1jYxcMVldpULlK50ib483MfSN2paJfcz8UL50wjoUZ
NTQBUih0P/raxlAXsVnvU83u7fTCOml5WN2nRZ4zIfAa6bjv7/w4Qgbe4PxeE9aLImQc/g0nZHjb
zvBolD1yxIGPtIMPBzAKv2qeP+nRXcE6OABlETme+V5LbwaIkTL6sfYuZ+YHbBPowLbPMdaz3ryX
WWpcNcXerke//uZnLndNqIDFPmfdoY55HW41ckpXcM/nLm+8wK5+vgupOzSaSiLNIALbesYnsa9D
8dQegd0Npfj51hOhpLyDZZWMh5RGzluNOL9bePzleEksiPEfEYB7B22NPL+sfeYWCyvq2p27iDll
1hqcIKbnW0Yu7F+ESoDIw7AT/dox93SlFrQcVPqs0SiC7tMQHTGJeL3zv4Cx+U6Ulv0HFZ0ebDow
sQxViUuwOgpIvXS5d2LikipEyu0aGvswEu0cgAnkUwbI6136HrBkcogiSjHVAJ6JXMncSzBizJMr
B7d8kKua7oDuWEJAk8cc7cqS3urYihaMH22YF6/vVSw4aMIT2cuJQyDocDtMZ3Ugxt9CzdYMviTH
y2jyke9t1Iie9LOU1Mml2WP/bRCxPez2uj1aRlKxiXkqCVOr1u4UrBR38GvnyNDKR7OExJ+BSnth
/yi+wyTie5dQfAlcP79+8PHYYVoVnOs//VWK8rILye+tYg+k+WwmjdYbX8P8g9HcF2HKrFtA05V1
88e0jHrENxnBOZ5j4JFUQjAjX0JkjBTZY6Wq+zvUW4kb8vpF3gI/DKEfzLRqS8bvhODmttsDswuM
gke9305NszZGEAf42Tgt4fiPXT5t0qChWzg1a0POFVmkmjTciI8vtKLQGkg5yJ93xNoI4R/+fcjJ
bIS6V6+BpxsjYT2GU40lx8cIpViNgJhIAwlPDcYKSVbzb/ZMLbyauxENunWkgqpPDtTYlrHE7QDo
xm7YYsz0taQSeb580bhWpznDxeCkZ7HkAVAqu4dtF2YvemwB5LHwUX/E6zCGZySUIn1+uZSCX38R
9YxwSTy7i0mc5nllJST0F9Wk2/6SgI2apv3dMTe3cu/poshcrouFWAB7II9auzIVL51CFHA5jCRE
ZZMT0DXUdyMQwVy0GAnzQebuwW+JW2KFsB5ti51sRBh6qMK1OFWPr8KvaoCZo5Q+gaMHNkEfXRj0
0fguEx0Inyl5jtK0x4F1wTvZdNYIqzpi6YyzorBiBxXVSjyHbKnkQOiFeeI8ICzU6WquEQq7hrJw
qKkSoL5IHtf3qTJKuef3MfqGD0lT/99Kvk4wPsXT0ItsMS0DatSu+wZ7ifkBOAXe5OSVFLgLw6VU
z0c45bh+E1Yx+3YJwoKPpvQRpA9G5/3PgH8ULM0P6IUySBwOfHMgUYcJoqqcEMLhwBT49jfysENK
EVQ8Z5KvJ2JjnRF3NicNyA5SHgeMyNjIBtpUcYXk6D5VEdORWg6pI5Y1A+k+MTXuT5Z2KkERxrmE
gXyY1LQRCXvyPNPaBIfXAlvkb/oU8sv8MtSxAQ6Y8TC9ay8voXhyYz2bOI4ejqCBWDedZcalxuAP
eXw1nVddBe/UGrCxvG0Ao2PWWOhfMk9svgHx99T22t+NSd/9+Ee1ImM+3V0G/UGyX+k0x2gWQ7o3
wAktWxiOus5TZo1YkL/IUiTCqgveeKdjw0wEPERSJoodR5BO3C1XUf0X2oe0tuJK6W9d0O8qISp9
CZbaERwpKepcg7jeMG7YulWy9mVrzsnv/Q32Q/OGPPisgQQiVcI+UpUi6Sa811BkODoDQBedhFHd
BtJydHHSBZbbVwqEJqrxTUCrXGIu/fdzjZ+R3fhx3vcGjZMiAW4Zb3pI34Gda0a/dmC8Zb+JlQC4
jUtIpJLI+TmhNvgRbbqOeodb43CDI4ja/CY2ldQy2giTajFL6YixCF0ChEIZwQq62LxhSdDdWBJI
R8mEAgShznybvLPTEbPaU4mu36/wCKosB9P0RaZZC8Vo/M/A9uBfDMeIidCGpNwByY2+i4VmAp12
yPIKXgXYRF4+joank0jSlJvFw4cxZr59vBAi+f4H4Zsfg5uURvDN5juZK1Yekqw/BKd2f329MmT0
NT79NM/l1XBk999VYX1KvSsRmUSwvrLkOmBt/h7VWSpPsrIwDgeRDTyKQEF3kKl2Ooy3kWd1qOWX
on7zUcppSy0wR2awbtS1vPPgMPc4A4v18VA1UCo8Q7JhajyEMiJ4lbTpUNhC+QW39H59ys9DrilP
3a9OQEEOr8Zd8bTO+mBVMncAgoxfeo+QCXcoxOXT8Ppmu3oCI4S6rJ+e5GSGnFbRgUdWDWbL5bqZ
ZYVJFp2AZeH/wuwsfPgwCLiPzMf8v88MxSqsKCudwRs/539DNyrA66YalCGuDATKcBPs1ynBzCwk
k0Gp09SOhzr7WnqrAHXHS1OwiKRm7J5rtFoO8zKyX2So+F99rJbTntDHPRUgsjtekG7GoQxKWMIh
dEGLt0zsylGmmw8tpSdvKICX2woMzZSrMUCM4JyNC8yXdktRu/SCuIvHqFC8IASANuV5qlJa8WdV
gSEtHgCxjMp9iIcMBjIte3CmmC8+pztHpYms/4wlpuUbF4fXERgBAqQCB9HojQ8FBewQjnsgMkCZ
29X6nSO42BKqMQMebxq50dSrMMvxBCCmW+XE6CTIoa6IkeT3HXC5dYXySGnIC3nex7K+1c55qYZ4
R3TjWHafpeeLcKRDktvkIK2Ltid1HPEGUGlzUkpyCXAXfNHBA/3nNPZ8vtlnjbJ5VMitT9BLLGe8
je3SVGaokUdyus4LLjtEoaPQ+6Z2gTBdKsLKolp2UTxiGehgilTgY92Q6plnulQw+6Cfi7Lf1ytC
VCW5rZR6DsOeqyCptJGRSXgTolIdMgNGIbif4MPHEvzYCCv4d493kXpX3sjH6ayS0iDiRNdxIl+x
ZjZb+7a//RA5o7RkmPg4bVGay6Gcg9to+0xNVl4in5kjVzXH7UvcD+YMfXi5eLMMqy3qyjei+WLx
6JJlZgUZq+UYsAZj8onV+uzWGnEjNtb4Hnjz4X0Q5z71Z0VUqrfb4OgU4PepQH6sHwc6yyc+F7Xl
mQUizcSuwbG3AON+Envkz8BYesFWXT/fofqVgptJVDxrDU49o64Zs7+Upx9S6UKB3ltIKDfHuYIU
zoyhyQBQ0vOhAin+F8DCo+QkvvlLmZ+oqkIdqMIJQqXLacaz6Hs6dLwNDCfeER2zF3ertC3TJHf+
4K/8EU9aHqqTybqCbFiR8qj4Zf9cYomtDt/nDAeczLgsAgyoRDZakhYLM60i+/6uYwBuTVGTgrWE
530L+KBDYkN2286oyS/AKsvFczxHDyxmumPSQ0Eniy48nNREMqqTIYU99FSq+H7LahePuSXNnScp
0IZNFJodrG++mAtFoqpW1CTxDa9fn5dQ7i3iQt88mRkSPR8A7vYXbYfKmz1dK3bGESGZsCuZRuAD
g9eQl/AkLc7ORxt4ClStS0MFyiWpBjk6oKLV9qh7ApOLzCND8UJnQ55tZjF/NfDSMhDuUORN+8VN
Zn1r+pD1datRxIVIX7Z8yquLHwsLzDHnIFFT7QI2nF3an7aGnPJopLUU3a1/H7zavnAGtPsRdOue
CqLGU9VZ6hMseTRR86V7zrhto6ixcVqCWutVcID3R3Xdflp/4ezDHBxZuiuc1++ts4vqJ+yhq4YT
ZNolF8PoRrGNApuOeQkgswnZAIhdFuuvxFmWRefI9AcWSuSwZeVN6rjgjBJm/rRIikW5GY2l7qpZ
806bPBeKX0lhZTIAVOoeFa5T/3yF0iqn3OifCloHZGTdW6KG7K9pHaA/FllkJ1i5dEBT62V9QU7O
1Mh2OkswZlqlQ4OGoARdgnJ43nLdggU9dJTNFZU0+/jniiKJInSNQFul/3pzApJrEk0g7ydI+VH6
aIlZUPjiCjSa2PAdR/avnp6h3hD3reFZB5YQNBMWiW7E4MKrwgEiZxmIk8S4kkeisJx8BEOgOWM4
jMVIf2P9Qgn2k6dQrwRb6+HkROJtGi5Rv/oJ/Yz9Wwp6flCu65a2dacXQAGoBCGUKFIgtFuuRaxr
jSVFytY45i2JGvv2blRvJo32moyR76njATAq2wv1zNLiJiuMjOxr4z0eBV5swrplM/RpzaHZ7cku
XT3jxA6BW8el4Yut700yYifavOsqhkmrI+NjpfjlzDvNQEgThLNT2jW/1chG1V+RBO8A30N/OZAk
seYC+F7ZMDrSscjTjxxLz+BF3UEZeYPT1akq+FiyUeuxCLvu+/uJOhaZ2hR6L2CaVga+avdjJ7CB
P089fzfFOeDHbKiwVR1+NZaUzXNXvnFNdjuG0AQQcW6bgatmFkXo558Y8RGJ19WbtwBcILCZe5wY
+WARV1EZflTN6LPC2VyGy+tDNlXDJJcpyNr6m217WemFV/qRohtYyRKACNO5KMU0U8i3GUX190lY
S7vfeD6+5MI53GEGsKEzpjagIXiMwP6fZEmHxzAqfTzdfJMzzRCaY6/rhf+o3rbwIP8Osa/3iqhy
iWld1Q2wBPaSOT0tAcK6QcA8oTycZBCKIKigWibZJtp4S6nnPJA08U/2DUdseZPQRPD7nvy263k7
MZ9k1a5kkViTYNhblwiKCtnSNOBUzKrRx9RXgKXUqI8HIPQZvzmK7MERMdBFIkiDabeGiNr0djm5
csglF6g4zpYubhtwFQpS37RA05wvD4Vku65fg8V8H/Mh/ZdhU6qelU4X5WrjufZetNKjfSokXyPz
LZHY03c2NwfIOIMNzbsCqPWMGZ8DuOKMqdmOwRiDQSmJ4ud51gaWT/mqgVyCRWpjWqnwsHlFXp7W
VFxuKB9z27UGZfqPdMu1FZ3byOw7AL966M1DCKMamPaLwoE2YQCNunTt3c3YnYbdIwsRfK6wS8c9
w9SQUulnl6kztugftu/lIEG0ccVKsv2Hwp6VxGt1ezTajNq7mWpQY24gxWgSG85rTX5i7CmzhmoP
20hPujIAFxLt6m6F6IuFJgOiTqdA4exltA2yWcvTXCImETAuG8Ej2TBfrq5XKWCe5KR4fzZI2l1i
YJBEsGi4WU3XbZrWs+5mavNoOmDqwDKmhPtf+xUGbfaTsMykibR28oFXWHKVtD6LMtcR4wCvCm2J
78pp03//IMOkvGec4rBHOKSPbE6bzRK1Z9dvMmMMBCaE/6ljtTYA5xnyUqL4tvmKE9CnhrKuGWF2
yf/Amg2g82Z5vkg60etxMgDfthGC+Xc+hLjz6Gn2+J9zpmZsYu2j8yajGKGA2PdlAOKcBJNg20DM
F998S0LvCGJOuhNYF+5E6YzsXAPomLabKnCkHExVoSbHfNp32dyga8mpb462MqFIz5FZbX5SuiPQ
mpqu0Y7Wn7PTIuhO0nrpqXZ4l2u3IGiBLsy3edC4jlXo4GFHCvnd+j8URyWeTTWadCVlM9kFSJjY
ZxKNS62rWp/yPpnIFcASNZB3XxoObzLy/dMPZ288weB5Hck6sJO5hFd4NZY0wW8fVynal/LWHpHT
IFYtEIwZsqNUXDANTI+TZ/W9YZbToJXVsg9adSQfNMp8/cFrAjVGQT83YK/IY4PusAkAfhXFlISP
IgARd76TuGWr6qMYRHEOlZMvaNfjcE5ik5xvH3ZEfB6btKB5dXjyFKsDPE8VnvYCF+4VPPHz3all
J3Urliz1FQzhdtxdw3Mv6AjMlJKe3mwHI118Cx8WBoAByNIWHdYhkOcQQiESP4fI0uOLE6zaGTgk
GMswfYpu+/ahe/eOk8a5xu6iNBsIZa462Xprph04OVel+FnMI/DIrws9TDvI41pbvYP87tc+41mE
rYtTMZI4dLen2IhNYWyGyGOUj1lPp9+Lj703ElVN38oVsqfuO3frFwIhmogaJaO741yz2Z+YCW9C
Iwqlk8hpyzJstvOK6zib2kFb+N+x9uDOnEcwG3mEFU0cP/4DLlTBsIpbs6LFq8HW3tvOQb/8VajA
RTkPBVFSn9xJ19p1qMWTJpda4TbYbxpg+pMJ5BBpwY+XVl+E/qkn2e40RPEDoGPbSEQMZX8zNuSY
gwsB1oVKWibakViwPiyNgcnXoRs8qOtCE0KZbNUXLDdPYyvY6v2LKLBL1e49yCtX08U3wO5kY4jc
l3dsCBps0HW1uPT1ueTmBxC/V6ZwEgu1VcEhAhC3dITrQmdYacIJVJJYvuSAmQ/DzrfdiIco42sa
8p/YmJw6ploVGLCWU4sw4GlEmNRSRqar0GZudVPSR67hE+XqlRuD42abRw8ITrvdj00Zr/XYmQJB
qaz2Da3M62XDBQeLtV0WZY5yLt/xK1mj3Ubs95KgNt3fjxn7Gj1eSIT/26Aajki2QrVRK/NpYZam
sMzFb2g8e56NPSR2fM5PAe1YdV+XH4DiLqKstWZEGKGLdy5FvAvMETbPTy+rLip/wmqinJenFwcN
qmOYM+18W5SlH7GIbSvXsdzYUbszWgbhjEkMPe+1b6p5pU2FGG5oItomOWn8T4/NR/rM7drlsgF7
DNlnB9xp18Md9xGl3k1AKDJ1+6PbinuDde9WrOFbpBg50o+MyFz13ZkGmpP+mY1GcIPkM9ifufTH
qLp+Sqj9m2x9l8loDFVsXQ37ReQ2l+xvV1gtM5bXu0OElw4WOr8kKnN2/PiAQJ16qHP3z222grSn
2FcKozmr1qVQF4iTJ8oJd6CJLOrOr8oHHZWDjFZQpcyOx6CxF9VC4NvrCGeoj14ZXxT8VtYFBpMK
5veD9g9aVDnkPKSMECgVF/mkbFc8PZ2fmedQfz/xxhtPCfSazW/eV1y5e6HDzm2IV9bm0d7GFX/f
n4aDgFSGSogCtJN4gTv8IeSDcRwW60pYKCCrskNOSDj7UnB/1jNOgmqDeSdT7iRTI2ycFHpM/ZiQ
QomV//gAxgJXDC18gsCQtkFbOVNjWWe0DNRL+4RI5M2fc6sAFZB202Ot5/MCemRZtykSfCtuaF0q
DV3yY9v0hyXzsSboctCEciQQP6azVhXdBthSkgtYG/9oazT8g2VfmFxQ+jYZSyquAnj6WBBYxMX/
Sq9uxdLzgT5K5IEoFCq2jlJba9bWYmFtF6/OrlQV7zORcH2sxizScdeAuwerexHuNZ+HZTumoA3f
oLERj8KcQrCZpQ5WrWMSxqdIB2GEkMeJAMg9SeecCw23bVRMJCghiE+6e56eHeFsQKSz4Hh/OT+o
u42gjsjQT2RPwCWBR+RLvi9brFfJOXege67USerZoga8vJuXhcFbsS3N4YQ5k13yo+wfB1A01Kzc
T1n8sUcjC/GasaIE/XpxLdyFhkaF4paVgRVi8n8/yFM8dxKSlMNwboVpwjnGe3l7aP7SOaQOdpkT
u0J921taXeuJ3wN0+IXdpV1NwVMTMiscNxzwI+yE3B8P49MjN7c2WHk6c5I0w2K8/aIxQGvEhynR
IP1jdk3uhkXRX3ISSyMPu2fCXLeVEVAZRBPJNKjiWGmtKiIndVl7xTs0AaGylhjH2wTh3N+YbJf0
gOQx0d6ZLecFBW3EiBh4Tkvy9TOyzuNJLZHhlJhJ2Jqg2+qwTd8iQeh6q5vt2ydbFUPjQsRQa0SU
jmGixrMi57zKcT9mye5E7fgR3fdOXPAENaAZKS5EnRUggugXQKue5Mp+KiNZL9Z3ZlilBDbCHAoz
pDy32QG+2+HrTR/1B2XyXBZqGJO55nmCvKiQqSKdmBSJo+87/obfu4k7WELeZ6oFwWOi99+lPnqV
vURX7EgSvEi4llLNei4YJK1nyTeFaqzZ3rsaInFJbZbtNEkMnCJOG389QaradjxYYj4ttRWiD/Qh
6ABywg82yCw3BqCNsNCK0Hgf4ccUt2KJIGJOi8j65KmySLjaL+rTajUES5HrBSSj0Nud3WQ0aGNV
YAFPLr35HG7ip/bmsSREERffIM5VfiexoBi2bBKF5jPmSOzRfTGRcBEHQoenk5HX6zWyz56e46PK
AaMe80Zox+lVEjBt4YeDUKLHZPcUf3M0yuvk1eoR5euMuqYYWyhXw+OFiMoK0YO7Yt0v55TJGFKT
G2rClGcKlsllFYw3PrLnBr8E63b7ooxsuV5O0RkRsyvHHZeTnwPjrZ35uENmKux1GoFwVfAUnPAB
BaYl0d9JOByhBEhO+XVd0mbBokaPotg1TLGgP8HhBO+yfmNO7fsSNTfGOjFc7oP9qopVklBkKH7C
YxYv+zC4Fxo5mx7ezpiDQ3wpAyAR/6f3XgnktcLeLovqngsGQXmd/VOcwYx6PCcEU/I1KgeAKR4J
5FPAHIT5BD9WukCj2Rdvd7uKDnfWF9cmSCM3Im0Zl4FjGPu72di83moNvRRIjevKVzMtHKnRd9zS
cpa0uB7wQL51c6hXBaQ8G+eNGwHEO+c4GP0IPCLmal5cwUezwXBAGQkNCCDlimndOtgRwj5G9auR
AB2nlA/+VOCB7LuwXE0XQWXQen32gG/MHvXjhStXOjpwjYgZMAHkMysVJHU8LH/IaVK4Ucm36k9L
4Y/KwiAJWsRmsI3qrP86T5GAj//m1aNgDyAnlhs3ZONboux6MHv0okSWINdznvsbZzqAVSd1Py5e
lvv0801ZfNgJyeJ+3dm3+KXrZFpl+KsGU5IPoLVtyzIoOtnQyfoC7dEkoGmCkxf+YOHHggrabiDO
UeFcSEm2WmcAR45ZOWVkM053s3OVSfIa/1+46oZevPo93dnlnd5FMby4w2ARNXymZYr42aOVWwDO
l/vk8oP+8h01wxi+WL5wX9w+Gnvzb/aDSrC6ssQ7rK/tNDJBvZm9AFg+WLQKvBUOnuJGtqNFBpPW
wIj42ngbZKBDPxc15gAB1HApkZHpRF+qhntSxaxDmW1q0jOghAp78v5fbOf3oKmyCg/DLDNnwRlr
jIDXBATFEz1HOBgp2tsorXeALyRSdG8RBYXfwaJRfCcEbveNFZzN5bRDOCix5KH41uQihLNsjH6O
K19+oi09diO1rsyg0UyHFbLXkRmdRNo9eDNfuPPODfA9kJj99j6DMQwBvsRx34l/HYNdZ13Krc1j
e6l8sRRiFoZ8g/VLubgHwgnhxbXBd6zhOzbukG8SdAP3PHMfV/FXRhAuUGHh97mjQsH5CeKSTF4z
Pr2n+J71pyjcDsAeA7Tyld8fHDFqtOK5OKOzhmfPYxibdq8dbRsUqJ72GjwgsQ3TMpQsCbrwofXI
TyaoLlycG2bqfccxkWnHD3HsptBc5ux5hj0x7gUQ7UIorNXtd87J+Dll2SCXjoN7GZMjFwaN4/rk
HX5mcrVwAWsWAGSgY+oBo94ttMQV2iO2OypXGNJSIf/7mgLoeYlS6AzwCA0VVSljI35eS0o62oYu
/uO3+CKr2NiHK5bIWjXt0GLxHhFzicU1+8r2xX+Jpru2N8RDl8P9p0+ZxZRXqF8Jwz7fHxoVuvAu
S9i/83ahZu8GCUNMa16OQRu4EZANV6KwoUnpXIpkGrFIcxJVJTyIMbMW/mVfXmfKYhkNV4QJVVKM
jfxzudgC98dqrJD6xYzgEwHEaAZb+utyb4m6avEoMk5eHwNfKA+pfl5kbUC4kuBfdy2pqrPguMvu
wAVY6x5+WiZWX9y6sDaIbksoACtAtn5+s/4qeYmcFVRU7azbbYBGIBER4ljEf6m7SvIbeL56BUhJ
zT2sZK/fi/HznxNVkQr2dedaCJgGD+KtOdy3v6uVE8zyCPaJWhlx0IByCfHRZAZkOzBMCfEyHTMg
A8piV6VZdEYtlTeIM4cw1P+7ITdvLOSBGy6VxM1P2iCHurvAtsnK3PMdI7LynieZR4FSWHnJ9prr
h4ylmDrHm12xH3fvx6SWLVAszePDbEsF7zXJniHvt81lBn9Vnt/iep9cvE8igfJBocsoL/quD1gw
DPjMw1LGDIDRMQ2JovvZUJm7qKR9v4GM6RFa3ehjbVnyvSBJnd3lIzvuMcKJtHyoQkmm+TLl81Jk
TK2re50kdtpMJcOxL88KgiUdIjiePDLqq7WUZVFMnGCHJOxPO8hp6e8NrgH91/pbzE0bflG6yHyk
EaECq+w+jkNRKf88vS4RmwkXFz9dbxVj2itfOC7lnKtP86Yj7GGFatJhcncWrelbNx9ZEXcABUGt
V9PHuaZyRkZB9Aob8Jv8LNYO1PmgTcHZgMcdEPDPet/ms7/KSpBykVFsia1Vu+LWmmCur1faC2I2
a1UsTFrnkbEeZCPQPmS2knph4pnl/0axfNf354eemGBy2e5fuK66++ag0AHA93NvYlXdWMab5JPt
Gqz+UAMnhYqz8Rh+oy4fGJH0CxS0wgck5gKOTeSA3aKwZAU7GMij02lczlJztOQ9ujWCQDb0esuI
jwDA3fxK9/dlJocuHQF6ZqRFXGtxvQZAJBGMYKPZyokMUNtmxT5EzrQyLCauqgs0A9bjmbN0VNp4
4ygyo5kYNZKE9m8+K6+02z3K3qXbDlVlsxGkQhJ3u+dNV7bj+YEk0M44Ip0cDGK8jf47k+2u55LK
kK7d6hpGO41CSd+10v0JmpfKQGkHMwa4XCT5xXxLOFxF0QfiOyWKIcGIu0HZP7tpds2bIU81WFS3
j1NRvseeMnAn/GMQBXhXN0b15oYkaZQRrMrwcQMpGSV4kXUC9bEftDbZzA3uVRPQlg+LiNctGxhI
3W6KhGUMj9rkUUZEMjBpy8guJLa0C6foEfPaafrcZmrP24CoEnya1VRpuJpCsYif1sLxv3Vfo0Gs
i5CvChURNi788MOZIgkj5q4+vol0b1/vtP3oJZoKDtsqVSDCBsseNNGq1yze5icw9+WkXUeIXPfn
Wgs4LJKTrvqms5thd/+9GDfnSkSFaZb5sIeIukYsMenyipeZo9aFo6ca4bN1VUAtRB7nlR+3SiQ3
3XJ8uTbZK2gEPpeqvt8FV4engehSb8hPWH5ACzYgbVSiGwzjaeaXTCbMOjbbd5Kz6G9u+5fTtesW
U+6FUMLYLGzDJR/pHbTRNiAR81eeGQe89vYddZ+2bLlFX0s08AJDUqkuebsy5/okvGHX2iNEc73M
18rxWHCafFHAwasHzCgsIPM0Y6A0BoeV8d9zIOSNbCAwoKHYAuKShJXIlpi/KdxpLNml+gg8M/v4
E+wPGMbndfbYcGDBvK+/evFUun729NgBbBXx70v248dCHdxfe3a5JR8lbAi7vja1ovuezTAlLjMH
w/KC7s++uSO2oxDTv3k5LbzDLkwJBipB6BQybfR6tXPWzyUn770pWFr30tQZ00ZjHciLk+kwqt7f
nD/9huJmeYvuzbwWikWYwwcFY1t9xTW6LbDfjANeTyRQLRvNMzamVI7eYooVvkW7vE5wXjUmleUD
WDkhUXt/nejrlcSaGeg19yPeyuhOcYxYJiGBIL5W/Phs7evZBivgTn1kQwZ4miJLkc0UV4kDFrJu
XgKZ22d2p4nemc5mUOWXZ6XwagYFqB3b+ky9GrRBTox8GDyYgzh5OsLttK60T8KMas8JoCjjKh18
/3WKh/WoyPIAMTTHxlJDZjlqxBGo/bomPL0IWJ92MeLAhL1pXpWSHjpIbq8VofgUr1k7Wxymldu2
kKDxTcjg6CdVrBJbIzIGyTa2oC6CECuCVXPOZrg9KhlTJ4I7E0zKxuY5ImMRhP9ENSvlR5z0YsTr
9iQEohtKeXJR3dlcOnDjf1+4xqh+1oqTQr0F+Ivq5zDnobIHV06QkGB9BjNEBKoNf3lVI/urbnXg
DvZ3G7kXuCXlfj9NIe4Kwe6B/iQ9LuBUDYAj+TF8BQUTjd5RloKagTfn07waka8esY16AWl44uvN
fqdcQs23fOTrRCf8wEH3K6uq+R2RYV6zpXQiGJpy9TU3RcNtlq+QanDU/jFZEcP9gdrPy2d3ZD6q
EFvTYXSZ+71jeEufYKLnGVUWIuYvVLpccQMySFGsD9uP9sqHMH6El06xDJ0cM1SOr5+WSoOVDkBd
BtQywJUqkrG+4M5kcX2Phw6bRaQp5Az+AJlPOB6iALFVzf0EaOpukgebKyMSPV85g7U+TuZ7Rhns
MQRB1VlBSnLMvq1rWozTkF7uw7QfZIA9q0sbkhWgvhTNWptPz0vM+fhiEXio8ADOlCTDPvINqL4q
GAs6YkA+h+Q/GI8eOAmOQ+bvLLx0DBHPzVSxusKjz55UYiJOny92PkVG+WIq2+DgLePZUbZLywbH
apxk4Yrb6xTySzt7K3mNYkol99FjK50SWh9vk+5xfxFfg0E1FYZeP8xyBrwJ14oc8iKJtvK8Bj/d
M0ocMCbnfMrlawUxm732Biwzbx4NH+UdhXCI06wPCBSgS0bSzhTci9FfxIG0Kw7FsncmT2UXG4/A
7qVUZhBQYQnEs4gYSlxkiasxp+hrxsK7pUlnCoLN9Ff9q9wt5pNMW7RyL7SKVtn9fUiXvmZVgsTc
p3cMN1vmuFDfy1CQ3SiFxjqq5cPD+ySbQ5M6wFrJjKDFDMT71fUDKYLhUDoMXBvsnhZ6AFXrMewY
duXTPnVBHLGVm065KwoTZkUkTlBC/YO6pW7HEEJJF4XfqUHK7YWCuajeeY+AVuUtsZvgvEnN9+6i
2bRVPgIwoCaGFJt3ezNNPtzpQ0Fi32DKjdZ11jhA0+Z3j+EYGaCoEBb1F4EjMIE8SC/kBckU2X6w
5rURcoaEl1eQG6fSfXAysyRpnoMVJJkVIhTIntxnBxl3FOeeZohIjtq1YuJemsqZkPoUi4/Lnu5E
xQE6CLugT/NqI15R8qyuyZU5bdNeNiiqDTLnbUH/M6A+y63lZbxJ7xeRa9+sCZEdGLokIZYU9p5q
6MLR0DM9cHygJ3DVdn9JddeCOH4PXjmexo9A/mrruf7GydC1Ql8x42Kd3P4zhMqrcAGnOBNjtGME
Cptsh/Y7MH2owon/XeMoeqB4vmsqnpTAcVqqkNeLydZ4vBmu5UELNjHKpzXnAhzU8YwShl/kCGUH
bDYGhE/ScDD3+kTcNBbALpbtQJ4euxtRFtkhd5yggVa1KkyQPBfGcEtqQcaFyUJ9zQ6VKRm1F549
dhpBGV+LGw9vzyynn2QmhINL80ymE5R/Fx6Ze6QiCGM20G4g3mqGeH89Vd/paX3LA/ZLfO5pctVv
1KT7lb9P3gG7Bd+vOmiMU3Jv+CcWyTh5Ap/mbcxnaEDWI+b9UyDV4Bg+SVIPdkB+cJimtfN3fnd5
wbo0Al6pX8bbUWeor8X14ZglvvFsgr85afuEQ38BkuibpXxPodF4E5zXwa56QCFDgDU0ixk1VaXG
Bd6evzll23JuHYH+kwgAvvHwKgxIjqP3Gd1CdUT0+h0Dhf73ypSzoelHVwAk90jWZJcdXtxkGhve
rqSObVZKs6M6Jf7fCMkg01pAtxIRyDxN8Ks2xVVa22COWcc651gyOn/ZB5aJCMkfDySijSLHp/GS
+W/SBSdsHhAxmJ6TE6sJ0SeJu9XjxR13p8wx4Lavgjt6Yg2pQtCRcjgONWf740SrvPpK2csL5ljT
tv4h25hzIzd7caIsMwcklGTIgPaJ9cYh+9b5OZMCP+dCsSs3EPB96iH7yDp36iK8/w4SFUDy+aPK
FSrrTQ2hdE0Xsa940xrHLIDifAXAwuLZdY2NffxjojMPd7Moks2ufQL+XANfpG2J5eXJkPbUT4zI
N8rCtcoP2cUAPj5KtiRk8EUpsp2hzIEimHD0FNX53Q/0Iwqim77k4e56HVZc/lMmf03GDLPfc2od
4bdl/WkHVELlnFwPGkXMoLTZPPlYSfjCBp5OpWsKvuKDgTF2eEv5R1sG0SgKzHaQOF7nhbAdc+wv
gRw0HiHuW7+XFGowC8jNqJxRkL/IfGLMhXs3GrOI3W/qstfffNvKKfNRd3AAb6Z2dM6NY+HN9Krx
i9j05ixT9E/pYGrtVseovF+0EDlcptCssZmrPxMHnAzVLfA5X/PDTS/aRRNx+QpnCqF5T3XSD3Rf
UhJfLriF3wK0W+MhEtjtGaUWTVjN7TdtsxRcREbg7GZ0Fd7hdMOSy8kGUvggNDWu6F/yu9HRjiUc
Xtli/1gAKYSmflyArErAY43r5PHH3i52Nkvfkh53yDx/V+ULsEp8j1EXv0Ochi5oY2rNJ0ZTGxVs
CGqJDZxoslk3v1NPnL+zLqmDL0GZV+gtLdlpjSBU/E5Cv4YIeIWSnKoPxEPcVDlKcAWwzDSIUmIf
sr73qY99KTbCXs9t8npQShR7G5nB/l4KxH1uNG+yc73XlC2KRPF3I1E/+sxhZmksoUjOTC9M7hx0
zvjt6jhlXUVMRdGbsl57y9LO2u3lsGdcFv1M80SR+rr/HO8IJpVTFTxoRt4U1TPAYzL9gYKhaHa6
z/PJMJr3u5Ts5gUzZyxJyt7M/CxH/hiLrAW6FdQOG3eeMUbexI8Dfu66aHU9HHv+4+93p/YVAvGb
8E5XtaYnGKdL5Suvo3OeF3Yb1X0eV66LqH6MmiVAJuACwLclRUnrrWO/eeWpbPVqW1JiZidQW23U
O5jarRW9UwJxLZRsRoJ5fgBdfXeaqDAJfhB25+esggZQJuNXG5gfmiUVs9MKeR1RhpgFrPGoeyny
mPU7d4sUVEX0t34JvpMS5k2IHTZEbbM1STsqHfFbluWu7iGCczYB9GqFViEu6Q7VOXTBaewX2ZKI
8l05+gBbMp3xVDJhAfODulucfDcEogVb1zVas+JfBT5ZJ0BbeMQNWqKHK5AgqcBx1vAqHEdvfhGD
YmtE7sV/iWUgqdY78D621Xh64oot0eDnwHgy3M3s+5P9HXwfv0KENfoPAyDU20myoIrRRDVOyss7
qBh0+QTsmP41PQLkBiq52qSt1gmVJUbH76YVdwKP/vB/ppQSN7zUyK8cTmZLi6t1BZ6H5fO+jjMq
lA5xwNddzX8WqTOvNzssUF+GwQNtJDoq51n4PCSBmOZh8C9pnUAaZP2i/aqc+HUFstm2YZYtPork
RQ1QGOGIO9Pt31mIjpVv+Pa6+qJQuECurZdnSan7EdCOxt9PNdWgncvt4kc/Kqt2Q1aN146C3606
Kyp6plZzDHoXuBWpDWP8CdaT7Z8avsQPDtk8YWWV7EUEqDw0gFqMb09MDIgiZvQ/oL1SaFHebgpP
ojTgQf7iv7OdUFSYIMFqUEJlnwLNhAZDUelP2C0Inj6lnTBPgtvcMsH3yeXoKVKLhxMUQEUFhsLl
Q9naxKh1xkzkmbsQf5EzHWJh0eD0dYk1j5SqxRIH71B85KohXhqeMjjwh0pumvOFk+KXoKrwQuSr
jVqKLxHXyHfSVKUmvAwSLl7IKnVrozP//FY++LPyYQOwgMt3nvggc8KZTZj3HURZCRzBN09hPCOH
tKsv1hDQ+uAKeu6+o6h+Il5hMYeTwZX9Mop6SVqAHQUeQoYI/35UO8HPGXV/5hdxhc8YurjzqcWt
h03Vt/BxBIteFoCWs8llzYki+P8eb2OpPdlgWDEGcZOOhx430E/rPAO+RZQaVEYroN8uSZbhb4FL
LZS/M33JSrZm3AJUcN17h8dkihNG40IXmHj7zTf8l2vyKVkgK17zzHGidk6b1dx1F8QC/drobVy2
9B17h1sLZxTpzsQnqqN1oxKQni1TseFVG2Y2NxXzZnsqAoIQ1LYo8guZvysG1+3wUwC10JmXCPFg
vkJzij8+cz4n7qozZpg/HleTLOKFPHoHDxeQ11P7mU8Rubmd9EEHTBY+dIznHehUeZtaeN+U61AZ
VFPKM7j8yktGAKrOe5p63fqWUDB0LfCSnrcveSBz9L6sPQFEIDs3kb0Uar8U95mdQCXy5FEIxu1H
As6iexzAq81tULa0XRip6MDvlQKlcRUvXXrkrlvFVG2FDieDqM+grUjt5VePGblNelt5SnSmnMms
oAIVNiQU7lKbnx1ThMXiTNZe6sp+7/aFkquenNhYXIWeQKYAja9ez7VMbpK/WtGzRVz2jRjrYNeF
6cyRIx/tq3d2sd3c5mm2TgYZU3Ozd+m17ijMVeVk0DS5/B4f+YgJJT5qvW71CLiNLuBstKJk994B
uf5JJ4/y4Oh0ygtIYp9xQ8VfKgXk+Tcc6569TAoulza6aMriaHvArooDWvqwR8w9piKshoytX5bt
FIaXMiftE9SOJe/okhCynRN+vIKJGLG/g1AFi0GsBfaaRJVj6kdlSpCpUG/VvEYHmcRmqVDw9ixh
0v/7SEyhsizrIzg/dAT1LustHDLMZG5aI1CMHloqsOAJlqrv0rnrwkp8mKSCGwwqqNVvPRcjjVAR
eAKPzAqfeBBuknuMKkbtYZ3UYQMT/yUHXDWR035T6JirZqv6ZLpxshW44hSL1PlTaVuV9j6thqmK
m73O0C/UqG5qKORB1+9/mqwUsfdsHLL/c3lmtXXXbDQ3OAbFms7HT8skCz3XAjn8ivTOk8YUS1CQ
MzQwjp8aWDbW6l0Shu+5AR3+9sNctFCJ3GMLrEzHYZOM04I4Sdw+9SDgPrc1kW8Q9JxQJ4HBushk
xIZ+yZQSPBNlJaINkKCqqleLzcbqlKzKsB3A4bkZId9V05IQVXuVCLC2O/reXibQs76wRH3jhAaZ
ZL2QkqqIUjfLhqqcvVXigo9xaVPfRqbtsG0svPspLYZDwPpAsoj7V1LTqhliyGmdmv5YmVJUsHzJ
BaMe4qd9A2AKU1VgZgaud8pZdDRK0ci7QuYsPrEoU9P6zNhM/kdwBjWgGodPjhuFwT2NAnvBBLDj
IDoAmsLKUOm1ouhjqIvzWDf7NX2xRlxSeKZDz7/yVcevi4VF4oHM2zKy6vvV80/3WDro+i+bJldH
2wxSg0fhIj0Yyv5lkJ0TCL+eyfnxnOxHccunFRRVd2as1aT4nhKjd3MIYuEUny10MndvV9ltFdny
2DfOgX7ODRR2OjH2YoSSJ+nEcVPkFc0ak22kzjevtcJIhCChMute41n7cGHMOFi877HA7Mg8Jgs9
kX4h8yGNv5Bk29ej2ZoBwEREiKgr62wgQoFmK2TF5I34bEkgsCldvJX0sg5RQ3Aikg5WWrsaR6Xw
XdYfmn2g5cSt93b0etWliMwNXN7RKJKmgrdqsK21pEPRSjBOydWSM3k71p/k/mEmqAYpWnZLqNxB
3sAzKKpMpraRur/rGTPS+vhs8uj3e7k1XDfm1/y9pZRymCqcrKgpVKDrfRnQ6ru2PJ26MlM8WA+L
r/6clyNdGsenMrsmCJ0BkInfHFImozJjfnjUe7gZjkhjNZNjjoeV+DrwKP9qaVxra7VC6rxXzWfC
CYi75G1WpY6b7NfrvWsLH9l7sTpuzx9ntbKnZmvzYf6I62VAWoMyOGP/693Jqz2sx/tHAhE/hdEq
8NapHG/eLZFZsj2J1gSDS6TH2mDHgmRMlFohXmqyHoFZMnT2ufWzXCBKbiNKqdBUzhHpoHXlDkuT
3OLYkNLeu6eztwKOtnUE6eqyrEb/5qhneXuGAROD/enflHaSX1iPjNFg2PZpyu+c+b+2I2ESXNpp
D7O3JW0TUgVax6mDrInWvhpJFnywyC19PsL91EGh5Xad2dETPbw6FANKcTK8cgksKd5kWivxsrCf
Jg3OCCjLkkkHHo6l+6/CrGU4ItY5+dBmoyLKn44q2Zmt701FTbrGvuqcMj4aJHLEChY6TH9UCP9m
CtrNNCXNd/0iWvWzXdQP+zGuUyohk0amEVQLdCvfY1ia+8EfE85TeW8VjlCkXx7yzN94xKnR1oeR
tWxcnlvlG5AiBiNB3BM4RAUwOo1EuGKqpqfGF5AtQClAvIzOVPRui3rbMdfgJJKS9wnILyYyn4af
ut5nWr79xrCebu9gpXQWOiz+mcX/EUVUWoesET/kMdNlc1Kioab44TILOu4GYv1i7iqzoEc/c6sf
BYduJbuUZ5miXR5LbOQ3LYqrJ/ygbTp22FZev8+65tyb9EJOk9sSssAjOFlBd7caDBtN5oC+nC4I
T8y9J2wDPXiLGChbAXXFL0vV8ArWW8DflGCJCNfZM/CFNFMwtWmY42uHHIUXAC/3Bnrrpp3mRWIo
3dC2ZDJxREYLwrRteXqoPL68CARkxWnAYNVmIXNzEmmWxsyEFhn2sHaGA3hac4jxst7Teu3MPxTK
M0iL9UQJKFKZ1rNH8Y+/t1MhFxyrZwpEvhCQKdfWkPHi5pRqJtdAJf8wQkNoWLr7GeDNz3vghXAr
+w1CR9X4G6BdvifW3y3LyxYvYXYY21blzsYtAgDqVpTBk6M4LmioYBKfJRA8J/pPMOyxPdEiNIuJ
Xm9pbv0s5LIJdIK/Op6S3ERIpmpGi7xDh9X4fDNCZW6ikPwslvlEHwnv0gUOvfc4wX1VdSDqRUxV
em12JQWHWXr/EevnoxrxiLHRYq8saiDI4LaFL3MUPVyMJBT6RVlMq9zgpJ35dIpGwdpbzZVJWXai
llvtXR9QWcWW6JsVfJiy5U8VAFxTwQcirzq1t4JjKmoOY26ElETCJqLGuhtZhd3NBaAYr5wPSk6U
hzxAEoAcxVBppH/++6FzRhwSIezQcuLdMv5F5yhQClvly7lY6HLVpyJMUA9zE8K0AwcqapWDBvVh
QopG3x+8d94HYJQgIkkDmpzfGGaD04ZY/sLaccfJPn2+OjvJ+sKFknCp/pLUaR3bt+lFMJVQsF09
E1VH0GvdlbN6dCdyMsRfY0fqUn3UaIxJWfkguwCCiu0aZX8gws5r1vxzx1E3EGkjpt2MbBdUOVXe
HpwGr25uIVlWWWOYDImlMaM17FJLarK6dWll1ZOKn6VvF6r3c7l+6YBwQ0PNcIx1tQ13nmoVvzMW
et1JwqEChQS40rCljHXQ3pRzH3jUE0ToSH3ZchC6/Gw45AGK8sZ3f1rRV4JCTr3P9scXaCcS0ePH
VNCoXIwyKHDEYXD/Siz68/YRAZZjS8cCTiWMEFbNRd0yRIIl/B5R5ZnAA542GL8rUolKY6+Se9Rq
HNNi8Zrb0x7QprCn7O1lgg7do6AkdpyNnf9rsbFx7unZiT7Ju7GtGOl+fc+RzBpacFFhTA1va5LE
bpGEnYNbiGYRgxVA7nxjWU7ssVA3HfNMH5OgAisxtIQk/FL1wJHhL674N3EdQ0r2D56zQxGbfpyP
bNitZ03nVl9/GdFNYKxDCTxKbh0eLKUJcWrSuC24iuxNNCKwLoARhyefClwGV+TomGfUxDgBtqoP
1q1L37+2sNF6s6xTrB9nPTuFgHkozGbp4gUeWgBnbKzhiJGIgj8OnIkN6JltcjxjpXhOnDZlDGav
aWrhCj3faujaD6nCf5VaQPDAExg2YYXUaN7B4HHIy49UDjLB0M4oHl/TwPWZ+DA9EdZQVhMWMZqb
ibTMl2w+CMlWoLKEdRr7sLY4YRzMrmOF+S9RQVVqNg7ZyQdgs3/GtI5o+zRruw71adweG1laacHF
ReVqXI+cX/g8xLHOqfJXlozGFggJqv+PyKMh485TKvJJ05fAJvmpciqp0K9oJwBE5LoOEKHJdVnM
fvMPgcFP0hZmRabnUQG37M7Oo8E7BQA0tlVRFnGrVtz+Ry8xmd3BmxJlY+ISl5eFhrU3GrnCeNC7
ZIGCNXql8EfYtLJrP6yqH9ZkMwrbCBrDT88J2Lly8H7uAFd+9jeKZP1w2LvRxu5MpeuAV5Cma7SY
FjOhMy7hK15epFP3moNhxJ2dJ/vccgjwn64BKXAfjfWc2a9GB9nSOgzYItTc6Hw74X7LxIF4wUvl
/qpei6RzYjLOC3wD8Z+ATxtw/EhDNIJ5PzQZ/B2IkKXPFR7vYu0Io5R/EzQPcbwH6X58dGbcbRkl
CTt42UgCxaIS19I/a9C5lLOWnK89kNdu8Y1hx7bgANfJ7utdnuK6bJPN5vEnS/Dox2q9Y4vKqMBV
Ah/ty4qvpJToNKzGGa+/Dn2iNbQ/gHMFbQA7v3kfs+MMhty47y3krjVQl/Sl6yBGENj+WusHUzgI
/4DcQhrx4ECUe6R3i0gHfpy5Qmyp1FebjyCdDSaTPY5/NgGcaGuoNSBQRcayGc/i9fGy+SqluxRP
uMBOD6/52C6o7fi6uAx5gtGg0f3AwKwNti+TC6KZjaoiWS1p+KoJIYC1CHhiknRqSxuRlzh03SA9
veL/D9EkuaqHmMiYNw1V3q84ba6gqFCFPhRPVO3y4PyL88S6tyg2fLNRV9iJaoLzC0GxCb36crxj
KP2XklWinBYyvnc0s5zs/SltRPNByUuTjjuJnU2Cl7Cc/dOc+1SKED6+jp23tINyEVExs+VSvl/b
x1VKf7ZThGun11iFXjrjQAAwxd6DebYf30zQVNP3T8h+ePBRW9kOrLIYxWV4lsmgTKqTSIUTFU8M
hBLRlCij71ZhhYT/C57cLqmbC8UcLt1waXWSkW3e3fIzHbcPmSe502N0llMDWZqRq0lgueBt7+gb
p48fUKPgrVssfkKPsGwfLdwcqNvbue1KoCO9622CVjoxli0kjnI97SP72AldUFl8mPiOf37W9YOu
nX1TPKF2bGNiGwgdb3QgtaZLIVRpQbyAkdWlExHWQJMxo+bPW0bdZOKLH4W9CY1crJNoD5EMiOil
3EsIjudZYoAXyAHHmvsk2Nnrb2PTU1LWCeL5SvNJluAXTEY4v0dgY4ytkhMRGURBEVoGcPlmKjNW
NQ27RXcAWeI0Ta/pUi0G2UEZdTc+hv6+NunJ0sCyhpmcFjiwGq9Fd9gl0gRf1YxGFj/saB2fK2aQ
jzFBnj5v5+Sl5OYrHhQnD82pdwZwz54FjmXWARB43D7wMtyGGSyCsqOjdbNUNFiXe+SAQNCrsrYr
ZJDoa0mQCcCpQ/pWA2LBpZXsYmZOI4JXljdCm+16d9Og6aUZC9hk1DS+KsLbmOhRoPZ6FkhvAqXV
3FEuCYfV+kPz59niHfvWDTSc1tKmPQt4Dc25Qs2F2q7s4+LaW34lOiuiTPpSzg1XM2FZ074/YoAc
br5jCs4NqbEP759jHejYHHU2r57cBiiIGjylhBd63esBciEwt4i5Eqp0FO+RMU2/PaQtCT3wArsm
5By9rnfIWPCNXDPay50amACHQ4yaINN2r3PZCkO4MrAzmcI9w4DSwJQ/0zivj9jB5X2Kf+KodGAZ
9YlWGuw+Mfb1VYRjOEFcvWqTjraUYBIAIp4e6l8aRAEECiBun5ATKuWQGbSqSMQ2Eeu8zDfcC7Le
hgy87MMJ9GsZhXSHh5ADZn0cmLvbRJbYAZhelysKbNOI2JLekZJT2Sah0qmH55YfHUjJAugHVKGr
1WcjLOXuiFaz9gy+EXUJuV+mAZVcNi+aUmCsFydCBl6oEESOeScEX/FxiETp2Nf8hE/M84JYobIF
L6MFP59MesWZ/hBkkv7mI+zcUv462maz+3imvxw8J5SjOB8tCHEYHFFhWCMEIvaDnW5Qfow40bTK
CO+fc3s9ReDonJ/4N9zLiYxEcykdysA/ZOClXg/LGSTFqdNA+x5uHK1BFkO0oXPgMwdfJ9AiWDxJ
oB/rHIvtuMEz4tIUR4Ongygxypi3ShlYFX5Es/RtSYdVh1xVF1NnVTAVoLZNscsPlK3zNSu2FBlw
06Bdo2moXNQnhxFq/i0DGgPrjqxzJe1ythnBsTOg5MizhOlRADZteGHAzgL9C1T38SrZeRU1jdFM
mhmTGhBg7FF27ewchg+xC/LbKXvmxTiDY1AWg2UAJlaA7j0yq9/zBNvz6lWAk+EizsKtVMMF+JUf
R2ZOIQ02W75NespERiiF532MJjzl4i0NNldkvKUjwiXFGPjbifHjoHtZ3IwTCzlFNt5GXCsYf4H3
CoYhsyaAWK3kSPJ9IRx+yfXNk8c72eEz7b3BSjLlbyYHBY7O6oR2uzui0GkyyEKjzRT+HPrgw+eW
KjRZfQHZsHKMXDKWaDapKAfaZrFApuU7gYe0qpxemMid993nYDYuHeqs7wFPkHsB+CFTaeKFtUkz
4l+W5eDcct+Kp8hyCiA3BQ+1ynuXn5A1woxRzOQn/DyYRpuXIL8szO4co2X37RuadWvvnc8I0E3U
sr6TD3iT7ub8PyS6ByS2SFWyJdc0jmiI6pPu2ygmERU+LT7u6R2nrpSaEn/CESKZcdvJ8iqVn2/N
hAqWUPe1w668PkxPFQs84DfcSDs+5Bw9yb20cgiCQqFnrFe6COxV5RoG08V4Le9LBjMNlHdfoNg9
vefrJS+dJD7h/aoMeMSzYz1oRQatC3bghMBvBVAQRUhfYZkIGjsCmG4alNaFLkCveMiENn1Df/8w
80QlY0q9EDNlIFP0FXjG2vYNtfq9qhRgFK6D8jLWBJQ2kL7EGSJVnrX6RPOOHZPNShy/s2TI69Zw
cv+mIP5lMcYpnqwb3pWHtJIgWKcm3dZID24Zp66xsgJhEntcRgF0hfGwkIXqeHi3BUuhdC2DuIJ7
+QNv0Y+OcCotkTfj9z33G1kipYBHed0WaTEXziZEwCI0jytkSQX7RoEGgX2ad6ZtOXv3YY0esUFc
9uAhk9ihYI1DVGgwHTeVqBIzqW9mPrrnHtvyWm7H+UTFQir5EeY5y17J90vNtCt9CRZmRmPvEhIK
0i2I1R2h/KD2wOOyrwtZnhk6MZImicdmXB8dWtn0C8LlHH8+S4ugAlLA0JQlzAE5CH1SRfWb6whI
wpqTJxY4iD1BRIn5MzRhLorPrZCEU35jSRAq/ipBcPUVtpf+DN952MScI3NXIPk6eUvYB+EVEpLO
dI54mngduwDYtrBpSUCkJAMVQ1NsOJCYhKcX6gdVUcS03nRrrrq5J8jocFGGatTp5myskhuEuk6o
4ezaWmgajgmhmY1cfOSfsOIWLq1n0//Oolf48WWRo1NRWhjDlBXciszrTwrl1Y7FrthEntZ2LM74
PC877FdH6FYx1gNWTj4lWmJEqFEBS5r48DLk/6ZMklchmPxVSscZLyzrUM90Pct2kF0RX22MSiuP
agZEGjQbCl2XiP3k/6nQ+JPPAYdWjxi5BwTFQGwX8utvcxwoSvrq7kSQNkz4ccTOQZRbyVpGRSXc
eurMl3MYZHRBZlJ234rpyysn6QhUYdaoXA/om8KRTC7U2Bdwrmpc0It5Ou3DvbkxQGaTzzFU514h
GkG7P7EAPWagUvxRY1NSH4e6lvZuAi6cJ+TS43MUOsSRV6OTwUElmWyfS0Rric3cW4YzYhEx3X3h
rWecBofVoY3W8jAr4QfO4oU5nXUYbGdz6l+PVnUdaLeuBmYSvPnqVoIr0cnturWyl2BmrnZ2ml34
Wnmn8ZjVDQe8UhLADdasbal+2ySZCrOE9cXB6N7gUBjnwkRR0Xx1iMcmxmqTDa+5X1BqrZRW/ALV
4IczM9iVuCEkcQSD32jtqiGfuHmu9k/p0NcyFLddU8YtHjD/Y8akOPQpLxU2MjeMZluAz6WbWPcJ
R3uxiCpriGCvyZAUo0EZtA+XoQsRROe0yiO4bi/QBoGghv+Il4M9nWCOu6ZRhO7sVbqmlyx5/ZBC
gXWlniCbnUq1rKTWg1LCunNgzEyBF+dA63VdLQszB9OOnUK4ox8aEmPe2WgRaV0aG8wleGha/vtT
Nk3hj2smL3XyCg05UzY4AJmft1v769Cdu84bxVIxD1ONhRMDODj9zkGL4+aL4wOIphQoFHw5a7QS
11PdBRMsq1XjQ7IxDyK1IGaBGRbhkF4K0A1nPJA1GyEQnzQhiTTTaGnj75oruylolRwy56AwqRD6
XH2QoG6ejLywzihr2v7msMADS3bmi7hSyWOEEXyZ0xvD3+E/t773dv2eu48zRq39kd3B5YpfLyF+
reeJ/NYBRYVv57KgXHdvrhz205U5dD0xmjRwfr9QFEUTnfplMoXP8/CFT2PFXoxTY2to3ZZr0K5X
HxySZ0oogM0g+d3tp6/NK7hdkKqbe2ipru4I+usJd4JwiDhn7wyrBHTZBKGlFhTWoKG28eYemJfT
Dr9H1/+KC6ksRQp+C46RwwDDkeNM5fVwfAY9zIsImMAJMooWm2ngbe85hPpe03e7pk3v5oVK+m0W
LuM08tuTgeLDfaj1R0UI8cA3iz8IMNBif1vSFygrdgMimsUX+Kp6oORJFz4JL2cauNJKXy3b01Rj
s+NrssWt4b6nTUZCXeM070M2NSW0RDb/CiDH+1rNWwADtSs0Fiz3YAJmQlFgvLdzud7w5dulTOqd
LWvWtFmZIgGkRMhVSUna0+NAd84mxfdHKvkvUz2usEnfQASd58AiVVPVRCngnv+6zcAKUYlb2xXP
7kHDpqdgf7foFZzUBO50QRN+DosVzx4uKHfPRc/+s4SmikNOB+Cfb6jH3+E+NRDtWPDocFcSJkwK
x42LXnp10xsdVD1kx8m7893T31ug9MA8RAm8e/W4PK23o511VPGgRVrWuGY0+sCPn7b1jD2kKJKi
wJ0NoFEWqHHIUcrGvGejoNAI8qnLjsHcy+1NbE6S+rSCBlVLQJZyWToonLIEkfSmFxcqhWHYE4gR
2eqJcoLIgIrrXch80/1VKj37lbjcjmzeKLltVoaolYEfGtAB8ce+snn0xtzu3G8gLzmgv5i4K55Z
B4qBuzCwxryMpjvpIfnD6Y6q6b4S7dI59ICOVYGds/7xUTyrIr5cxuFYRjJcrxBSXH65D21RHKjh
cL1mHH1tLAtQ1X7Ra548hAjjq/q0E9zIKwHP5U7Ok/68dLUjPTnJt9L36gdUOnrKbHCqWQ2sU7Ln
qtOKdrVa80yY1jdzspNp3whxPO6tm6S94OTn2xOaJ6UxvBLub/0CTv0vz+jrENzVKnhxm5TStFsd
bV5+Emo4PkTmh3jo0tvoxo4smHIvdGRKuUkPcq3vCrYPt5B6ptBQ9i5Bvf9KE0JcsUDTUtVCcfR+
pmEL98gN/Cml9ewbowwGMTIFJLGU7aBx/KL+o+97a3zspNXMbufUvTkHInz0XVhzZCiqpMgJU6aR
xnVrn81VOSV8ZEoURcosj1TO2VUr/FX085pMiNpXH8PEmJLyrPeXK7I/29xYBcRCYqmPlaEQzMpi
0VyksOMs6MH3Hv9aJATfM6zbhzFW5G+teQCdjSbCTu/e23nowUGTgnBwT4aTrhD/rilk/08SKtPt
05M46OV96SHrF31a6t3C8u/7NNf9cGgfv27PznNk+f15ynJScxpPIt85hHzPlJKFjIqEx9/giTnF
rzcNCrOyw5mcb7f6wYHkC+0I6PnShyprfS59CTcOXV8EOJTQMxHzaf5vpwGUz2bvlrl0oHaqo2T/
neL+bjVhKEablGRALiUkXs8w3RuqEUqm3iG3C6m9/11cmdcfM2SHRAfoxWutkvhHKsiWYjp8L6nB
lb51BWagaC1SdZOorGMvSNc+4gtX7PHQ+9j02iiJX02TIsYpooQQuAAbq8JULKPxid/n2dOuwrlh
jfv4j95BO6ZSxe5ciqn7/uU6Ir/ADetXbRkrQXzg7O45TTuWaTdQNsYOJ2iCNPDfdR7MITTNLr4T
nkrYlaQyDncRKwpwUWJmjqjIAcWwi7DSI39oUCQ1rLSb+IR4ieWzD2drpUEZhxBa+B7rNegVLm2K
esm7WfbdQXZY5EEh8jKHQTBq5iTNv6gPGJT6CP6cEGTddM1TvALiKTa34Lr+K6wb2n73/OFUUfe9
TpRBySxSG0qmWv27nyHBes4Z+k2FosW2oXGrRTzTtSgpIC4KnkTi1QntlOCkM6sWvKiVaJoe7RqU
RZXHnjVjOabQffNPfiQTTrscbY35IPCFbDsj7bvsqrFZNz7w8qyg4SjgjkPySNpYsNUC57RJhiW0
7rQE97Kb7CZXsxt1bpXeOGyFRtO4Gn4c4Y9i4tgT5Dwwot8NzJKQQcsi7ZrppCHy8h7QpfGmjpKH
OukJDlzYw9RHI1ttuixx20HpuG+50QXzNbb2y7u1CnJ+rzJP75ftIsXKAc/Ld260JJu8OCobQ0ON
TwfNQQGO96XCfxDFsDOz1IsCVzi6pVXfPCY5lTG5vk6o36Qr8itOd/ZAfD/qF6IEUOcu/z9W1wxz
5wjh0LrsVwIpYXacDBWdi0edcn5A7H9FkJN4+4/erg8duWyWnRTha37DH4Wa14kFuznDtoYEaFMd
gbayEP+iOGDsxj3N5qrnyQwDHTBXa7B9r+jZgvo0Aj13tF+ikIOph2672QWIOHvoF0WNN8nDDaDr
S2Zf7ku5cTH/xXfLwabRG5ted+8M0z8dRINj9UvpGPN5zuuQ0VrTqxSaq1J995kMADsnfRVDtgMj
zEN8NDz8jLAyZxJgj8jVlqr8cyF5zOKI+mPuWSK8IXgkcTlC9hwMKoUbx0IRoOwzlkK0UlCIIzsm
kvpym/wjPF30X39A/PCN079H/iUOGW7P9+a4/a1jr0+NXN80vCEzSONzTYJQs1voTbdT4BUTB9TN
76qePa4H4QDo5Fvfx2OG0pvA4WiMd4q/20+iUWGY81K8O0fWHFLa7NU0HwG4ebjubzWGOAIeIfk6
u1TzVNNCojXTOchsNk6T7zYKjUEZN6U1XVScAWw62bgeV9v2cFysEvfK0tYOnve4Q3dxIcjMW9Gf
bW5UIiAItBBBVwrkyeV2WeekoVudExqtu7MAi3+WEJ73H4p+OrTC4IJ6r/I7/gSUFfTfqZHj6Zyf
sEt1tFANf/LPMB031aoWDjkiyLMu6WHaVRy+4FbYmd9NRcYjYtbvtKWjVv52XAL3lI7J21X+o/wu
VwyttNUg0LWVT8uhAYrKpYLOoYbJoX3Uokp4QyYB60HIMI8GpoF7vHLBAn3HmQXxLTJtwuQqvc2t
B4aEPpekCfzWP+PASQfxXDC/Ais4rkdOXwqKod+ZNu0l82NfsTGxPkoavw+sbt+b/m/7mAT+es1V
ojcwVU1ctWn5lAXi5JnRMq3pE27fX1m81gheV0AhkOHiMRU23rFj2XPjUCI/SAa/cDL+jLAuvBpx
97p9PDCMyQU5KIxIaGWZXA5VeUOUR7fvW9+pUE7KHrQUTTCXSwOuPYwbvEv0DKGDr/HORmhqzxwt
qUm9NFYS/6F9R2XPjHmbOSj8jgaX59ly+nTsSjrRL8rL5176w/Gju+u9lxbM/vljl6SFunVmJIip
xJpSVD7ECCtFp0RZ6utaNe0r8+nszPdHABxSJKA6sPEaehfoR+pyqW4iCjNRs6IpQRePZP96Nc2Q
2Nx+JQ7AXuRDnFngediNe9bRD8x19zwLRs6zwjhL/1dMthMHq4+m71+FmcTit34eILEmsXtFdLrL
dZF1pM7AokbQL9EYSwuzwpfwl/9QjqfQiaR+IUF94NvJZCz0fimfaDGKISpSBPpxSXHQPfoDjgtQ
h4En9bzRRjWHIw2otkDRXSyOwm1cbqsfCpAYvdCxlJVrG0VASfsG0mJOeNwvt3aSwyVBorJTnwVg
RANLGNc6NA7bi4b2QmC4vKKcvcafOD+99Po0b7N4AMG53D83qUNOxjMatiQfJx3MvzdP97RG8cy7
enaJT8S6djLUzPrkAkkfcRTnFZHjsDUkEJmLO6muq7wyAkAWWFIZkvWXBhAoD56Y1uaa3KUrl54U
a5xIMyAzdXrRm3CgFLWD41VUiQd24Yu/hFX0fbXyWv5F/aFhxd9zqUdHJ4uXVDM/QzLaNBiZXNVA
MF81iRyK0lbXCns6fEEcR2JjBa7+t9aqcXbr3DY2I/6ohl26kSbsg3MvM2K6KaJbUZvLSwneBJ0d
aAgiBOy19roeAKD6C3skacmq3oBvcgUeBmYmo0lJIAlkP2/5eTykJYU+qkEIT4jdQ++d5Q0q6MXW
IP5fMAfimdGTyETJQVu3Awbn/AW2Qtj9BnWWEBVyTtXafakgPD55Ilf7zUprVg1jQdLzQstl1+1Y
sBhNZOUSJ94kss1EoMaTyq8Ol45wPdvPIbozmkqonm1/cgoscUriq3DD+nA7cLHJO8AfIUxjC92K
pJKr/59QdRe9KtIlSKjqkzCpaMNm93lf7vTTWWLyqABvN5JKLHFiJt1SvZ5/xebAspq9See5+vfo
Mb8bGAtUsUvPrvQM7W/64ylHE3Al5d4chMrBjd+K6Z1a37WXfcDNpBfywVTq6GHreMGSe7bnHXlA
J9KmjN7yE9exCKQGD4cG80QZLLYIvZdNE3G1cMPamUoNdVlAa7JC7TAfGMVrq5re72jPhEDV0m0F
2Vl9VWtSHctZ4kq/URx8SzDr2ICw06YyAbmfdti7z1s/IoU7RHiSV5NJ6K1WNYx0RH8wBXv0dT/b
5ww6nojR1rj5dUgx66Cqna305pJyOlZujfOvqhqtt6zoAT7vwmECQS1cp4lX+MPel1b03/aUyvAK
fFDN+YlD2vK85WMq0w4S+fOFX473h26LKM3ScuqPsWKstc2RqxqnU10rcCMaE92D/nUpd11RU0XO
gq6aQI9VyFQfPsFEBRpenFiBF5VJl+X8Loto3z8hE8R0Q11J2J5r63BTl6xw3msIbYAmSns1pRZW
Nraez/5rrqJTb68H6xkPX7akX7noOpjJ5eCQDILwUXDByQ+Jhq66BfULNEU8wuGMWauORph11X9p
3NQWS9os2Wz96LYdwmgM483im1ikHPinjvsb7bwdj8x8yXQt2aL10mOAPSygEPxKFXkyS/NQ4ojr
BjTPrupGNEsqVC8BwF6HX1/l6T1ZXPGkwaPlkyg4cNdPruLJwkve0q76pVkE/b2TWJ6JrtWfN6Z1
715TqtS+fh4V95zuuNVvOaGV7OPVyQTw+3DpOS6SNE6UZ+CH2v110tHu/xcZIp6CQpuVR4Uu8Vy9
n9WBo5aoAOf1I6ecOCQzJIZRWH0ohaWbh8K+OvbtrOAVZPFPCybI4IhqN4bYdujA4Qly94W++vLn
m8g11MsKgYoKF/W+9DSkt9Qrtv4FGW4TApaWKaWcQfTJ425GpRuBZ5v4iZhN7HlETLtxSOoBu4C0
bC5kztZKK0JUTzHlZ2r9R/v0b9ZgNJoRDmTqcMWrGXgH1WjJFSeIBjtTy/4SXEmd/r5gBIsO5NIf
/zyX8C9hm+GFpckgQG3sXEdzLFcHoY4cUN+VS/1SpUuGRTke3/Lgi1DXn7TutMvAtpPxWxi30qJf
cQ1qmOw+jdypSSMbrJSpE4j5YZH0fjnpoLdGmh0y2+OBV1RdvMtW5kkLwXRnlQQn/lLoMeI3o3z5
eN3FyZVoFyFsUz+0/xIlyZo5gue6GKI1bZ+Z6kF8xJ9EUm8cWhYr+0/aTX8rU8vruHI4uYbh0y6m
brk+QXs30+o1eCbWKc8DPe3Jvcm+Md6zHKXy/Wa7dHe+nlSahDTkT3BL5twjWeldSwUbi3L0Vi8a
RPaRFEI0FwHM/JdsSJO5Rd96qV8P8/wBU6uQVfct0LIDjJg9EqOj/WXRjFultvY0hipiFisa848L
W2bNnsIKzY+uUMJg2aVTzSfXOoWnZS5RvRZadwjsh5Hqa/UppN8TUhNMtB1P4/mrhtlubtgbFs4k
P8YW+9ep0T1r3nyprmbBQpo7Upo2dsv+YqRYVEr85cRth1KIIOiai5F58XFVujN25+IeOkFLNsoe
V3Km9vL0SHlE1jZyvIn950xZMmBzbKc3tumDXJcW/17ILG9JX47547VBOYPN/hUS/3+ftuwawHFN
zOzrzkAurSEy51AjPWePqJfwnNpw9VzmPVFJU3HIz85xPNTgaHYGnvrYMTwcpaq7VN8uQuqjbOu4
It/44Wr/dLneh7Bk2nSNJeE8cn2hEuYpbypNl8sAZTqEfcIpU7C1xNX1CY3oooHZLXlSnDFvMDZv
lAvlsf2TrHJzIXYfvbsFLHQJpzU0+w5AJ+mfZdOWjk3MaoX7OuCl/4M2NMor0I9PczSVQ6bg2b7K
qQE9YFtQf92U5NHgoe4Rldm/Pe9WaNUzgrQ5cGaAtPZF8kx03DvOwgizOh8wCM9uIAbBZdSUmIeu
zezQx5fGHwsAj/wAnW/AMAamO4+1bnwYoO7I97/+sK5nVJW5Akk8dAuuTcv6EOmdYZUrgUReqMZF
NpuN4deGQ7+2Q+Q90+jbyAEEQ8gmQgFfDQk7u9MU5/PEn7IrQqCIEcx7xlJ+u4KXPtUmQj83CH5G
2gf7M+eliJm4SLIpekWwWsX5e+aeWHj1xMEEngrzSX4dUAXOoJklg68omEzwFFB6/aXnqd2B/Xv0
V4IR21wf50Djprfl04M/l7wmqcSn8v6IfADbZcGz6Vyy0D390pRS2jXTeup36JeYCXmqLKU+7NJw
UgQZmuDgP/opai+9kBFbaUugzsgJOG6V0cvN/mkMfQQVOMA8l/TsFqz+AZaUS0saAf+GweTZ7H9u
mHryNThIjIa3ay9UbjOQmi+VoY1bRN8E4c9/Ub318S5jME3ZvP9tE45c6vxW22I4hHA8MuuItq9c
8nuVDCbk1IIglTDyHq3u6Hn9k9ofoQaVZ4We147YWfS4Hr97RLrVLB8QRYSfp4A0sugQ5vsQDeWk
UD3c/9Sdm6/wbjPiuLUt3KJ7RquVuZdX5uMsCbit5sbiacJR1xtbw7XLE3sUhezGOY8zoesgosUS
/xwtpyki66kGF1fm49RDZ98e1uyEywl7PdCv5HEmDrAvVouiqxx+Qy5xjYc800sTqRiDU7ZUYH30
jPZudUiMt4WcTlJRI8gTGRbm8GGDZb+4eRYJn/hmgc8ua0xm4EUSVVNiJYBHs9vKBD8RMhoOgvSK
s/r4fem/LjHrTa/a4hcXnweEelQ7ii79l08/Dl1GH3uebguRnJYuxTni7gUaB+9buqvm9W8gKV2V
zhXBKkoZOhDZc2w7qt78yYhkKTZn+irrBPdlUczAgQ1s8SkmJVMmMWnMwAuRW1FIwhvWlJoYXHTK
krBUeJwJ1mErSV1G919BWlPEPam//Oz4sLthrVqdtHvr2FCv2GbdzK1j/Io4AAOPCLupMUkkUn2r
Tp1a67MO7uzabRji89F0nxi9Zf21KgEE+/SaS9ZIwnsqptEwJK2qlRlUhimtc9zDxJwKYLg7fLn/
zykZseMWpxRK9A5m+3yfO38k8pqpBcmViN2kKUNgXhDRH/l3DiA6T1GecpLG4HetEzUyDpQPLC2W
lTS7Ne2DE1sc84pHGM8Pp4JG0x0qB4Iw4TQNXvu8AmgiqNrw4/rLqWao3WqzTWzoiC3rmgil05wB
D38Pl3C4FsBRwDiY597xRE9v/uY/kXnJngwIyIoEIa6L7oPrgcZKrnOk/VO1cnCaj3ncJ7yaefFH
NZ9lrF80Nr8Wbosed5rBkfDCkWNO8bG1legd5cJbtZDyPWaJT2TRyR3gKymrYcnTZAVJLxg3hTYc
Yt+vz0SRJnHu5EVNM+65vbZDIkUS67e7njS9iLMxurYVh+8XAmQpKZdCJaYjzt3/Bl99bwqo8I9h
MOJLs3gJGfmqdpCJpE49PzPUzdn8owgo1K/TmlHM1nSZgu5GLQ044a222b1i60HPXMexZChcM5l+
nH3I3llZX4yglomfS7RLmghFli7poAfgM/UYINtRJc18iN//6VAcVqf9eCdXt5rVFgJj8Eq6BnNe
U0B5WgaT0CV6jrAYJTCrawg87ZWludVM9O2qGOZPSypCkxxgYssLf3T1orM/mf5lVMAe+ga1ABt3
GV1I8xiE105RV5kquFsoTA2mWPfH1pb76gxe/1rtYMRMnGgxCMg2o8cYxzuYcKIWs5P1sEeuAt/R
keSq/2OOLLS9glR0Or2Mb1Q5SGYHQ/9lPLsbjlmfNSYrzZHvAj8llvC/Z10xOv1ZGANiH3KS3vwO
+bZuvU6ZfnjeJLuVZyh5vh3tjpdoaPSK9pedeEO+JD1KiJEVdfCxTPSPjhHSaWfKgUbKcTxfkfxI
M2+QjsXeaXT/aX5gP7gAVGhCns+sCze0RG6YcrUj/R5n+/U40gDOlc90rtb5RD3saShFxBumANBn
Mi7VOV6qo2nzbk2DD06kD0fM9ehGcGPcdQ5cCHXOetLehO8mcF4d/UN6NtihqZc1Pyzaf5BPMp8U
+5QInp+RM3ien6Gf/IqPqsL9PzsayayiAyKj1/qeho2FP8vvluaUX2+kVP2G3S9RKDBtVhq3Xh7f
g2hINdHprh5/PmMM+yyletQ/zX7yVmmGLqhRVruraO1V7rLR7Thc8gpYd9doiGnZ5o00gVnArr8T
naAyDc2KCzNLgB1VOPAV7c9m95D3gcRLWADeGKovsmmfkavjw22kTURtkqhT9jc30JXeykOKba10
RkxMWKiG0DjzVlkEEAczPrTrcEr0AEyqutqL2aBfEfg5J0iEaHaBpaFcGuyj9p2LSmHVCfrBz7io
NjDaffKLngV+Z8AfCAC4noMIzLZJ3GHWro95LgCM9/qx4bsQ1r/djbQEqBikBwVg1Gt4qM87WlKL
cV39pMnmAwsDBauK9E6n8lps34gBI1COItEpjrKpPz2as2FTCR1QGZyuEG3yBGRHg7D69mpPPJbX
QB9prSJdJ1kLSOD9hmFk5r5WGQ3Lv7esIMiSsAmvo/vDvUGE5pmSKuFwS2kkoNW7rs0IyMKXatIg
8xRklMWMOfcKY1tBymA4BZtMOA6qoCGnBjaxW4DldGBl/wSg4/y/oXeaJltbQ7iCV89bsftqEL5s
sz+XftlLbqLpd5vNqMZ/KQIfSp7hjst95vQ0+fOmZoCVqiyfjYZg+bGuJUM2nQ7EASkWCR0T9iJ0
OipD1xx9GFbSS3lfzlB++qFZBERHBd840YYZgL442PnKg3iMgp+ocwyUwrFPkwh78HgHvCWx9LqI
3mpijjeSzgSDY5mU0C3LLkKGRI6ha/sJvgUjkJwCHub1wfxT8JDFmwbgquXN2fc1ywWLFr/tnQCf
dtC94WGRgX4TGw7wLwvsV2+tCIItDbMq4UfNkDA3RbgwMutyj3u7ew+vubXiOdeq69HrY49Fo4A9
7T3M9nM/vztNbx46fRXa+uc6xEhxblDJteMejyZr/RuJwhGmu3Ozu+s8Rt3JC7Yulv3htdblYJkv
yyRXLXGtvcK9Hy5cC1ySQ8EvQLwaCmyleDWkqno7C156J2yWAXifiY9vr+Alnx5vmg+pu2EMOapU
oZci6E29DozpLavTKRJ+0s2rEFEfE2vN43x+8GPvFoQbNImCeQWJes/BmG3BQR45yixZ1EUkIqjs
2ndmunJ49X7DseV38uAQYIf3NZk2TzQ83gPiqKVfldVeAIFcA930G4dmLmP5DenHzxvqWpnVzz0M
twNgNWgiQQ+2yT5lUcqEmHa/uLvgzvrIhg1Apx0SGy8hWfT+NiL2Nj6DzkR5EVLK9KFRhb5Mr2Xa
Wfrx8iBPFRDHvs51BwKDHm6xr1HKWC15yEp1oLUPOAL6ONuICgV2D4bH1iW2JTPYFpfpAVQmUigO
RbgbMhCMqWARbn7JZHfpMvBGufYxUnHz1YCn2Cik6eqSGcvozPt5GiLIoWnSbpClTvzjZehio7ov
icjNeGApxBV0feG9eLdhpSy/c6DDMlUmzns6iFZGkP4a+X4yr+sy9tesAZc+Ghw21uexD1icNDFM
w05z6RXR67kHOtudBaEQX6i/Dwy6DPZXE4DPgGJeKvEH10XI1FiPwHr94XYrhULU5VCZiQXvpCjE
Ytv/pByoZKjwFfOwjf0LEKUBFGe4oC49aQRnnuSB0zyRJR/mCgyRRkuHsTsy4EMDXHYHAJF5fWyE
+4se6LSPYlObjHZNI8WNUI4N3+lCZQwnvmRuyrPGizNkBTBH6pcYjwmFHosqyyiNul/VE04hdiO1
jXDnRfalKjvUfzNLc3MCTG1cOE5NPM5RaIIwH0MmyMxuljcdHEFWVYHN5widlwPbFknxVEjljqsn
9nEEs5cHjAIsoo7YnVvlvwZ/6Kwpngt24ZfSDNiuc/2N2j9hDyHpwAU2MOqUMWUzDhnw9UnL45pJ
ACK+X+s0GjTrQzhb3hZU838gfjtiiZv/Mo9W9eKVgkZhPP3DyAMaVDzLo1qYN9w4SLMY0Hoa/VMT
+73gUdGWC2S6WD6jNSwdhEbZvLZIMwbyHDbQ+TqphtLgxBh7dmtejAV+1Xg67PgA5vcDOGRdgywz
7kRXDNJvC1UIj9le7wBm7gMJGCO1N0nXSyRSbZ+dbq2Vst8i2qayTnMS9Z7hni0qMaNjJu5Pe/4U
tRRzHdRN4+zqyXdsI6xUvd18aaNZiz1HWo6yxCWlaX2F9ioFWxqKZZYX0eqzU1tMrSe+ZWTRRWKd
Hm8TY2ri8hPOajZpLYAPbnQlmQO+2ekAb7GekLPTH7kLuQPpHM4XvCTnjr9/pTU7Xy/pjqaFxcDu
Q2QH7a3L/mAsh30sXmxdB5JTaqQJKaZJbygJNF+UbOaxQgxXpBw4rJEc0KH2CvZIBsDKR2XmI9bN
L5tKN1aQ+GXVSJ7Mh9yNINYM8EeVKOtRqwIAQoWRmuld8i/luH8mU8CnUDeYi50Sy8Y9FcRz3sGf
pomO0HyjcPhFr3YfAQ/BeucR5r/kBGfzPby30gkrXBl1lsEWYcHC8mpQv7E27iDQJ7CpDD8DssQ+
po+t4oU3YgLtUmHVH3r59FJPJ5/0FUfmGs/uzjWXbKBRP9V5KVN2N8iwheYNiZVpe3xLUoAxFEbg
tQeKpZYw8uzgVEKnY6DW6vy3Z8WfVG3VP7rOFWckbpyC3UEU9BIGOoMJhsv7M2hNg0pzmJ7TGQTW
jVjQkCgikRg14ZxEBRZmmj1GP8237Jf9z6NwiwyxhPVLBC1kntw3QDCccnIlrStq6W5b3CeSNPJA
XStOuydECPxXt01wvZIgm4ZZT6/jX0We3VETQybjsP2oDL82joktVk7H2MCNFL1JnszCCEGenSCI
2cdqfKtk8z9bpTaGDx79sOHaxaVyxR4pqN51AYf4Mqov/p1gyXywN0oFvFtmKFINnUwDhOBGXoeB
mNriZW0RBXYslqHjELp6I7an0dzqpDgs2MC8qVNndsn3F/q7mvCU9B2O2eBcbuhyOm+1tpZx//C3
Bo9R5YRFrVA/g7WChvUCk0KlIrVJ1uIDMTJl+duwJ/T49lQCKDaC47zPaRrIvw3jS16xWzeBxIkE
q9CNZJUCLlzyq+zGEZHoJB/7dAghb1oH77wzGu0HX88nmCdhW60pMHiTVzKYS4rr892Yf3pgk1TG
7hbJEnCDq+DLJLrfi1fp/E5yBF6gMCppulYRczK0v2bglUAvcMAzWkqN/uSgYatkikB/K9eCa81U
L8bADka584jwXIz4uA1r9y+ImcV/aPxItabuD0ykK3sCL0WQAWrMPwLRCgDq/D17NQU6UdEsvRO5
TNRhuG46tCAWwCvhKUA8f573Khsy9Fy6iOkVaM8+wdUHHSMP4mTlZ0yaYmi0bp7MAPcw1MfV1X2L
Ioy+yhOr+l5O5jD5ERtfS5CsEkpB1l7xxLHKvUsBiEX4vNWOQOSAepEppkBwgBwkNXCEDkHWoDMk
CdX9JOensY5iE2LBYisBqvDsqdr6WnAaV8kNW/DxwfWO8O5o245Fmpz6suQTJ/EYwQ9m4Iy5onMf
0c+Up7fyFVgQxd+PVwrj+uFzSO99SN4uo0s5EEwiaAyFPYlk+P4YlzLXd4bn2BQBn28s6nhJ8Arp
A/Sznb+yLTNOGoiZZkYWED9BuXiVy5RRu74H6CSwVo3ZHo2B0Xt7anenD4wlzpkdU8t/puxt5LGu
IbaFTVlcchFo6eKXhdUEcHRq69rzNkzSOS/BWSwxgZtczJEQVYzA7ZTPeN1GIyL+08s0BNKViZLW
AnEqbCu6bFfesa3wBGptgjRUeDnC3ilXSQAvpCcK40/UAeyAWiEngoQFbpEJi1fjLa0r0BFhI7Xl
MvLI7+siZ9Tv9pIQM4mVItBDXubWMkudS858Oud4Q/2UA/phDc/v7HVeFGBLQhjMwGm7IgFPR5zb
nosWW9QzNFbUMBVZZXKBNy9YSmO87mO93PadjDN9dWY35rlshP4m75LXWzHskaYDcFcqI2I24zl/
7VfVM38Xw9btbUqofWYlxrUsjZVRgTMjfSsSKjPhAyrid9xgNnmFHQhPfTR25NnXaAwo6kqkd0pM
tj25GVA+9Cng1M2wPTzZljW3XpjbCNVCRX37dxk1Hhz674HKRowYLZfLiE2jVMIklC574yF+bZV9
/xSANG2kAdetr9mdoWMvgGBP/zz7UsoHzMRLLltlMnFoYyHKrolNhOBkLKci82X/Dpm0Ibn8Wbhw
n9KUde+K8iAH5jZs8lz28seSuxpHd5zazrjXhv7ldXKmpDYRrmRul3rQGgXFJ4PRtKMPcJS3IT+Q
NcEMOBBEvPpPiPStgHYBVRb/xY9REsZOEtmx5RlW5vOM+GrYQJF4n7RWELVnEkzZ+jNsGBVaFZIR
9NVhums7naPWaRHp8stCAM577N5BOfzqhIJFjOCreaSwE/qGPyOf2AHqjr5oLxnHKEsDatQXNIUJ
rNtT1ZrP+ljxf7hXd7grX2McOMrgTDJhyTxvARi04KMANOxx5WpPLwfSmyKPLnkB9bnYOnufziRM
M6rBxdkffAdLD5FVh52h71vSEFydec+vHmUl4MpY9Y9IvSYksyY1aXAZtWLdRt2bEkblzruZxOhz
3LojHC1hweq2M1gZmolF1B22H+9902S4MWE3pefT0vU01VtZte4SftkkaJQF2UR+FeYGQW3jWjbE
Vb0IDoFZtV6dh349gfzHKVrGadySn/EznRV1CAPHwiUBy4NtFUQQStKQY9y+g1rQKefb2BwOz10T
hOknuW3kAFmV41q0mTyLeBQjW/R/Oa99Bn1hn7OXPHkpaxWv3Ke0MdPviivVlOs8PsXffKdRkCSa
f+iPbwSNMg0ouLquwA1dU/UGoIMVyVl83qbma1o++Jacs24f8E7csW4vrr17Pil9s1+EApmy3LLF
vbNjzNsXbJRHx9deIHiR0FqDIlmBaKAYoZl8Sn65u/grqflMBsJEx8+igSFoCAAuqEF4RTOcK+5A
Jujpd0uL6omoIx0ZHD9/zXOL6fBjgQGrdyXPmmbQvQFUxR1iBFJJeLkHUR5/H5JHCfDPu2dTy+uK
isI9nSaQi58kSDLERTW2hHaDJTo5tbOi8TgE0nMpr3+g4RuO47D0hgpjjmJUR1/0AGyejE4p8gSm
QCn9qNpLHQOMj4vTvNy55SFYE2dMsHWzTuOZb/qiooOTTyZbx5cCxXoYR1hof6iHMaqy0S/uVxxA
XzUr565rTUnYkhuRiH+TeJC/haA3NagCsrfHaIE+lGftIO4hDnbIwRLtFDmPU0gFr/EyXp7DDgcX
7Qun3K5NAf7YRnEDkJNf+mArlHiM6qoNqt6RUJ/EF2zYLrSul2WZACwd5RBcysbd5SMw8xyizsSM
D0XnnAAxz/cak0fW2dbOr2sHJ7V5Wgx4YlRO/Had/OrcK2TNn8v1B4p//KwQJz/WopElBpopePD/
TwW9TYxf+Pbkm7lluRszk1txyu4yCciD0HWZdBJI8FG9t4+ISaEr+9JaO05tVRoxr978TEMmHrVR
FFh3mUcwY8KeermYeUrs0G6hoKIZeFhqr2yTQIm7tVOAfulRTb8NatnlZ+CXn2ClEKXkjwtEbtiP
l8Vxn7uAhmJdoQQVjGfOQVA+6UOTIbqWhVGwD3EwYJt5r2EZ7Gb33ZQK1jQFz5JK9arm8lR+rseR
8nlnNpUoRjmJ0hgTaME4sCq8sD6H+rVhniM0Gr/HuqrBozptITOia9gesOupNCoJL2yulZwDG4fu
Y4/EhFHDd4dpB7gs6E3Io6GeQH2K6q07052w/y3gcTpKBapR3X8x9/hyMe5jPN1XV/pgLaUQ9DFy
cqJdyaG2ERvP7ZQPQBNSIymUjSSsiNSTg9PBqJaCpS3Yli/4l6K/IscZComVT9ZcvzvTOx0KFoHK
XwBTxytKzrM1Rpnn545gTVLjyYAJTRFsAeBy2O88TuwMnic98Vhb10wKvYcuUGFe2xhJI0IA91pN
M2Kdzh8fA7Vp362JSuNxcoXyaCbdphoWJH6p4IgL3x0tMs/aPrG/AMT86KnOUam9uVVBnXIHFKR0
VyXfGHmNYxLPos47wgEw2INeysbGwz/NRQspHJureGyJATP3/1xPPXMnQZLKoMf5J/3G+9d+xuNo
DhMEIQrQH8yeiSBMt6tTIoybcBQ7VsQ5yg1ZidfsSHCxXAbqDChImdb/Mf5xaSwT7MTVNOgzcWgC
JyFFwb3/v21nEmGcvq+KNUPMPAkcKfkFzf1yuWphDuPEHvJFYYbCuX0g8rdIjhr9jSuSpErUBTcs
1O8NbCIiuOoyFczs4jMSOzDHvEg1hpZxEmMbWwHFN1DjJWQsRl/vDYgdHOCV9VzR0VEevtqn91CG
KZ78fWFQfR7n3aAxeULe4GJz3MIV42QdVkIG3NSXtW9ulcw1wv/M+ApBLvI4WLbpKp4z5nefAVbO
umkPgiOxU3eyiGEafTbBgJIaigi+mQYQs35FLWCe+XdU/E8GOxUsbLg1nAppSrGXpwaJJOJje90f
ralrXab88wbhL+VBQXCjeI0L1094UFz/mUNK7doE3rA1X6BVnVHM1C9NTPZq/JPFvjKyXuTL8HHb
wbPHZGc+m2MbN7VoiC4JA8Belv+m4fceV0HvRr/Othz2a6cpZCwlTOSWGihBcKdQywiBpqM0nVI8
f2yfdKhlfNnBGJnMbWk2SOqIgAv+ErvGJqnSBWF60yi0WQ5nOYcRk/qIkih4W8/dA0DrqpAvpvlZ
dkwkz6vrv+9puVj6zPXXceEm7FfkOTFW6X6tOhnv/jWb1qgDlVu2A9624xyNWtlSGj9qBl1eLFsw
dr2prc74AFIlfp4iSdCFHghD6Ha4Q1l7sg1L9f0q4x3o5im/gKFtccEZ5lQRgHbxq86swwQLbOz9
E1c4prv7ta3U0uPxuCgWxsTN8DElefNBQF07V3cFYwdheGICLJovRAXMK8brWjOt2fxVsq3Uvj0c
9IzwcDzzNTdKQq9gfRo632J2ggFakRDhQM1Muiz7XEbOGURgaH4cEPJ7ZAGo9fd7151V8HIozdZb
hny6/vmCbAHleMYrRS4pTKHClcJn5uE86KJ06THMfVjLTg5kQSz/vQRq4SAvr5cGGcM+s/R77dym
bMzu3yL2tLpwMgx0+C4R19a07kwXJy4zWc0teZzFTw1REbZKZN/WQsghs8pFjfWj1BAf9l3383yG
7z0Zm3YqMt8zEI5S3/G6QX+a+jpQ79iO1sc72A4yeQGwUPwnTlFxHtRzk2UWmQruVZK1GpXpQjdH
MCxv0Y7OU/DEDQDqZ9busKA17LO+3n4qD9rtGMBSnV8198OAX5d248OE876nyPH98NGHg5k8qHrW
Oiw3O6LzkGMcV0lzSKJiC74KImC95ALvPeinzyl/iL77/WoBDjU74Z2wdvJmChq+qjIvJBaAT8sO
EB7wbMXnCLnnoR28VPVTLyklcFTIFVei/00JSppzjKIy4kMsY44kkirJBpUASAWKdhZIssQa6Fen
Ip7/bIqVXYwfp4SLcu+Lon0uu2YP36bIoBz135qtsLkzEEnIBqA9VaXf4QgcfQDOy3Uj1owsUrtl
M+6+TBXjRz8fcFzkJcT3KwcDLAD90ip0u+we6n0W9L3GaAqA63JQJF5sy8mNAbbnuIXt2UgKgpos
hm0PgsqWrX3gwfex2IkVvE8AUVZ9EpEVXTqJYRAqbR4RqcHE28tuQLmAY7znV6OydPEkt22NoIhQ
TEHjE6Ah60IJZ8WcvGrUE4Ourwr1aNGqvjys9RnWU71iOtbI3BlL91L/4Zf2P8FbaKrRIZx8Iq+5
4p3PPStsy+kJR+Vdiiwk9q1Y3n8zL8DBxURiYNiTeBqfB9bK2Phfut/1/naGqKCW4ZjjwOjfxN3V
Hu0usJ57LwZfvcSn9Ls3PIY9C7r+HqHPXaX+/GgsKOyS0nhtnydQlr7qW4IQESEtFvWTwFZVP9bt
7ffXT3ul/aMe93m8olIUd51PFKdGChaDV0Y07NCP+yNLyvnEnyUPpvSTJLyomRW7vDKKSnWX8DA1
xWbu09tZv7qDOMPKi365E7d0fl/WC/NwSnV6Tas4TOK2KXNkqYbNtPeya1jdA2mCkosHyTrMjHvZ
gWsJaftq9GBH5q6/7kPlwIDzmj4RKOgxu4c9ULov4h9gcjhYKA9RFCBffK/sHtn9o/W/1lv1Zuc+
YTGwymlp56clVNg73C7NGQDFDHp2I6Ykj3LuefP/jHnKLbOnmWmwYkxauqVF93PnzZMmrqvpP79C
/Tn6S11jwbL3tcFZQ0AY+nFNSfeMn95w1wP4c4U0pmU465B/boEemdigI0eQCqrIReYf+N7Q5BgK
0BT4RkZ1vVTGx6jRIvYh58EVvOtCbkm+oyMOgCIGJ7heyZ1c3s0gs5aWkgWS4SySdF6TkI4BadZr
uPEFNHlInsyJEshFiD/Dj2RLi48RwNtyEPZdZelTnh6/+p4+G4hkRybJeqIGHyXmH0OnJY7ZdcRW
A4W/81q03LmjPVyiGm5VZLUcxwK3qQGl21XAzxrb3x+IrJGOorCYFWmtxFELE8seN+rotfSxyFwP
U7BKf3BIh2/eLrg+2ZCPkFckfXmYIGp0iv8ks6yqIunDdmGBgrCfX+KgBcmQhygQVF0vik/cDhp9
2TaZLHaoIZfOdG3/kEoMDId4RdSE0J9v9R4E7m955DipUGXjCla+68aSKfx7ui/GHCAjFr7+CIDt
YOVvNsVqI0N0HCAal+dSZLI+K23idehWS+q9P+viz+Og3xdWXZKWlHCSjrMTw3oSFRE77zKhKCR0
xaa29WdsRRsC/u7KPq1Ig7xgTe2gAyXMaPQA4CZcWCJQZ1Fw6JrTcJ32yyqG/Ef3xSVMmUdAp1KB
4rF2ODjOTbOmvzQfJIc2/o8UPVUXBn0Wj84xL1kQqDvi05L1DCyiUdXE3q7G8Fx+7Rj3TJPtkTSg
e829GYOY8dE6nuq8br/Nife0mNyqU0VddAdyMGMEw6BySOjh5f9TNvayfkPWsFirEUtIHVfocvXi
oEg1XlE4ojnKAGEVtbICEBJefIKSsC3o+ZEyQ0oJamPwVB8uGQjrUpdEjcsCJUG5ZgwXOf+KraV+
+rpwviRr7a7GbX4zzOx2RpuNP2I0pr3TC0ABoi1+BUeQxoyNf33Z0bRNM5UaBaqe6HL8IP+poV1I
qG4zC4EpOm59XGl7hi3VtimFdJkB9GsR/dn/0TKX6X4om/AF97aNAQ6zFUpRnidzimeaHvEWpK+P
fJNOS3vWiI5gVSAIeEyTUvMwQBn8EIhkP4zUJ6bt3tal594EfE5IsIOZoxYIEvNY10zCpE7n5aQ/
bzcWB0OJTwlKFvF4AVhFEYQjxnUd+UV+fplg6tiDGmsSk2SbKFOdzS8AyGMIfQ1NoYMfOKgUqvZR
GPL+F1sIGqM7OFWrD/BEivx3zoTWyzW4uPn+IoZVLks42d0Lf8UCSP2F95zc4OdoWi9tgrGhHzdy
wMrT4SjEW+ZmX1DXlQ8W5jrx1S7a8ecTzTmtNYXghVjB1Y7cua62OovsDSJXiJsVmdlT09HM1yQX
SutllvAwTOhcnxsfmN+s4tkcocTsEgkqLW41Ni1efpXwrgYFpWL4+f5l3LExuu1G3sQa656dr04l
aJbmNzYSSneAwfIEJm6CdgomRN/yq1+oJDLdeXnCtk9ZqC8YmQYFwaJxrdjXdKA3ChFdpMeHiusZ
s87wxCWd952fwaH159CJbklxLu+zkozTFRm5eLzSGijTTQB0+f5wmp4LDuZILyj1PtGEhGPVHi4l
S3CvNcCosghsMG9Ha0vDINsDswGyFBII3bV/sArf1M2KaS01QP9ypukcHs/9NDiju12TGjhQ7Jt3
7yyIzZJM7VUThD2KgRi8BUVNUHRMjcd8CLomFwFDFRr+Q8kKzRV8iTVjVnlKJw3rverPfHa9jeB5
Uauvvl6QPf3hOTnqPngGPy9mvp4G41RhgDDLRZ///oFT3QU3TaMziHgSrUOlzynIFWROhAV2Omyh
PTV8+DFQ0k09VtkUCGVlJa1CQrzr6J1vQcq13GjYSKKmNsEd03ub5d6r8L28ck+VN1u4kZZs+KU+
TmTq3z4FqUHdAAYn1FcqX93YQEwmNBU4EMnG6whsaqGemzNLbtaZ7yKPL0nJeABwoTaH18Quh2qA
CZfncOxZxjIbfG1tV6gXiUKUU6oaADXHs1HibjoP2vZPNR8B4OCNdTYgZfTCMjot/oTOejuVxzBy
qJC68JY8RuCDlbMITvU7/v4Bz0KsN4L6WPWu4wIracN4OttOkoca/4hWkdiA4RsufaA0/jLYNQva
w/F0v59Seuq3pSP3+He2cvl4V1U3d1xHH6+O94IEEcH/vjtuUhMuDfxZMPsi+t5WiaffY9W066fz
+DKtq/ZGiBhx8JIE/dyRzjhUQ8BuX385h1i9DYFpx1+MlRJTRI7Ik5X+hOgrbiA0iM+6mmhHl/P3
t/hYhs/yYlPQR6slptvUwv6LN/s0QfDzOLkBqTOUZIeAupFTZfGGt8scgU9sqRLWo2KjAg9zkgvq
dwDrzAo0YX07u6+jetjPkcLmeZ13PSxCJq8hKgF2963cucPQ5LCigRb+hrEShjtzvXO5QHvf5fX4
bV/gUciDChens8GMAUfMOAoe/lnZGVnE0Ir9gI8wrEgtY++amoN+Xt9d26gKWqAx3lGQicX6+zHn
yBCGoH6IxvfDhUbABhGR8da1tgDRFs5GGNhjnLBxCT/ePlYy3I8fp22BLtD7YAUgK3XSho56AROo
cmauFVdhpofMyhHbyD+fblM7wV9bcTvORHWKTfuF+I+X/F0imQ6hUSfbHZdb2/QfpFaEQzYb5g7N
JrSf9cRP5IlmfjlCR8XjASv2UvYH1ojg659cOAkKygEt2GcWRWtuN3VA2WahNLRQqzDMHBUftBRn
21Mjgg3ufFugg4ijCNfXqS5QHf2AybJ5WTY23oCnOi/IxUqx6KfMiONQYpMsg4S39Bv5kv1LBTZt
Y1hu1keuiOvEqJWxvzaB7MJRIUsVSQdY6NcE52lFA//OpL2QkgJ9TfAtCzOe7w3okIgyGv7+linc
rKXkFIaoCKaLHPg/F0Prxc0dHtDyYF/m3YhKwNyLSQ3rXoYeuQaoC6hDJnUeFBqbiVj0kECOOAQ3
A1Iik8ED+6OBbCdixKKqrm7keICoVB9oN+o5muQJ6wrTErU9JzcEWcoTB3v/7pO6vMLjmix20h4z
cPy25dP+K+ghwg+VvrCQQ8lFsQBaxBEUDHDw4twFl57hUVP22AT/u50sSeJu8LUaLEU2nO2WNCt4
4BFUjemCHWj6rEhEIyleaPDHovMW+qZCvEdEbRZasvlqDh4J49r5fk6FSnNjGBTVh/6vCs4P1fJ+
jEnXVajstcDYmKFfVFLPzwiKd8z9p9WLXd+luilqwT6PVlQ7NIsz6rmzfWpNXrCfXHkMz9jU+jAl
bBl2E2H6fMpAz/M7JeYLB8gD2UvHK2jKMtaIDpWO7Awha8lVgmVc3vP9vSHUcY9B3Q9EQ6ZOlQIt
fmc9ydkydzPb/nIWLqn+B6VhtWQP8HpeuAVCZXG+I0PhG8zk5eM0u6KgECTkCSUpyQTWZlIU8lz4
hHf2QN48KqVvx0smSsTvP1+PMkFjmJKHrDpjB7Z0OWL3KbpYTaAOBe8DR882N3q7Po6E9oLREE6o
vZX7sTpJe2J4/8XoH++Y+mjLqk/TkTWR8iygS2WSCN37gj9LNggt8zifJ5rQtinCB+HheBAQLyDk
EQlvh3CGaFUKFP1zESCzFNK8WI58Mb7d2RY7r/6ATUSu1mVOQvgU1SDrWmgzshesEGHaX0Ew7s4N
yJBGilBtmznZqQTLafTc3Ck1xOEoNwST2mSJMzQsL3LzBeHWIdGkA1K5PMY8QSkoQsg4u8YxGqok
yXSTUYKdp/hnzh7yeqCGtR7Er4cGZSJDn7smSWkr/EcYQDoFnw6vE7RhaF5KfIY6c3CYRUZGcjjX
ClfdSgCtGyQgf7cF0ed5R76h+7rf9zkLilACIYv9L0ns7yB+KzeZAmtpErL5awC1/N9XpKP9nZFP
mNQJqemk6HrB8vL+6p8mCLp9D72yaixeHt6W8ITe63DWoUFg5OT98anG66WFsc5m6YVWxghIQwO+
V9bg7XMc/Wnz86Ygv1cj3BudsARiVbAQNXT5D4q21Hfaaer4/RW0f4G6Z1eRxrsb1OAg6Js9CBu7
QwNu+5pMx9NVXY3atRpvgUpRcirhCMw/Oa1zARKLxQNW82BLHEtiGOd3fcCQ/GvAhWZKrzfhYEHe
WfzObQmLm5LthjXzI2gHlWok7jVt9djBd1OL9Rv52SKemfK7YOqcJxiLGeJ9grZfg20HRs8VOC3a
fY+whFDIU9BIU6l0GGnuCrvNCC8B7U7jFa7B17C+v/6/AXgxvgew1BBTSY7Vn6hy/lxZXGlhks/N
vG6xLA5WZP7j2La909JXOXH9syDxO/T1Js8ypf0XY/fG+3J9FKiv/OWRhdkYnZZHPhUm8Z0/UGr3
8b9ygv4z7hIohX/5CacACSOmi/2XsLgneboky4dLCQyv8oBzaIkn0zroSN3LSpKaN6N1PEu2iuFn
ucEpgjdgKYWRJd/2ioLrCVAO2w0ZR1e+jde06v3lN6yaZbIJj27s5EFwSR8SudFwuaKHEouhS/AD
PtNawO8vvd2Byz5CS0ySIqy+Y1MtiKQSlPzv34SccMFxtkwFTzggu9FY5lVkOhEhNKPx7j8cT0AX
MJeI2Kj4uV6gVM7UMCw+VIIW7YEEjtNn50CgIEt6IA/O+ztKP+hQSjSbyrd5rB2+kjc0mnfttUGo
pfS/0t7X+CsM6+zw5zJbgaZ6amwtFcibppWjGBj9iYHoL1TsQMpLTKPC6zlCYWoQGeaM7r0O0Iuu
O95puAZqkHekShG78w4xX8/n8N6UJZ0TtxpSr0yZDmfwj4H+q5FM+X386Wk4cOpm1bdXijByc7if
d004z6Xn2Wd0m3KaRepU1EZK6Oj8KctUA3m5cNc5rtKeDnI+bV5O4OwlP8SEmxPJbwM7BBpSMRdB
5oHpxxc7yw0QAY/qN0lQoMfoqyNnuj8ZSNuMRQVGdsUi1z6o1+NjimSlhyE/FJU01UWNF8Eka0ix
N0ege9XHfCwfED8O/z5WwrdvRcySkD+imxL6gconN9PzudFAFaEsI056WOpofNk6NQT4jWng6LCG
y1lP61Tn9KxFipl+ahdhxLKUmsrgQNvzhdZhVnZifkLR+F4O2J8/qkISLLO1dc1d/QngxgFy8ZH2
fQyBscKoQcksXZC9igC5w6AHnl9eEdgPoqILyFuDXMlpA0FEAPrTwm6Gz6Ru6bTy6/B2WYaiJPjQ
9cbUOwlCYdTyP+xUwHHIUd8ubBPtKTPPcKbaGDyi5uoTzotWwVDxlhKdl5XfgrYyaSun/OcUwDuD
a4Y7RMyD5z3aXbMg7oE+N3fzY65CovEXhF30Y/wq/O+eDo/Mpkdm2TvkMIl812NpMAYtz+2kw7LG
yHRMZydOQU1k3Y3w15EFT8HkfosXnUbuw/b17uxHubF/25LPzbQY4wM3b4YW8Frq3UuV/l3/M405
WV9EsTpzFwlrE77Dtn5B8t4Pb75IwdecYgRMvD6NKYGAzaoO+K6pK9vMnPtoAfCn1nBJwz6E3n0A
Fwx0w4enKRko1yATaBvaOV3LGi9P+R3C/k5gsLn3sRygMMJRwH411vNn3TQ/npAKXCEcB60pQ6wV
sFyDCpsN0uoeoD6Vh9CpS6+/cIlZwwDlXv+KJDEjhLwThJsID9SxQFygLQVk0F5BcOSM+6ThVmQL
OKfa3EYFQhr7J2P2UkLvwLN9Zo2GB7jktOvteL535BgmgbShZGWLm9f1knHlqT33nIn2AdQWEKfB
m9ZioUZE2Ym8H2JnBaOymj17dcc1azHpk0JbwRQ0cCoSPYlczp8Uc8tk8YTP4tU/5nOSzGCf4NYl
w/X15zlv7Hc1PTFiIY5nsbGakSybRhnbIPX9h9MT5KbvihMS1V6b//U+eTmnSDkCENY6JGr7Kxrl
sY4sSB5lwmByaPXdLhjSWFOl01VFCCZeMQInpJukB4vjlyucsPIWyw2Rev8qG+LytBNXthtg4wb+
sGXjXgQs9v3c5z51JoWHGGXwoGRohXJCy7kezy2rulSGCSksLy8b2BjzUnNLQ5K0sA4X+tF1LOA8
aVgOj65A/em9Ty8PDeKFk1l5hauEBr25q47/44cu3pDePiVV1E41FDFblLSGEVE+c/D3zGcKdXKn
bxHvMyQmUC+jJcu/yIbPzlBTb5sBenJKWhXXkCUB/SwswIIy6Lgynxz0buwmvnNtvAiS6dc4iqM2
9UJd+dsg3JN4Snk6YD3drx30DFiHPjtqdBHFNtapBFZyIQr3H+UfPv8PH6QiJxUNiLJKUduIh+qD
RQsqHCZpQ+3ZnyVj6CNa+DsoSTXaDxzCOOysLdbUpauUYR0suTTZULNUY29128I2PuTJtJVY6pXn
s/5LHsgwKgjnDj6IAe9VF7cXTKYENB42oeHMYKJ7/UIWcS6tpXvjlMMdBNc3cOkGfHesmH7cJ/f3
9dsShYXtaYDO2rqFqYdMv8vtUS4ifQgrERJHovL37wK1Y63tzWCYxSAQwPkfNcCoz4HpN5wb2DSm
hpZM5UNuumH7OYOn6arraM+6eKNRnHBlh4ECW/QwiRI0xU2KttR0EaXVBxktkRnbyaXSziA3FG5C
vmKiaSVZRrhxUSNFKVouoO8uVfUk7lHUJvjjSU2prXXs5Becw9H4bRfcR8inx0skoEnF1fLffOhs
W5mBxPUfzE5HSSLKkCcxDNlgNWlDcTW2iWAs9q3qIOM+YA7AUwNrM88lx8076N5+5vyaKoRBCKlZ
hTdpee2hwXc0oxomqzP0HynuA14XsVqEhoJs25j5oDwPbfzEXxmFEgnoBbSsW1YDPAR1nboqAHNf
YRzYVe2/47ubPv+GDhu8pqGE9zwhUpNeYDwzRNivUYD8NStxOdUTo1/V2/BK1rVhNNXksEpkCAUe
ho4/iQeQfIRBIPJdcMhsYB6UPKXCKWPj4FUKDqul4E6NyzAfBHpvzRyuA2O2sv6mZ995pDN0YDf4
wLMX2m5XoD4VyJ/PA46x5w5KDyxZwfxE43VK5yMuu0g4ntRRPLOvN48Kmtk9YGzLMuf0QnZPCF+z
Xxt423TdO32drtL41AY3YUTQ8Js4lBHvk/5nT/nDRzCxkHwwDzaB4WnZXf4kJOEhNiJ8UWI35nPR
oOODTxcMyrBk7syHWh2ABkiYye/kgkqPIKQBMZQYA4liMQG34rGqFXrSfQW/86sRlaR5O0UeTUwX
agKcCaE0grcAXSBB8GijXkFJdu0BDJOK+cwxdTRK4L8kgR4fpiM2C13q1rEuDhIhUakoKuO4p6G5
mSRTaDif6zWiEQfYa8tamQLBIf+e5ybgJ4v8DcyqB7njHFh4QH8LQcGfIXDq9EuBlhPswG5n8f87
Fw6cb+Zv3p6yn0Vc7rCy39rfkaKF0QuhJAFlWvM7jS31qR6fqZN922NZNWfURWQM+hZ4qaaSt1XI
t/sra001BFuZs0rYKhUomLvbJ9OfsmsqGE7D59Frp+GOQBKc5dPASeQPcgiPwWCVTbjxIIg5o7on
yFJWUPMnLpEzHqDkYFiS5av3hsqjKrqGSz1rEyicIBO2JjNG1w5ITHz9vTjk0e/8BZ0371lZUOWw
hkU9U1MIM0NVxBpY1hjADDH1cY7a6vnClWi/mzVwkjW5I60CfbSC9A1JEVayIxsCZP8xY4xzZYfG
w+u3jUGeJxjC3nDRv3GBehDv42vrlebZBPekvwg/fyn/Ptn6RBoWoJMXHQ1oemc+KWiAmPouwRPb
Yt43jn5m721iANVoleQ8SddJfbSph5bnfZ5xiDL6czO7meLNJyZkG/Rcd8H089z8fPUXprsmiM1B
DuEQR30hb36mHCY8aJK6Lm5rhgL1MlwRiQICttaIhf50DdFuh84pg2eqWbYN/0OTZ5WEMfo60JsW
yut3f9IVhKF27zhkv2JuKuVUCin60lv4IHtLgqhFXS2LRkaS/3BUFxgNoy8i3W1xP0D5cusOHpih
hmtg6F6p/aD7SdcGsQHU4Tl7eRXEaiT+vgRPl8iRq2PfkpUaniYoHmrC/2BTn2Tf7u7+6DcAsBPm
OtfhhGYJxaURFDosZTgC9XAHi8SOBEy+4LkYYmwAQNoiFxMKUy6h0M5eU/qwzj0Qhk0lO9IFmqg4
QJTI4edkBvguLIOwERrlZyiHXmHn848jXuJC6Beu3HtetKJoSGmuWD3BwUMq5JDTOmAFxixIPbPi
9VrBxRX54kv/E3cP8SiNiRPbDb7DFwd3n6vV88TyxYR3mcSygSbq3T/SJkkC6uT+UXqm9jy8YIhr
YGP9YzdwbaZ+9/GbTja+3o+5tpv31TIa0Tt9cuu9c5yHIZ2/hh/jZG+AluxzeszXNjLNlW22k0FC
GibdrK3Gwr8XI8N0GLBUkI5nF49cNgDVi4Cxbbp6+Id2UyeA7IygIeoT1WKzsT30Jegn1aK5MAmV
sHI0PS3XGwqiMUnNmcgm1q5sRzn1bRx3ZR6fYHPwnt2lvGB5d/YaIx5xXJgjlXfsnAJietq5c1zm
8uAWPVQimfUgBNMPG9w6lbhBZC+q7QTFuyTZgPEtzVfuoR0nyOFZnU3uvEvfY54sNLvR5TUeE7/R
xRz1bkaMw37+WGvOJfCAm0U3FeLN+oBT5xfLFOYaQyxwvH3gSyeqzoqLeeOKp0fIGUPEdv+fJlK/
ZAMpv2ZkzF1sgFzceQtq6sVw3r9dvFzogVb9Z1jNHKT9zWPhrhDakFUYH7L+hGwWOhbBslb8lIa6
76NmZxB+ueNVpN1FTahu9xwbtlcn1fQNK9/RE21kHOWzETFhu+oEjzefrd12iiSgL9TBLMtDeibz
Rsv7LSmxuLvNWYi37HWIFsY6tkOS31C4JEtanH/OMzm0ex/Cq5/PQtH/J6UxFu/gwW57jg2OIm4k
oeaOa1HUKIBNa7/QfhYi7UDOXFcl2s/d8BII5PZfeJZmL8tzH4RxfxrIhWjTkyhEcHO16iJH7EGI
DwT/hoxNaYOu3P9VrWkFy0bOSniQU5vHtJEpozFJCwTl0wx24BOh3+ertHIs6tSzCJAxZ5LSVU7C
7P+SpAEGNExm5BfxH5MMNxU/Fbylf/o63Sd9Cxj5AuEoOxGSdgiKupr4Hz4J9SJfZGQzce2T4Qwo
pC1ncsnoq2rFA0P4ezabNY2a+alhT4VslEy9zDVlTk6jutLasJJ4VDPLzmoyHLEmwt6oSsIOhrhj
AImnIwPNCnA6n0VoHPuChI4dhTqZENjPiY+HtDE3I+jUtw1K5sAjMBxkJKiv4IA/W7FFK9IfHxnM
gj0KHmhEiDFVCoGxmyL5DCIqAI4/5sTecPSH31GvBZUC+VazQOZ5YmVQ3D3UtRDre1P2Moo7x1cV
uEwg6+02mYhzt/6rxdlIMpP0BVqbNOXhRSER8ckbD/JFrk+9ijstKFa0mSdwYx2JgARyefY1kMuj
nYQ1Oci2siQ88/SbjDJ/5h2n0JtLosry6QTpwQQ1OTvR0XKnpmR7v7NITTO6QrleUm3bbD6NzTKX
Fa5CW6fjnynjJy4UXLS+TBs/WMy+Vbm8stj2Qvv5QXyEL7F884BbXLtpfK9D05N30s+Oqj/z4iHS
bO+9rt/P0f6EPUZQXNG0OzAXKSJWkPYaxLftejEsHetfxCTWJf2PiuEYJ9gMRiMPe2L8ZpWu1UUo
XffkW77X4ezM2fCEiCrzOC+DL4r9H7Z9cAOudbUAzN9lJQ1KfKXcOVe0ZBIZ3eaQTn47Q03sibKH
b2WC2m0tPS247RYWeL1dCbXV9WNHfsP13vZyMSO4RXxIrkNhsiRRxl3n6do7jeFi2JTJk2phj7kd
uvyi7XwT1UxK+GxNclenpwExiIBlf1FnoyyeGlvgiA+L1C7MIp7MGN5X+9vgGte8Ua51fO7OhL1B
ijiqdqcN+f8xSV+s5e4thX2LlL8Ra/qq0LL0i20xp6Utt7qzNiGq/hnVn65L+4Vtv6GBEdfdojuq
fgWer9IAiXz2hEBPyOH1sKQU37Vji+iKtPQBB2OkRJiXMB7nMf46K+UzDs9+R3yf2dEzQD7dpfTy
d3Fo/Jy0OsCLBBzdP7gVEgXwTQlrNs9bVc67X3hp/8yNSZNghqKgev9HX0AUmoq56zb3V3dawPZx
47o8MWe53tAKvyc0FCSvak9yI/Dcd8UpD2QCdv2qxRcPqIu13tXw8Hic3X/Ig4qcCjAkdmi5wxQG
F6hR7e23+229UgBUGEilJCvBnqRasV550OCz2qrSwbCMut4NmVV9gkazcrnny6YudDayWdY/Xl0R
sY4AQnqtipnv7Hank3AkrNNLHAl5bFhXg/Csq+g6uNbfS8MHAkA36lq8JblsxCUNJQvQk3d/M5uT
0VcDhVar/Qv69fRz+tI6mF26QfHz/JEj3Vp5EXy+2YiqR7SaNURKZatx863BryGqtUpHg4Db6IIU
yU8YPZKqzoO86UGVVtvD16ThdsT9FmPSvH5Vng1sKqzLVVV5QwQijebbWDuZFWMp1GYZpO42Lh4a
9HEnmrASiz4u5tTfQGumxFe9zA77Ao89SuNkIy+Hh/23V3g1MVaLj+lIXrh94CDi8A/Gl4RiNqrQ
6qggDLcvqN2Gf93iHiZjSIFhd7gQmM4h1RZ6+5Z15DO5Q6wtA9IShRdRjk7vGsZJu1fl21i5C4Hl
u7oSyP1+obe8YvYHSV3WyQ5WFkkWqRNwY8pmnLC+5/QkmQDy/DhU/KGF/T3Anef7wCR4yzZsDRRs
mZaWqMgk6Fhhu7bCbMC+ALjXeFlxoETGRAiS5skr+bnjs4tQoo0DenWouB76pnHchymTa0J7iZuz
PktZqaVeaSYCmLQE/l/oabjGeXbD2Z3ExkDpggq5Vi7avXHELrbR9nhLPAufudnD9SqMYTmY9v1J
o/534+DZn2z5GfjS+Mn0poiIm7E7vnOrsuIHRvk1X6S9eIQOmzlDDWkptFAbaXcrB0k/v+ds6qIC
g1nSgXb6vhmXRyMWwQ18HLINT/kijAipmb6XbuXuQh+ex0HQkiB4tqiqolhAibee6HbIpc2tHheF
K60JX8/5hjGGZ4ax0ux/J+Iu0TsPs4g+7a4odaHRx4C0xRPJ8bL4WY3awR4V+OE+5pBEEL3uxQXs
DqMHGFrso8gZBqp5N7lbNNLWqw75o5q29Bf9LkZ2t9MsuGbDrrozEZlOdFKKmWJduBOweuEqek0M
jzTryJVjZA6YL1afuTYIpT5CugwcnS3LrYW97K7BatLd3xUiSRp9AqVngbhpcvY+8O+FdctY969I
VjsfEU1BSLdcZAIpUxr5bMpgjMsMvsRKqIsJEA2eW5nwoWdfHb6Vn6AFCgQdOOsX/jaeT/XnedBM
0VEbabD1EuYeO8V9em4PheI7m6PhDKxD56EQYuFEQF0xsY6JdWXcRxfPEuQ2Z1uS5juHvqcRKTZw
op9+YhgO/leAt4vvdlf3c6LBhMSTjiT70QUb9HFOntACUBPVxYfPm/OyGd9b55B4ncQaDF1CEWK6
XQGVbG3+xFKyH64e2wupZHxTVTMznkLaSTa1Y1QLNr8pPG1N3Fb/8qgdxK09k2HdRtBf2GECHqe+
9jP1cCCY0pQnVvqhHevl6kiU6JksCfdP/AefKJYmN5Vjml06kQ7qNQXcSA2rJuWKt2KBuX5tCmoQ
6SZt5DiM1YTXvUYQZmZCj6J7ocGPorFA872I50czVfbnHCvgZuIY/Llxdnoz1D+YohQKvjWaNca4
PoZJN2xONGEexvcDR2E3rbPgAx8kqeHyFHTazeofDpUymwsr3YNygfGxiaUheIFXL2JUFEfXF5mA
5PrzDWIH1N0INupIhWdPkc2zU2gUmn/rxipjZK1DhDTHuE5rL4NYKUkjR/EnL+RjVU2Tb9oT18RK
uFuSDQOtF9V2OENLXGZVGkzdNXZTYnhlU7f1BtwvCsqB3V9FLDodHJyuQXyipSLd0vgXWUJQJ9em
tDaScUPOXwzYVJHEm6i6d9/+jp6B59XdiE9zQwvfVpH4p/B9LCk61/rbr1kK9A3m4gpk0fbVp1l/
MFpE3hzu0NLGubhlCMQ9Z8w40D06w3KDQedugk4ashTDSf5p0bQskYpTCLunye5Hz9kxI4wiJ4kv
RIrYjqXSajXwlQCJuTj4V+ym5kjrYWF6mJiYsm1MH7u5/hnAcBHvHvU1Jn3xInS1kvK2hRLHcw2b
kwxQhh6khXY0HlIuwip7SSL1nszWKORErl+Mm0XCDCALlnoOXTMMgqHQvpTLZz8nSzWLpI1IYzxi
u1I0WeDa75YDA7tYsxoYBLl15fpj8cFwkAuiF07IpV1gvcP1HPYw5xTcVeBpc5yUov8PxQguOE29
P+X/6gwroJdJ2H5Bign1FTRNTK/kg38ebZmb5DDbMbILW7R3eDvha6N9Y3aJVkQT3QQAb8GWP7DB
Mxa5EUXyoJpwQH/sdT52HmSFnaFRWt1qNJcsM+tHhbQpJaRw+qqtliuOtjUFCXSY0YRQ/lA3TalV
jAwNS39SAFdpDD06PoZUK8Kv37pkDHYqnj9X8DiysCkh+cc3GWRu1OODM+NM153LU08djsIjXyT3
fuebrlX8d36Clgaz4Q9cFwgrZ7G3ZdH4L7ZEu9OI7Np32oA1DD8tAHnDNU6CW2aZv6BHYwyszxOl
OaEz0em3WorHSrzr+7+XgVaHnZniDMTw585kKZRkrqEIBFjZX3wPEHXN7mPuSydGOZ5FSAfZIKGH
LzhrOPTmqfLxOjgKJxRMRkVUWCydbAIxxOkkYP9gaXt4X/IUbt/Dh9I2dhW0h4ttocFv/QTA0wyp
d1E6YtH4BDoUBRqUNqxsOxvbCtqliXydar+Kl1QUlkgTIsHfScPBlBvxMl1qjJrHV6vUwZIiWGhR
uaB0BD8lHxKjqn7isHOxtzFkRHeJc/XLubdR79PFq+zE9M29s/GMy0N7pnw9A8r0Funnw5DpfCSv
PUOgnSjlFbt7bGwni43G1rw2hlv05VwWUeWulHhlGpJ36VwrjL/yMHDKU057hl50ZKapuXtd37lx
/famwgCTTB2GZx7nOe7rjPNzyH8occzcFM9RH7ZKYjDKTP8CMFb2whCcuWBXrgFJo8UXLKq39WaA
Z3cGNTZQp6ynwqZLR9suhcvGNjAjryis8I4MnNjF+zBPIcDAnI+1lG+EvUQqdQQH3jOyNEiqCIqn
OZWog/7JMriqMjnMu16F0JJpiJiVjNQ7w27nHr1GkiuTDfHYEdVz7YzYhoxS7J19IQN3S61mekox
7TBEu9Xyixg0UNe3dnFRLo8NjElon9SGZ5VzOCl8kKsl4qb1U+Ou+ZhssZ0KrqMd7wxhvkqPm61f
/KRUZouqDbkop0FyKg2qFVVolZql65xV25/a5/WPjR+VTMUZPhDF5GBIKbeFZR8306HWJ9jYAvjl
729spRwJgDtD0+IJFF/2tdL6G90+69FBM0EfX7cxirAycsffqe0yAlTn0UJYN8iN2pkzyZy8zZir
Ol4j6zJvYZv7ElliuV9SGs+e+yPSruQ/+BcZtFaMnhum+kVtRmLlyL3iBS/QDOjZwWE37A9A2Rrc
rUj0WB56VzIngzh9TKYJFTtzpTLEfE11DKn18hcN5h8eU5662AyKbKC18M1BtQyJtEUFvfeVD8yq
0dRtM//IyeaYAwIRvfBnaRW2qFOQW3ih3Q7FzZJ9hmB8XyoXZPl+OijsAMNaVgVxa/BZzznkxBDb
PKCx/5Q7Adp6js2RXHI2KUjjy6TooukRVUJyvSa7rLbdZmuCs4mwEFmEUZXTXCfhhe+HyTFLsGZK
esyn6jZUffZiqv7moWwNsuCadqSPjBK9EeIesH6ftWV601/HvK1ubXlhAAO2Q3zmtbFVbNAVozqv
Jj0T8qhq/V8mdGtEKKfjWqHqqvB6BPEqNTypNTKbIOPSk+Y8JIvycZzjBRS1DQq33du+4cAOl5FF
G9fT9m6nRtkLFain65Q4gJJxiBVII/IKZTp0S51eQN4kBZxlP2SXhGQo5Xe4y0PLRftINRZY92/W
Kob4zYiNK46jKs2gUIAT1qIGyyXlNbXLGOby9NffJ3amWpWqIDc+f0BYeaB4FTLIZrOUAoSzdv8/
FZjZbUracv498+aWEtgPe+9UOPFK1p9e5kGs6t9DMxNMr4qFlgtVjnCLR3+HEkpQovyj8QFZMUA5
ZJFMsuRDhm8hofJsRTDTJmdD5d5KYK2jh8qdbHr+dd9JNmaJ5XEbJGpKKH67wdx8rjKNkoRc4abh
pIXqoSqE/AH4etewvqgSYSNC4vReBGm84hPcQ53Wk2PJzR0EpmGJhqz6yHKTZ2j5lTn3I/s3tCuz
6uojCWF2iUgfFqLkTOOQ3FvuiMp4d2p04tatJW5y8Q2RuU4iMH8zmTQWDHKsK9KGtJki378cdMKf
OMumzEcSv+LlFoRGjg1VWEHCIL/OQoP5nBZVyJBOe/YpZtPftouMR4E8CyobFfXHhrSLy5kPKwRe
OvDlt+wKpY6gQtMt9Q6KyVxq8o02alwDStGMfeEBSwaGfTmbJ3IACL7AN1Q0ApqeRU56I1frEbMF
3AMMxgAuTPRyirt7lhwaA2Gy7KQ9oj4k/IXHb1EQfzzxs1yw4rbc0RNLsRH3eQo5xpV4t5d0pZa6
M1hSShUPngASa1GASYWi764zd368WEDg5R+yiMVYhDH0UMH3uujWFCG2tsUtL+kRfxo/NRhIQAli
0vfMRXPpXka7VvuOp6QQkWnPg0Xai+6kMVM09lVhgWg4hd8fBKJcuuXLewsNJR/D7ux8QEBfzIR7
nTkbOHKrDRFIY3V7BDga9+rupA08qy2Mwz/+vhmm2e4TOydJV+VbNGNH/rJeXzGb58wrNm0iuJSq
3m26o/Jj757TeRnphgigioZ7sf51tLqF2bPxjOuwK5/RfxUEYRobQlnNC98tV6L3GIqbM/rXsU30
ibLRZrxR7klb5s2qEtDOt6hdSZFCJ7WfwE7R1jjfx8Pz/vfSsck+BUMQ8eIbv/NOytg2Nc8rL/gn
do/2F2J3cngK9NbKSrYSjzpGavgV/ue992kr/8Oz3PN0ErNssrXCdnTdyfHR2f2ccyVujiVY+94C
TGAbpugbyIDvT3BCVuAat//4d3iEB/+98aQon2Fa2l7UU/p5NjoAChlWMrzeKrED4eOx2pIpNsx7
qWVxixSqxZ+m1LztR3d4Y2hO2dZkatvANsTiChnTIEBUy+3EiAYcWAaGHwEyERRgvPPmH2HhirHd
VcDi8Zqu5BnlcRM4yQpwfC1EWZ3p22kt/6k/+HC0qigotsg0XjKHDeTn9bU5SHj4qTwoDQSB/mhQ
CzzwjOmvXtayjikq1XFXDj6QctNoFA05eRcYXicFEtVbLRklRKrYyBkVZlkjfFq2+e6ih78hY0LG
iR5bX2EGl4fqVU/w+DEaaK0vZT+cVORf6r2sFzJkJ2oQvgcCvWV+WMRGbrbP5eOjHt5BLaYKLIgC
HJKA9PUe8h0Ru++Eh95BrTa4vO5+nxL9XxQAc0PcC5UkIxhV6MqoH1PdiadvwQwh+WIiafGKRms3
Gj1pgvSjlg38GV74fZR+AJ6ZJnBxtcqduP29DKrIz2ENY708FbDuBtp7vBrNokHlyhOfr+TtnyM3
6h7agtR3ClvOZqt4eQT2QsFRy7xx5Q5r5y0C4i/6BRrpn1TjHmiariGcpwiuLD3QFmnHIbi6ZKu0
MYyfb8Vc42whbgYdNYrO/jOHAVkgLiYfnl2ivDH4AYQzap9ApiGVBg9TZq9Ak/R9ode4Mgqf1L2u
bSUseRcrwrDlbYCuaYeQyndqi80R45G5GmzUptDyYZLhRYy65/OvGBCvyb/nXrSUsjiSToBNy6CN
0RGH0F1H1cFUq/JTi5umWeiG3NE35qfj7pdXzPsfo7DLZSupg9FeTiUPEfqVdoZ8FZA6rigQDUQI
pXS2COnDstoslbKgqlXQYkSj3osvAqKB2bf2BcVl5Sa99ibFHc4soDjaI0BrsTEF1becJHZ5C/Hn
Xfpd+DNbp9vdRXxi4q3sFlLkYzKdXZlgkcxkrs0RluKPnusrNAYKvlCXttcxGi5A2QNPb8Hhqked
fJ7AMoHoeOOEuQ+eQC+p/oEUskd6x6WuvrAhfctp1lRnMGZj4W6rvq9zxL7zolKvltaEWi5wCa/u
XSWq7bJJQchffiOrG65LpKXC3ofTxuIdYaFZyPkl/mXNnwrHuEBgW8yDyb4P7xOsgvGUGqxT+TGT
FM278ftxQhU1ku7R28WV60Nqqyop9UwZFJRajwcGpJSacOprdG8AsA8SonIRKsYS1jsZTBVYqJ+H
MNOSfBBFxb4c192v7E1LMBcQEDsNKe+ekPrDOg7/f5UpLFiOeT7Hg81A/XHGjljIANR2OO+RV6Sk
BYmQUU3lVwAoDQ+vAOmyU2G7Nf+vPdrwQnSF96HcUo0nczTjt0pSJZ2/yMN2l1PoWyr8s3Tk2a62
f9i9Go2BOSEzjg4ym98Di6kcHJgNHRitTWcGl8OtYhMM+YT3jsc/zCTdxci7oRv9TgwyeRuUFH2J
udISnYpYK8rjb2mmFhfDney3RGddLKZTT/WZF9fczMCheKWYO4g8jF2FcvPV38ibZKI2diJ3hqhn
29QFBTnlVzEedw6jiIL4tz+gTBhCrvyN5P2IAnHdSDQAU4/R+kyuvgEVPLRy0fyXqMl81HUJgxYO
3rDek1hzZA9obVVVdY9SEfAtkt9S707ls2l65NB0CUdDkj2cPda49N6YajCnNXlL5YvZoLMH4Ek5
Y6iXLXQAndG1FcOb49tn4g/RfNGbDImhWHHPxS+efdTY+t9blzhP2d+//QoxW5/yI+s/R1mYAxIf
8YphvA6+toEkdxBHigkXnCOg5oCf39Bxqh89HzhOD8k3ImM//JrTkJVBOGVpO8otYA224MIRcv4N
J/0bVUnM2y1qA0GwbbJ55nAtlgMpEfyk5Sne1CZHKSV307C2m7V8fb0S0fGFmc9YmFKjSZt/MfOu
H6dTQ4d8HGlpkipQH68koopHD6DKpcdHefPSUVbKmancsYRSoQgm+hemvvFhs1xZw5SKNWRCH7wQ
SUrNaDmu4ix89P+UoddbhwwAuZt1Pw77VvGuec9NKDo03WE3c2oFd0FtPPYpXS7boOtIfWV/Bw7c
hRwZkz5buUktK/Xo6jzuEyehyHj9tY1CWG1mzO+wfUscjSRF3zB7v9LA/EOOFia8llIDL3xA633I
2PTvPSa+Rltm2574Bca5RL0MJ7hz6L5411oyhc5q/0Pu6FUg7oV5NbTIdAUm5e1OV6f/36efJma/
BH537MXo4VauEuaGVfQL7TtVsSEUJIU5QxfowG72zo5RGe+Sr5NXJ7rJerO0Xs4zB6/+r5jMHimE
TcCd5dgmUmYiJk46JGIOLyUcTV1mSSMnBNmwocyH0BfH/0hzwRMm81RBwtvNFs7ccz7XL7dtnQQr
hrvLO4E+jte/tXgE+sUDq+5KS1z538+tVzzjf/fZmUUCboq3GRQqfCkGyeoB1EXXAkKhcwoW+cyW
hWNt2iCFeO6HrbR9fCM4kTO7e5NqBW9JhwpecTKDARdFgUOSBN34cYjJqU1/U9pNSOxMrkNHdLpz
Hpu6JGQ40NkqOI+c81SoE7O+6fh7gUOBkTdfwMtqYlly7OeYPllOV/JdKiArjIMcc+ay30XBluiw
v2O6nT9pAf9JyqsW/cnFi9uiVXyKT8YeQAJfDtGhIOQTwhb/0pw5CXh3iZgmzWEnGfwomR/9ybRm
EjCbjCTQy/MM0lq8Ptcy2B3ElInx8WQ1CwnvANpcwhoV/NsJdGOkbTkgnwCFKT6xtCk0gb2BkjRz
g0Drft+KKRvUB6SAy+fXCJx4gpZd/+/A8FbqAD3KFsM52ONFGoBbaWIEhdoIxk9ykRv6mzKhR+NS
9/YDKzWuqpVviLIks8g/hjEV/wEahRZ35jI4VCjwc6QURoqxLLziPF8PwQKstStvNlOG81mKc/Fj
DsjrUeukAka+4AiUgJ4qRkShpQJI9GSuIWDYsKb17i2+r5QuZXEHChxKK/4qc4MphPb6QuSsjWde
ykCaV5ELgZLvm6Sclgkiv8h1MKFjVgFIyQ6UgNfe+85ursZMPWROoyfDyndFwzANzpQGk3Vsd5lH
uCVqBMpcZ3t2N9xJ+V5hF5+E14M6d0KaUsNFFbI5nReYlpTKiwY4gQB/03/bkB1DDF7fL/FDoNlO
XRFsWPT1B53tfhz2p0yZJbp1rfziVy+j/uwi22tWpjD34Ta88/jt74z6QuDPzcO84aUn7pHlmIHR
MgMFHqTQDSu22SM/l4m+K3Gwd+Kz/R3HUZcDMb9jRk5p06imTa2iMbjXHwM3lJoa8ckZOKD4CGXX
GTyuCDsAbhL0g71SXrWSdh/yzuWoO7kVJHytctfrKMiNJ8FimAzq/D0n5w4Tg8WPKtCZP5rtUo4d
DVE2h6vFpb5CFarCEe9sEPIMZaHLiayCdPndqBZKV409GYfmj/rx6XzN7MRNmiXtxImOECgsnTvw
cNAMsGY10woUhcixxXh6iC46Vl0GpZtJ0AVnGIQWw0p+aQJtBCDNT2WDKfORRET+SJDePLCpPD4g
zMOvCjg1G50nFnU5zVTcdb53qTpkT6OVk4+wG7Pz+eQlDs/t+pDVdVMcsP74lNb3DwW69csCCCIC
PwqDRE4zoVuW0YkvwQ/pKSBC2KyLE09NnzUUDlSDMNXe1N1ZKtcFfCxAJgVeHKNnFXg04OMRJscg
eSeyFsrTbZF74s6bvxAZU1QepTUgPHm/JIph3CmaDg4UNRkP8zJAZJ6p9+ysVL6yzsUigmKhPgPu
+PO+JLX3X3gu9mWCElONQ0E8EDkedcl6VQ21JwDlF9JCrlQ3k0nIln/TEc9jQG0LncSnk1xvV/+V
jqhoZu4rUo9ZohFoWlhkeiERw/tqw+TSG8s0QyCnCJDarpP3/BZ3BHEqfOFZ1uiHVWYFwLPjRWZZ
ogcmI8rWHBOglGUCae8EBE5C9kQNMm4D63CoU2UmApxhJOSuhcToR25bqGRAVocJPQvw0DNCJ2se
xZQQsjEiSrJSM18/+HPSgUqYuwk2CSIx4Q+NplJo54gZi3WBC0slDOM3nCRT00d5sr4wNz1bwTSL
l+DZJ0ZgXMnGsTjKp4EWVCwdSksHNxadQj6ZgeWji9WjtXgG4LH4aoT4HIqNHALYUNr9+11wjJH+
YF/eKvh8cEP0rV5MTYW7V02LGv4eiVjeoKBqqbUQvcL+epusm4yQZvehZUbGWUK/wKv9M8BiG55x
8XnDVq113Yo57jP6vdUtx/ln23wAiE1MrLXgraccVHdTvcVUZXB1iJuBGsgJ8cIXlyg8s43ygQJB
WOOSfgpz/pgDGO8dwHJz+2Y4L4x3zU7Fpw5AOmsfk3kjfSXYGPR+yIzHWxhBqgHf+ApS9LP9hR0X
jnxtj1Xs7RqMDpTM10F2HxDOHttxiajrn9ewnNt007dJvgrBYg7pn5dPOzgMhrMeWYSqB9XD6M7i
/2apSEMkQxZPESv63cNB64mY5UOvbybQsX/gr9a+ewFxJjBSVNxco6hCYP4YpAa9jmQXRPws9TOM
rcHnvknql7s1isTan1dOLYrcvvLmayIOHcWOxv22icquXJuaFO09TzBMjeRRnaUFnl91joPaoKL4
1VP26pmpqNyG1sW+KSq7SJxGbISzbyknr618Fobh6CM05L9rIr1b0teVmYW1h3Jhkx5SRLz/MMBa
UsOd/LaMiuY4VjayzdHRIJqgmCuIc9bdzX6tIIluEAZNj+H/Z8bHHvp2VymqLw6M8x1p04FZTyH/
NKuRoXUMYSkAKEVOErfYNBdtf/0ExMCJLpfiZ7fs5/hhkPIFEFLugJsACBt6egbClOagyi2+sP0a
QLiGmB7Z3WMoj2oAMDkBGtGDTGh58ctu3d6RM5sfl6mcWKJvOOOUiIW2oI0E7gpT/KJG3N/bXNr4
d4ThT3iv3snnQRxfYvpUPIwD4RU0LGOkbBq8Ex++x3Lzmqg5ANpJhiNveXSF7nKs/T0Y854o6gTv
nHDHouGU55QbzDyhd+zKwbvgGUfLFaN0/OuvyLkm29Hc7sD5KTRCikliIky15Yf91rFfF5VN9H7l
Vm1b7zC58gQZVCmkQfCxkiF88CLhXFPS5LzFckithPSQ11y4wb8IHnVQqWUOt3DgQfFI8k2xRrSw
uEIdfUvZKGDd46OhBL6w9aJoko64P5eHDNm1SQM2xtdyzcsPLR+q7WCBPiSlr2ZPQVFZbki3qPuf
4G0RPs4nc/EjqByEe8HlYVcwCjl81oJXX6743MgbBRNoamKzZxtKtKYKfTUWSPuIX59ZcdCRb9YV
u7UQEfwOYtEHAVn1sTVdXkaH7YOGmrmpCbBDK8SNTxxlvdLjNRSyrYovdrxg/M7VSyYeG3mzVilN
78liKhs1EfRicZw+jeVxlU5rWzPUcSDdUAXay5XUcIGa1Uyo9Yv4G6RdaTE0CAlUXV2EXO5tLN/p
9XGEj671ARK6Ednie5mBfqFpykWTLj7exMXHQw39R6wy9y0sIkVUnsc76GcGgRF9nphSJyZdi/+m
R8xRJJlXuieGEihxSxfOo66kMfYLw7TXEbrrYdWR+06UBqYw7WFEMwBDofKebAPs3t2blIJzBjbJ
3xzUx7P25wYVJhpwbBHnsSDwKYgvXNZHpR2DTT10z/ejBVcxImXDp0o9Fcj21BJVGLtDo4knBnRn
5vxldN7GcSM72cyBiiWhXCSyI+4lViJ6K4llXZ7ocTbcNhWDhUqhlBnN84NkoEBkS3rnNPKnxlI/
4bWf+7TEJpzA5MLAdQF3+LEMFSSkm+15Eve6LS5Qd7Frg8MERk9JVB2wq16ly8xHhF5WdbID+cj0
yh4P1kiqMT2RjJG9OmSIVRK1mWFTtsm07o0mLTiild+A/gfJ6ZC7vSP5vWhgFrYM7y1DwY40la3z
90wfsUeqaoJvpKz3bsX5YpZnvYXVXkQfh2egJ0w/8WbBawxJBFa+Ef4TTDUGrtfJZp3rHEhLxEnW
VH1Q8ACS7W+joQF9LUzS9QxGA77ZP1tBp3UIvlJ3UbZCYO9iFUSlM7POsA7mtqoSy4UJ1vPjqioZ
8vgNA/unZl+CevPMGtiaPpPeAY5PfOC4ndM1Z1/T1CeBaqXkLaIJZQ45RGC32uwQxir1flBly6Qg
7Q+cPPttuiGRDCBSNZCqJpgLYMtkRpBmUuBeJ7aWQy4EZHDBgaeHte7YY0caPKIkGR4NiIAb3q4v
lrH9dAjvlb3NX3N3Ekq1h1nV2lJutGVkycBz1HlnyCxVZh57RrXJxxNfbk2a5lIKg9qM9+Ccnrpn
DZmBI9I6HGIhVod9OjWU8Fvn6L3bHZ5gB2rUVdj0mQCd5u8Qx+gJa6JjYOCNCpWyhmV4zA7NdZ7o
qhqfSRe7RYGmC8oDuVhAj/7Mri3dshGwaz1Hmmdi1QvFtiR0X5Zct+1303m6q89R1uQpOrmCE64a
cz28lo7ffrGoKLtg+mQYaiFlxf05gJUYP4fR5jrxh4D38w/rMgAGqFo8YeMWUKmoUSXfOlOiBPAs
On5CTgqn5dv9k0gJIqtnCp2Ds8jbMHEJ9NqlaB30vXpADGb7Tac193mQRFKjQc674lzOA+Gxj6P4
Y/XJX9HjXofjps9P7m+Sv1AECT6aP15Xh2HvkyRysgDESWX9Vt8uTdgUdfsRTo+ccrPivBDW2upV
FEzjwmvB8fhFNGN5bK7f1V1Q6JlUrr6zoy80s4Vt+DsIERF8zx9dA5zKP3aQfWJRJITzflCB9bTp
2pxpEdUD8ipFrnC1bp1M48fhHfC9/u72HffzrpEOs6GET2HDPE2JcuOsmOnZU9FnqOEw3xRArbMF
1exxs4IUd9wpAYBezCZGcRuCEnlt5kJU2WxGWPeHKcFwOFEyWb8wSTVzzzRkeFT7VB4HzV406/UZ
xga6wH+xFgEuR4/LDwpm8TPCbN4o3L43tBRPTBiX/4xqzcn18o0MwnTJKkrSCibI6XYLamKiBWcp
bGmft0ccTtZ1qfjMcZxk8DXO6zzGY3N8Rqjy/KARVquqvx7v1hRqtyPKqiQt5PJeYQZRWik6aD6S
pJpRRnHuZteDsjgWbznQEqmnUX3SPkcDe4irspCzkF/lcTrZQyuLUji3khUJOOUgh6ojcbHgw9F+
6RKDq9KiS22nVwl03Rx37obC4b8fFv0BiQrk1eikZSJm1XZwMNSOC+RjqGWCY5SqaLR3XLGTMYmn
bjJvJbm8otWo6uixQJUXDkVFaUvHzo+kPMuRt/PkR4c+7fke/xSXfpeIeJXKg/7QwSs5vBzKVIvo
CdMVyYiCDtJhqdc1BclCwGzvXG0O64nYNhdabcLiMzPBbPl4GXf92FEy/xY6/NbklruXwYkqGHrh
SA67R85EAdzJfUhCr10zbV0K0+CEVR7f/3Dv+7QW1jYn42BU6SRN1T8PS4VOM6w8NVmOzNnbzBQX
LZiY5LZSzlZa2prc72iT/JCajMfilY7Yf/VqxFPmlBFb1Qx2aXtWv4wnFp2KEVOPZxd4PoN4NZLt
pUeE6Eatp5185IXaiPhoQ3mU7a/YS15xxpdtWE7x4jSDGVhBK/uQG2z6u9zR4YyVp2r4+XZuwvLI
dkjjjBSKYM5p6kNClzjhvQ9XrKtGc25qdvryBOxRIHC+gA68CLxvzyCeDSR28gFXixKVzewmDLSS
U6h+qyUT7LrZ3Y/s8dIH0cdmufyL18fJMd3O6W//XkEgTJZFjcsenRwobuHWQhV0ZkXFVEdhjzAp
MN58zpVbhpvTB+DlDELrNRmM/AuxRmq0+pr/+32rob7GP8QNNc+a3wEZM8wHYiiOj8C1K+q6850k
zFMbuMf3l7rkHaf5e6AKy05ydyoDzo4cpM03SZhAvaGdw2wGOzWuZX3I3tUQzVADaXliJy42+gbb
VRyrDyiY1hGwCjXsayMgr/YKAcI32m6rM/XORFpgS01bOMZ4YstaFNFNrqdCHCDbK5lPqSYEQR3L
Xz2bhl6WtRTNLDijfzbj0rBrx4rLZifRcJZkQCmoNnycjhoQmQlJZ5bGJWKFPqOYEDZmOTzqGsjN
aHDUVvAPbNBom2vviaNlvLD7CFDCFmoAq9b/TvuioTbYGyYl0UyYu98Q9W3TrzEHU16ze0NGFzF6
QwCfyN4ltWy+dvcif366ISjPZPjfbIaHzzbeIoV+pSppXV8eSNY32GuBq+xCfjgpYr4JMJcADDx6
zWAWri1v++r0Ipm2pThBKRzxvTHPqhi2bPJvsMv5dY7+feB/aULY9MLbEiHnfQHeR0wpjg/ZeyuC
osVRCvQI7O6zOXucrZl+cQg5UUpJwCJIFdH52BIANgmbsOnhJ2dYoQfH8ocSwhsBFPgOWjx0d1xU
RDAA0m/d6qmKmxcgSeLpHGL991tCgVkk8UvGWdUwFHpgKaRCAyqHjOSUBSeCsavmQPbw8yiY+2q3
KIFRxc8ORabnI+xHOgYCP1Fjivzn0lZ9XXYBYOz7XvjamGyJqRIuU9JAX5+8i3azKoro2S/yqxFA
1DzxWK4oejg3Z9jv/mwGaUzBRqx9YOYr0kBNi6XY2Zb2gNKf65KFct1XkXTdR2cQa124kJv2sg95
BewtoGPw7XPW5BptvzELg0q9Na8lGF/KhGsZnNx0n4AC3UgBkw00ybMnFNuM29EmI4PVI2TMuVam
kMwonKAJuBpPH7n5oFRcUVA16s+gVkUiOqPKvEYQmzSLugmCBo3S6DdPWaGXiNNPIRvgZSR2XTUc
dN5zIEApGnkqYQulSFT1kWAkeDt7Jv2cXdQEW5bG/+swx7bmMLU782Rc0CC4bAjKv0V9aN0ykybP
3fK7NkzeP7K9ZcOKTc5nsQsdhxNnARnFua4GgKHkzmQZzILIcLpJ+R/7rPIS6jhLBp+CEpxZUk2a
33gqmXRoDkePNI72HfSWglTTwNWwvurIKHRaR44Yx49+haWAlQMX7pORZPZoCRUvE8XzTpg3EyyE
zLLjudpXKv8BUyvcQmoE+sjfa04f5NWnmMzNGhNGoIbUPQ4WOzSBH3miYHRPRZrA59PR1rqG1h/8
azrzHjg7RHR+Fzw9j2zpPzBdu+nFz4jK7kbc150SxNBcm7PR5Nxc1TgSVMViBkszxReeA+WZVtOD
pvDk3OuKOuL6nrlvJyJ7+vGuAPS5xl+GUEv7EoAuBqDAC6RfC80deiS2+bd5fotyFoFWeoVm+xZq
YZgrKpO8HyZaDFnxVdwtXohxLKxPf9Ku5iP5d6l6iyxld1pjBKg8dU3/WeoKswQBrQyRT3Em2Y3C
pVHseXwnwGrA6dxOaszSMkVhWJbKyGpK7uDsH8nn7T2l9Xf3ezM2urhFMqnA/i6Z29rHhZRt8v6Y
JwxyySdJKnqrN6AUZsejBmbOX3ezrJVGLMagW8j2VjwLC8Sga7fpSP3t5F1YRAyNfzpwamw8KG62
IPdC+uicUwKjnqdoniPTdvi/0HA6RkgzV1CBEqikGUGoMVBolmfVDI50adlAkNA+pH/KLSEgUSYS
TT5f62F1Cii9thZxhd5s/E9LRd2y14Oo4p2m3BeXVwzIvz/NjPF0o+scwHJlEpIikzyPGp0l+Zec
9kMrPwID5t9QHxd1ICSLGojLgyeroMrKtpYEXqkv7/t72WT+UfTc7am3u3HLYEI9au3Sf3vUbC/o
WajcbaBY+kuvD5hGrymoUcJQE0c73rOKnq4WxEBYNpbv6dxIsfe8mblSDyVXTGO6s1IcDZvsBRVZ
Hkyaw/MaQloUbKy7WmqrADN5s2rpYlLwiIcTKL+5fmogcaIPVL/lBE/Wq1qwiZO3YKaeNVyiNKho
W1qzEAHuFLDLmefqMQVkvX2vhu7VtkgQ55+82qcw6d5Qj3XV0dblJE2DQwYJlOnoQZlZzNfBXbGI
Ce2UFw8ISJ85KoyCx4t0MYo81qu9/1Q2p5f/jJ56jjNlqfajLar09Wk8Uzi+nuBIWTS4EXtMTVT2
Y1XlZC8x6Ex8j86NlIJpChvNV0IzRdcUIfhDr6RpTrqaH//dcfqmS9GEjWw46Qdi7wPsfkKJ7A9H
uvNXwj8PAdUTYmSMGeOCM8x3I9ErskPQDwsOChxHbzs7Gd7rSEBofioXw1XhRNOGX2ojZrviqKwF
5KgmZr6nVY4KT7kQRSuBZsXutWbb6Mwz4wMiQzgpdquQf/LwSLmf3mZavFo9tnKM98nx/i3SriIp
txo1+WwuODOWKzw7VbY5P4wSEsu/iHCPScHVvcuGBf28EUiI1N/sc55NOoBJlbkOCseB1eklWAMe
kSaIMu4jJtTOk5WbeANp4xlZ2AU4gln7n7CkKBpZcRILF6DJVKkhAdgNz//BUE0/0bTkg5CEliV2
ZXMSzOX3OFuHPg8WC+vA1SIZvpO1K1FDI02ZR/9v+RQyMJDWTBkRmDudpYbY3nTTJPGse+yUW65s
oiLMsrCAJW4OYkTSeLW0YYEkzjjgVzZ13ABGG5JE2I39K8MlRL5lExWBLxORimqjx2OcwTCuIW0a
o9yc3EGoct2fRx32O/Ul8JrGlz7ebq4WfrzpK30+aMmlsy98h2oX8pjW/fZvryw9qESTH8o5i6GQ
wtDaQcYbWEedNT2z1UjC0h7F9N194rn9OoRVkpi7yY7Ff7lGuFPduGeXcHSUKSdBGxTF6KMMdkzc
ghV2YXx7H06eg/3kTsJdL9rWpOMMClwFR6NejiJpGbrnyttN/d7Lq/mPnqCQsQ4y8cNOQuA54x0C
b/olAcloahoydMisav83FBBKc3WPiYTK2j+v468TmOGEwxdLxi77AMhMJ/7OQPo/yARKnmTV80i3
UEqnHv60w7z7pPJae3sbI8kSzbn8ZLLxnlkONy/S08l5y89AQIS68KGAIs/nVoO1II81DF8UWBDV
/ttTNtezrK53WVYHAUE5oLtjN8ZAQrF7CTutpkiqtCiinR+fYmwuJOoYUNxr/zhiHwaO1osYTPkQ
ZMs5OH5mNporn4CN7h6Twg7XfN2z/uGbuYgSRIPI+FMdjKbXfO3nmGQR7xOtPpGAaP49puYeIMab
feQPveMRoMh4EaPlEO8nVHXk3TzVydv9XNGD50yPl9mw/6BvX2SRyhDCFsXttbpz2jmhXeAUI842
G/GFi/eV3kC+8et5d/YajVNCN3h/5KdRgybg4tfnMgdH/vQ+AEoO4GiQ1vP8T2vfZWpYLVqfkbhe
PinDJSdKX5Y9Lq6dD+Grf5BYb1qSP4UFYAMcrbP3v/o+zt6ZciIDP1P60FBDnyRWeU+QDavekGZy
i1rr1I+x18Ya7Z9oUKDtPPsrr1EVJ4NB6bIn8EfyCEhH5u5qt5kcdLmZgcCvpiCnqfQbEmVRaHq2
p8bkkYlSYA3Go0qnjyDHVMPBawx1V/C9cNzHagEIKJQo76+rWfljSsXgj0/I9X3EKL+GtMqsFCUQ
o+g1ccQTaz/0wAAqmapdsAF3XzSaGU4q6nD/tprGk1DcIJV6G+VzystshaKQOX90OGAs7tyzQK9O
sCuf5f7ayhMWGxYTZjAnGTkvdfGGhkmLVPf6MBQHXP31d6TpBXznDXNeb2C7j+W1UerVZeH8LIa/
uaBalHzlWD1AIk/5a3Btl4HqklRi/52Hye8KE8B64+1rpY8Lbs6lI0s9nNbb/lJxNL6eTJfrjT8Z
sf6JuJCDzEJejWjO6yNZLExWEGqJlMSxEBtE4F8CdZXOM1rCchTui+vmLR+WipLh3/BFbnE0UZJU
XlQy267TN5QN1lRx5X7z+Ojn9tcnXBkaY8whoOz5Ty0UNfwc6iW//CjDObJru+4kd3R4Pr3LWzvc
2In4ua4CUaEu0eIIFVCZl5CXwulcq6YWc9VmhtCngd8GTMLm2D6Y259mfZf/x92lF310d01HB6iw
PA7LIdQxH7KxnjH2hRRYv5kZFtIM7Mv1fsCuPIbzuq35iRiNkLfxERzRkZ91fUoSCUtmSvltJcRz
l5fBnWx1pwttWn5vfBMb4IY9sLloaij3tL0hT6QQm7zczreCfUcRfIaJ3A1mIvo5JTJsCfA/WDxF
3TSn94AkXNJykJlu2W3p92stjTwDeuMhSAjd4SXCp8erRJ8CRhhx8JfduhnSlSMAzlsmrWFe5Zv4
Wr7ImG4IHduU+eUMM1rB9msNrv1TfbzY8B8uXV+bKojUK50t6yZstvvsM9i5pROnmDLsKgzrUx+Q
fVlIzbDDkuEmhzOdb/SLurl2Wi/UhVcGirCRg7ZT6vRJcfGXMh4ZlTTp7QMU7/8H7eFJ+0yzehp+
O44rM3qMAPjCP13B3ahH/Uix4ALVvkruMru+1Dz4qmxrluTFTvgIgCJC5toNdTSKn3zSKh1odtY/
fDrLHc/fKA6YU9eA5KmoixmiefZdKm6q/mEvX15V6PQ70urYIYD/At7QeyiTUmBjZ1IovAId+Nrl
Eg2Vi8hLISKheCZPiyNMgswZXjJZd8oEKcPsgnjSQO5aCdUhIMm8mP/U8BZvCTWB3ktk0oAWWv6J
bpkWXhFl/KxW55gNCwnYLPZiCT41ON+ElKTgWuet616G866ViSDFcYOm1bbStVBg+t7JKTIDOz7o
7VD1wj1J6IfkAHq7+hy1QP4NkzGqYzyS+FlZduweuQzMjxkoJ/PxQb3rLf3gzucOg2mr1cMVCpXd
ixWO2lUuuLk5sfm6T2zDofATYnd5zDh5qrkFvKZVq1gokdqCfJZCeN2hSydmi34fm9jGX/omJ9Az
VdT0+fZv74limgmuTWJJDE6DG/MVggXDt/wE3fOmpmIHguJY2/sY+bTDJm4BIEHOLfQXGkL33gTH
nqdxBkYYqKROAVpeBgfPuK+CNh2/TmXe4Yiu5jpyPs520iFnklUYJRzd7AK6qbSw5xrXTqDoNIWc
IcpiAGJ61TbAEXqkhiga4zjiF6xZUh0/fe9AfCVhmCmrHvkVnGmHRTQmkr7TJgb4ZLDzURuv70AU
zP3U1WgJuWicpl2DZhVUmz89K5/W3UhUDkhwJHqzkk+bvZ+bYgTCGnBQpea2T1qmhRPQgM534MLj
O4YGz6QEQn+p+8VNyrIZfJYJFfmFpUuLh3HciEE04SsbddvMPUXU4rpBr6rlHGhadyrW6q6vJ3dK
pCwJ/W0eArynUtI7LREc936h/0nJd2We+ut2gSz+Lzyw57WD+0354YayKlFeX0A0UTDqjJNb53RH
P/o8AlHy1i8sz7KbW+ljbBdA5kgZla2PqzASX0ElBa7azfB2Xg0n5laLngUxA2gwmGYkYj8KawPj
2+xsmF3+/ziba/mO+XWDT7Q0X4ziMMShjmm/wPchfU2jumyRzjEn9NgW5zdjAzNW7RpHmoG1ASfg
vAmqTHKYmzZFKcRxeSU66szJ/oGwaQ7MYtryRV6iV1uZRiaWY+xrtkegzwYlxUl/lXLcvgQER0Z9
g5N640Yar2y5V9m9Nw4fvoXHkGXoDLwltsY1d228Pz96EwGhdJDWJBO26KgyF1NMguRMQO4EVrcM
YAO/ZVjro7GPZn/iaxn0zEVghjuaPFgMeOTgtQCR2BFksJqvSHHIpcJwg76prjI9LYhKaQAFQa42
kalarW2gskHPWKipL/dZ5b0ilvgfYTD+jOvedwXAJrkG3uUrXRHw2BoLMsRpXdXhmaF0MUlo62Ga
S2W7NCbmimnbhfRhVUUl/EzeudIKDhINm+jAC+Fg4o162wjpTNmmyxHDwTrFiAF5yZZW7RK8xxHv
8hJKx6+uoW8fuflRqWPI2Ht8O/zY99EuT0JCp9eEzP8fs8oVTlA8yA/4NiVMqTO3iyM/wcyyt52I
gH/3/09rjvyDKy0D1Y6HuQTwBljEtD/nI+tQLayClUhiAbhAA5e24UZbSCHZ63FYaJHSUyR0FG6z
wV/iXVLYZ1VeyQdt9WpFZXI6YBFBp3MsdykcVN2AErXi1+OET/rea/VTFSfTVp7qb5dpCUK5DCpu
10lNIbVl4F7dTPQdhZDwDQ/uXrK3RPxD/m2JXzOresEhSpiRO/Epjidx1ne5xUaNZhK3OsDkamnX
EK3MIbaQtbdg4qcr2+h3atU3eaf+L5erEpF3FaWIkB51kd2NS+fDiC6CKKOBe1ee5Ufe6sReiFS6
VZ2GnUv+PI6JBVmALwwH3a2FqFMdPeJQn14+Q8cc/k/iaAF41Z/qBLTTelda1AcF/9bAZsBuPR66
IbwvOmYmKjajIcJm8Gr9W0YSIhBvLVy+nPQckd+rcGfjMxNXsUlH7LK+w62qFhUEOgKd0RQxvYPE
+HGhVRNOiy0G9toJahdlCsUr8mfSAjEwQc/tJQNC5xl2WWzZUJYZpk2o9zdvme9uOF/folOakvDC
4OjRSVuXdFY/TaTW/v5sF93ASqjnLUhgPHgJPTWtzlu82tPk4Svic40eTpg/EggLCtxpci0afQiq
jQ+QroUhYYCneLa5Ed49USnbteFNrK15psnnbVitzZ5cFmXpAVb2Q6/XXpkGatupdYLwaGslRgMR
rrDszcQUOLUH4iFldA5dcJBp0Peie3qwpwI7F/JSQrAH7cO84AJf2jQhOPGCKy5v4U3XL8JTgdsS
To8SQPIVK6vKs/FRQu/5unraVMYduk+W8Qn4XK0Aa9zRqKggwwxQPZaq60hLQwDkg2jmGxSgnUWU
x9Q+xTjb7FvPxzYF0B96hQWR/tasGZZf9ifPF4cxqfm9BUksPcFnkrRz/SWfwWJNfWMLyqxYUCnp
Fuko/U8MZ7nl22WNPPtMCf4eTg9r8trxjkVkNfRQwGL7HVAnK8Vp7GQedL8wmDialgxowL9fxPv+
IOtmWHZckP81e8uxbhF0PR3AhFjGRGJmnB1mUBeXseyKfGGRcUlPkioq8FgNAokoKAFUm0fauoKg
yx/XFFAbXV37YxLeRfkfsbpgztLRfhDyx5JV51UIYZXveZoamOlIKdCwaJcPYT+gXCWVAUHucoOm
B2YF6wYuaBKfeg+TwjO++2OyarSnAfv8J/Ip0wW/74+vpno3h6+cQNyZhxMokX5AUEei3RGrk64s
BUqavuIi/g7GAQLdS2v/oJ+X+4gI01zy5I8aSe3ks52nR7AKG3+WHll4H4efzcKbJAe1W5EGNMSV
jNkLt+p0+TtjJSSK7PMjn/hwqN1FwErPW41h3ak3wHU6GeWSEk6Sddd/hvK/XOo3XsakM7LZAkjt
sc51icwfeKseOQJSXDf2Ipvig4rT236M4+UIGwn6viTDa2N74VjKF37/P87eTWat7329xkiD+kJm
t1eenoopvYZdZZOgtP2NkJvmgeHzMQ0SQ4G8OUDvJbr+GG2QglurVnP3GZTb9GKZKetIz4HXyGrS
+GZKm6B8fD7df/fvYUz6bt0S6uPenUD+JyMlDZEm+WOumiTL0TJjlil/MnmyWDSKnJUIGtZAmeQH
QPHSye3f7ylZYqEYpfi/YJ8RmU8taadc3EthPWFjRU1MoyOtZxOX9rSelkHtp1dRGQ2nNdah7yj5
Cq08P++JoHebIb4Kuu9yHxshQZLhshKSo85lxU1q4aPEJALQ0cSK0o1czl4TSeJfuY7v4m2RGuB7
bJZwlSNcCbLN7v/FmIr25RLEVoacCo6DRA+mgCOn10sY/atEcnpLR9uegz2S2waEUXW6dBxBp5o7
NZWWE/Zy77h9G53Gok2M/PWUJTqp/PG3krHdbtwnZL92ayoPXHxcuA3ltOVhV5y5jWobpwAFr2uz
xvX7F3Z5YwvTs9D2PWyuZEwnLB2s9ckizaiLhZ+vxT/XcpUe0iciH0rz1IZFL+vxUA3r217aVNnF
xErb2xztRlHu4xFbfi7TFtwzhrZw3CwSSp6zDiyfvlHces7QJe1mAfd3AoL09nR8+LAp8NoJcl+B
eC36y05Hs8U9/xqcBHSdp8+XKuBNIeBqR/tiQhFlj8ar1klefPeJEgLPlK35GNEZIMaaKO79FsKD
JSym0iXDnXXuf0/EpiSEFuiO1GlWcE8XCYUqX18obwTtAim17rKs+K7g7HU819GDa4889lCHAc6h
ZjelsMu7BPBs2pYEajzPI+pkXHw2qMOoWNdgK8vY7ptm9eTWPfnnAStqqG+VS81XCJVRYkvziI9X
2Z0bV/LrjpURmoqP6DXzTkf+U0i8V0mg0D3NGJApMjlKnFtyauonGmnc7ruciomsd1KEphG0Srqb
N5Bi8hYqSxuTyV3ypkxLlB5TBlDOyWIMADTxp4/Y+M285dx64ZSL6BicAKIDqtHHPsLYkz6Wl/jg
F/EPw7UviNTfsBErtW0lI7lF7oW5iQ67dSWJyK6d/U9zm5XcdPCAFyuOrtsS8upn65DWFUP6qKp3
+WxuiEI5/Dsi5Rj59HEEbT03WYelu3FuqiBL3JHXzIYWvGrdyJjPTCQRNLr0UPjDSv6OTzZYXY36
+sa10xxSkhz87ogWwtzVnYgM0D+dr5NnPeU0jjbcLnHW8AH8+3Bi2JDC6gsNo+O/wb+dYvmKmayV
NTJHhzBIVGklNTsOIv8qXmTXGVFnN4INkaqPgCj/tGHTcNTnxU2L4ASqX6YElGo1umPhbSv9+iyX
UOcT6yOZi0CqgoXSbqj8vBzkaSr0oJ35p5kEq8OTuPFcK2Ke0ANyOeujcLLuehfc1ljXfpPf5LPY
kjZwYj0QThbVT/hNEsltw+B5Pr0lwZamRm0Z2FOzvb02qsbWCdL8/XywzGYE6WG3d6aaWY+ApNq0
tLgq1txNCmRuS6LFBURkL+c/pn5K8g26OGOaemE/6XXkrTxPQPWiiFQCfeDlpL9QQANCOV6xnlfd
uCEfKV0wet7zXk7voS7Dp5Jn8KMrlNcQsmEfwA6RG2Od3o9GVevbqTnaYpWaf+JhKRcBSeIoB1Ii
8+hiyTMljWiTKyj0XPGA4yN5+NabIVDT1xKgd9xlBcfAWhNAU9/GIuNiBf6sy0Bh3nx0Brcg5d5J
iiLsCMH/4BUFAnf1vVTbdRAw/lWOZVB9kijkh3/jTpVTYL72w+ErLEdgwHVlvB5lQSIGyMWiSNP/
d5Y/GBpLFKRxK2aXi0jaYrQs3aiogpFK5rZ26IbT1rhnsROpo6PTthF9f0xJ6T3F6aQM6JRMysBH
vHqLtOqmJZ+O5zjUZl5/IZ0I09N00ZhPktthrAc5UGCvTw6bdqjxcIKNfPEMcxSMfySN9mEVEG0F
CGSGjVUKhStdPZAibFJ1T4MlacS64bIdhzW88tOQBW3LJI1+0pHuoi7bBpRWVNZkSar/sVZQLQ6c
ezzobK1Sd2K6BCAwWqAP20X7cMPT0E1ZtjELupUqpjMvDfj+YtH/nnfs6ErCtuXqvd/mnWpSdAAi
KHneiXZtwSR1A9WlztZIFcNQEht1UGzYf+2eQoxBXVTO/3Stk637LrSFpj/Zj/DS+TdFywe6qWjz
KwPropVLJkyspGLYsoZ4ybVj8B0GrWDvdSC9vqf5zBM4EbUZ4WmgcI5csXKNnkdKy31h3VHWhwLJ
vlbpkpwJY/RRySAh3lWsO1ElGBOnryF8XzKrBZB8wiV20WiWv0ChszuqhbIAcpP/j2lGaAutOF2f
C2zCCZ4bxxrFVPXXb88BhaUglCh2eexg2dnIelqGZQlrSzG2CrU+H84IQxC9Hq3EczMibfNz5uO/
4cyd0fB9VXbRzY8TGUV5Rv2CJKPoOqhnpNkXegPCUOYjvR3n121gH11cLE0oYL6qZzIVRs+FXkBu
R+Ky88usKYwMqINcFByduZFqpyhd2FBOCbOMIpG19iB6ZXKDQs0zWKpymqLq7rS9JXfDr2RxfNah
GL/COqsZDe2HF4X9g9DhWbySoh7WznKzE7UT9FsUoy4woGXMqOMP2FZftGQsOAuSQduDn6lTxElx
VUTsJ74+Au2/DUcVTsRWg59yA0ZBcDqqJhCQc3XgLsE6hDRLaotWA5Y5/IWlyNwTrRjDpU6yEA+k
lL53jBuCvZh0XouSBz6TVdD7AoGSLhFjubIL+f1QAHBf5CmD5wE+QZ1EXso/XdUTOl7Pa1NDpesn
N4HfZ12MZy0ufUuHehoZ5fDINzHIopj+Po6hvM7Z4cQQPceUMx1z6VCIL0ZyhkAK59gIIDUpNKoV
pELg/LTemVIv3UGBbq9+ebXjhaCmCvb5HqGURDtihUkZy1fAUVrhej3DSK2YcDTxGah8ETx4Sj9h
vI/uGXQ+TI/9TtROtEf8xFyObEbkwjIZCo+PmwMetoWrSXyuZ2RU/KnlS20+wFNNSzIA09+vFW0l
ciwWU3ONhgWH5MEaTf0ihP5TJqko2pRh6OmQUvkjQXPFfhUgKA+EEiq1SnA22vZ4KPfHAc4PA3le
XUo8fmO6HIL/7OUtZm3PYn4TrwKAEmJDtdAbuRa6SktnUsIHu8C0uVsATXBSemidy0ysPNgXJATI
PoY180ZNQVgBRliqUVoozHf7f836ZP5MVDv2jiUUs62cuVFGRs6NrINx566h/20XhUGTNvivRapB
TobQW1X3ZumXw3yZFCg4Sy/4TFdPL0pwTm9dfaNQPGVu+OjvzNTGTSRQOGg6wg7Zz9NTOlCBWU4k
BCAHqkyFTb7vPtlrxXkc32eCfz9zCzZOVM2pHZhBB2hBRIQ+czkpalq7+Y2pbJEeiLMWsRsiyY76
sHkT65zpxJOmkLh0PFZbM6JNfTXmSSu+a8GDm7hlOyfqh+RmA4AzDpuGOcXcMhIBwe+c8NBA3GZN
mlWi+71FMfkeosq7NEzpznL4GE3alsuvkUSuWbo8xZGqy5E8HENguYWK1GNO5VszB8/BJH0/rKiG
St634DygG5krfqidWrjuHZfdcbL2REa94gcDZE+M+3pBkSJVtNvOVrGT4TF2sWInvqWB/REpbX79
fQjcPvoKvoCPLkzfAEB/lI8GmsLHlnRoiywrhkn9Z4NAnKd+zDvRBFnRrRumA4bwLh6odecg5g5s
eArRu2lVdcMCJzN4w6rIMw6t4jyeOKgdYPVxx49uK1QN/k6VrYOyflWaMgKJJt2RFc1LmnMKEfny
dE9yZc/wsAgmy8Qe+fTfTCQIdB/OBpA/8+Y0UqFSxkA1gKIMLafp3BhfmzQj/3BQVqRkFhORzxnR
5zGvVnCVO0nvkuMj/4gTC1zi1aH89DhAiNHAo29XmrGIgOp2JhFWwYkTUxd/BUCoa7sQsudc+cqr
5Ta0ddb+jn+aEVJrlih0AfsMg9gSZyqeUwphyImMNEti8RV48BIOyJztsZG1DwPZnfmAKP+JK6jV
BsoJgWNopYLVEiLe0XQTeatjPYSd9bRZIXOxP02iPwAKIoIzOY0MSJo5DKXNDivYFFbqHcCV647B
aIkjwDfll1hyi3gC/AOmap7QDIQ9cjy55z/HKQPfpIUCBTRERBJVpdLfNvl33zkSaYWXpaCH71iN
Bw1WYUJqicdi09lRMgfsqIzWqtwaNrpZdlqiyfaz1Fbll2tRhExVisSXqaIX6p4lUXwyngXIKMYE
Nu7rlP4MwErJqIu0B0l/KbF4e6QWVSzbgIOWG/ZaDTHLQYc6yVsKuiu+pAt+CXxHfQLgOcMEvEhD
i2zGrTThy0fW3JapJtXWI3uCeRFCjC6FHfSg5rl0dChN0jqfTVPdAkI0sWick/XXsgV+Dwc6eB6j
aoyBIwI6YM59De+di24AguHVrnrR17dJ2mLbVBZ7LzVQMQqlyrD/d69BEKCw7OvnarbHeHpdMQET
SqfLJ1epXDuhmz/+VC3z/CtNRLkWSNcpCRcWBgDvlJUo8WvxYXW8EOQlkKPkSBwPQ0xjhmF0Y8CY
GLlkeDNvhzUrJbqYeX4DKYkDUPTz3BzJRWhMcOms3hISauODbJgAW59SJxE+9zHw84XkfzJ+tet2
Pqc/hFQN4U8cNJd5QLE3OXdR88L9IzAIm+e0gZkklquHaL1PANdcWmyenU+TKDpuSNbJ+ZlsidLI
9ahpOBZDuP37EWz6qLmTqCCFNM0+4soRgZ6Lfz9A1+ttOUiruHtB1nXveEGNSJ4f6xIDuvYznmzK
OE2Hgt4TbqKhsHt1YQPB0hspR6d0h8xeueXvEXWxZz1XhViKGfRNMxPxT/E6HQmEaHNmiiWwTjjn
B+MxTBiD7w/gxYRrH3sR9ITo07+TbJbVmlpEMdRXys1sYxp95HGJwf/9ye/fzYVMnLwt/WykNBYS
9xYvxr6NE3w5h0lrV/2ybJkMZHGbF2PwxTzeaFqhIm6gksF3aNt2cWlPIIaQTOIv9o6Rosmyr8Dr
8udZvcmtUVOoC803N9+Pz3NSGE9vv8hGV8oSp52OoqeGygIp2XxMIGS9xWN33CYC7MozxmxioR4v
9NVDCztkmmz2PVSwgW421DLJBiDtkEMoW41g4BNOShOOZjXL5Xp6F2/hwzRV0E4kYFUXWALJzCnr
SmXN8jrBFBoDRJZ8i3h8wPAqX5R9+w6BJAL3uoRrAw+HHPgAyy+fAVef6ym1ZTg1oSrd0Qa/A83S
j9hMWJIDqWe1kynX1zz459YvWgQ8O7nxaEEhqOXJuoFvzqfflz5Amv1i7zwwewl4+zeBDBG2RVJi
jLwOrly5LJBgjCF7d+ZMa0PAj2WJXGhCXnahPWgXLcnUBdvS2FFWFs7xhLh4qA+AnVsSDEFmRchV
t6UcT4wunHsGmkqBpvDVLbgH4zyjie/uKR8mbV7BR6VOmFviW5nnDEN6G9h0mSZWvQx6wCVsRff5
QupADYaWyOYTss9m/YzUrN8czHqvXuPOkiDNHeVWPgfAvfb5IaVPju6+9uTSD1wTWDThNlX5OmQw
UDX3a9dPLaWYkSju6QPvlZNm0X5XGF/gdC3uJTctwoJ/4VO2yasSBhrKYJjvzW1nJQha44AiQy1K
VeFmGvOHX5nCUBMZitPQ922rPK1iUG4VfsLI2cG20irfnzidWP6QBJuF/b+Pc+vM5AOhnZuXsNu5
3oR9Yllq9u8Au6uvtgjpT42pVfOa0MQrk0iniBnDsSG7OpfVAdcRdHK6J4gJCmYKM/ri3FdelTfD
LEhktC/5ZzLRlj2CVjNP4GR0Ku2Ts0TwRsDsDe15Ynq5+L9jMO2NjDjY3g2Srvc5fG8ErTOXJxZQ
MReXRo9tcYSyJ2H2PENMaVGZnMvMr9JW7f9m5GJJr9SPu0Srca/DLLGaEMcCPkbWeTqVdhwqKoMT
oEtoiIe+8Aht54MLJFc0xv9CGolRS4LK912MCdhR2g3gbE6XWYAFKz9DhegaV1XEY5VGAEhCRqd9
zLJCriLqOpy68Q34t2/02oBJipNCPW+6cF97HF8RrrLMEWEoZqBAuziFEpv1ixJFsrzSfFnU6ZDh
7oXQXAzwgimVKkO5onqy7/IoIgS0MjzM+KSi/mdgG54w5Y/oPrDw+SBmB5orvMwkRnp9ewZfoB8c
OSGL9qZkNroDC75DIlr/NGAWIy/cDcOLt+xW6OAJoj4RhH54dXfoLx1Z1peRxnCbFgvPYLMh69ft
icP8dWe4EMh1D0EfOyCYx2nkEDC0xOcQiR58nHsU0kItbXXMgjZFxtK3kor6XhSvOCFzt7OxGT3u
BtH0A+bQv4qnO6Dsdq1Au2hNbrHXyWrV9SCKi2/WPuXl2oXLv53kL8XqJOGLpfWym86i73rkX24E
BvCwS5pwnDcNcFiN2ZNg9u/eBY4SOajt/tx142xv6joBYhFtSrKIGiDqC6YCQXwElxcwW3m1R0Bj
FyuHEl3aJ/opdsy4KbjAzBuAter+TW4TkFoyWVbeOZ+Tcp2c5kHM8ConVXCbESGC0jrdwMgS708e
pqFxOy0hFkKc3Ar3tpBOnhdaqev9pT1clgsRf+hbmeQK9BdBpPxYgcdp4t2W1amwKxvuBUQjdK9F
sdMMhc0JAMnPylWmVEOfB4lTf6MIF9tx9LHKBv7pXAoe/DZ0g5wSVxx7mNELBV+YXo251/zJWhps
K8YnyymcXRfTlSkkjssHHKJ37t51U+idWJ7VfVd1T+VFO34xrSI/PD1DnStp1EtPM6yA9pLj7bSG
/LXNp2n14zoiWlpYFXgDwTOLbAWOyZmeLcs7qUwPx3fgjVAhKsoZ46qRk6Ny702Vo9XdI1rjvHcT
lnK1hm8y4aMDh2ehnXLT0JajOAZOnPUNRWRwJYxLXeIEOztJ0/3+6Qn201flsezIpAmY5YTZUg3H
m3MVodaL4blLQLsnAfFzK6qnlQ+L2uvXCt3DOzgS6Jv6gHiXwwVakWSFuDY37OsDXgL5V08+QkQo
ca52dtT0jzWkJEaDHnws6XQaslujg9nMQa/Fk4ayUCcis4NlayskiQCEPC8bcQrakSxgkpmptu3J
ZhkulDoZcHy9le4EDTij0wGsPL5pvQKxV3DQ+DTA7gPbgOoI8Jn2jFd2mqJikAybxW1MmU7yWKn6
/c5tjOYZPUiposkCg9jygYc+EHWuRlEzWmpJWqCUbxC0fgIeJ+zs1EZgqdjui00q+k0Qv2vmGeFO
sMXFSSR2EUp1IHOHPZ9/V+XfOVgYquIj7wSis3T5ow95/OMYX1UYyKwKhRMAZI8nJHIk/owJKjxv
XeWC8wsWlOumpxswUWEYOmAyoIT4gG2cGNyEgxGefQGl160Egwk/wuy75JwagjVjyHZojMpefgZW
dwZL6mdoU98RTnjUdtNdXOfVxptWI/AoA+/TgsSQUn8DWwu4OuR01e5Nxf/GRZ+7oFqBsTbcWmKe
vwBCvnBJ8/7myoIs3AQrdZ4qoeHt5fxygPVya4xzzw+LK+Lik1wE8WY847k/SWk0t0yL3aOkay8Q
dL3+jJFXeNQI5B38A1q/Q7s12sgZQVIhmzhwz5F2Gi6zuVUcy26iBPAXaefRhYI0UrWMbnN8+vMq
ySfN2TSNvosI/jaZqf6quCfFBwe1Ab+WHwwssiQko4wG4caekcLRe+i40LcPIOBpPfC4FK9J7bG2
zQlMD6KeplGR3WRBSnzwSctZA+Cijb7bGz8fG+cOjTk89Sl9WjAAwpeu6ZQL17LnAp0tge1qSrGG
MNWoSHlezN8PR4Yz8rvhWoG9i9+kRy6E16/xYS+TsMVL7i58dTCxAHiFyKX6LG8m0oxKq5uuq7iG
RBg8aW0ffLfUvxfhyG84eSa/MhEMpDj2R/BmyjducIiSPhDMUGC7eeRdpGcEFp0IudC2qj+1EJ74
onhjM0yC5lFdlMvgJ3lFfupIAkjLqCRBh0EPZboTVak0xoetbBDWgtqsaSPA+GVOR1P1RlWtlz2u
c2o6vH0lsOvTZN3Xkq0Rd0NJR6EycvZsFEyI5ijL5n0aONhgukvWVjjK5cnj9nMDhGKYgKMKcc5E
JMsQYuiE2K3so2fiIpy+HLHllmbE9n7swnd/LIdyiX+UrqkiVwTigVh2WKT2UWSl5UJwuwfQQY9Q
03xB3NbP7A35oteX7cCvhYFkzVn5dDY2YCxV9G0/sd5hQ7BmR57/3JUS6+ZN6dD0oEGppvT0Vtll
2ies1cU+FzGOorvlmQEkwkQTEdupIdPP3Q9jdzMxUo4VijTXAOMHi+ySoz+3dtDzwsDHuYMAunpV
YHIaceNFw3aJ1ye6ILaXXEijeo4naLPEBjaF3ZKIrXqcySSdqJmMrZyv/xakyPWqRiXzOTrunvdJ
HBM9DCXJLI89tH6jiO+TaTIYYJ0Ftql5VE41B7tbGAQIhV+JaO8ZFw9oOm1xLe3PFH3omqbky6d/
zwswIyzZl0koWSMrkuOeN+ZTZB6IdJcTXkSjB01WIbznKkkdS3yrn2Fz1vNnW1eMXJlSvzWR/Xyc
w4/zHrdotyh0qbbeQ2d5b0NUVyI2P5URef4R0n2NgKb1qxk5g7VS1QPTcbzuMEoUKXxI+uBzgbBL
Ro4FTHsHd0PWBEqcZjCBmq2M5N2KzzY6nfZzPqs2EXiHX7VE5rXxhCMTeFvLdyWNH1Mz8QHde5vs
XV9/IseHgvJr5J8kd7AplXTt6TIQT4z8bY1R1pbSr0BRflYvfMAPdTpMOSCKzgIzQZkmUFuOQWeu
99nkBUf6NVlC2bECv73mKymBa/50DlFUcoSIQOH/46m84xeXQZollMSR062KYI12WUF90Dic9+wX
z67eo/CoXYBhRlj3LIPQA+IslXtIBdPKZwmAEzq6LxHtZaKlH+ShWdXIddLHNOGDQo56s7+jETaE
h9HoQYz+PZ7GN8u3nttNgQ0tJyAe2JyAW11UOpa49jB9gU/64lsjF9f5KfewsbX8eMg+116IGhC7
4zzzI/GQkAbc7z/2+wf7Mr3TPdkeQijA6EZcC+15/pz1Gi1hesP/DIcfeOkbsk4gb4Zf3w6ltkIw
wxP28dzmAK9pXjGbNm/TlOyoA0rwNB2W2LMCqZWRyS5oNv6kC8cC7FP3Q5a6Z/B8cyYGq1pbOSe6
JTFnieRAiakeBhvxQpddJLTmxTL2NVelywWBbwD6Qe8+UUHjKe9zk/Vwbl/55Kgl103pFDvHA5Pt
6TfDpz/b5sqaiNrJav82bxOJ7upQf0GWmgdcvxkMDVF1/7RWL6zoMAz2EQYbO7T8O3NHUzSDxYBD
wGdmMGXfLWvKMzFasHhAocmoAejhVlsSWeQBW0RP3joYxbUWx0BmFKjCsZ2dWjnyRVN+iF03+g8W
l2mOn1jrWsxtR/bk8yQBC0v5JKa0NAzJbfSCIXc79hymzWS4eQ+0vpeqrWOHIVPueLGkbzsd6wWC
AxKDNLT6+1R2MxUR3S/43FCSOje5C3FPPaC0XqzttT3c1CzbOmpJdATGAimGIV490eakAeuzLYyu
vaHsWAIsfPOTqY7qfvBlGekiqCzCADMlxoWF7dmllUJsoG1y80OCZUYkbKP+iYGy5gm7d1WxzuzR
bbcFwqdVZtKv7P5JdRMnCkkusL79Db08wUTks9NJGMCF/jcKXda7Bxbl+P+7pNDNjU7ExeYAiafR
nZRMzM4FLbuzZ0lLfYEV2B1z/tb70GdpzIfEoDxeFWYtoRAEBf4VntuEJBSCuGkOoTp+EZiVE3Yv
d67wyVv2snvcQPM4cfSAz9kIyyGpw9Acp5o4lHXee7d3lR6P3xNDZiJ9MCcOcBjYbAJ/g8W9iaL+
K5V3LVuwtiKIEC4zq41xMFB31UTgq5s/LgJR73AqVOUzr2oPVw7Xs/n1Xod9X3o91xGNXd+nd+rV
GclTyq7PmDv9OLczSYAY7Nqe8J35ZvAXzRcD16M25E9KhqdtO1CaQP8NWLtw6oVKcahTe7xL+YUs
2fOq4GP/CShLDiEjTYyRt/IKa5gjKCjg6eMMLnIsMavtJiMDNZrJdso0LDJSvHoE5Tiib/tgTBUl
WN1ehWQeTgXTmpK+QCnGx13KjJjhSiaIx3WpV7atLWf5DIj/lAcbBEjan0TTuDK81826iCkLbQxV
ZxcpZceuKU3lJ7Z7tnsMjBKQpQ2anxpaJ4+tPs5rRjVwD0MySs8VjsQUPqspn0ZnkFv45zOyRY2G
7+8DZf2DCo/utrVhgFmr6/Qwn93CZG5663FbP3a+52tF8TFofq5Txnjrye0/Pm5rAdYlvv2ndqnn
8WEkVAdIhi11FEmlQEc1z6hOjN/fDA/YshHgvTcYsHQAHPxHUqdhJB9sD8UIm0yvOEC+RSSDB1T2
UfKaKYDJU5hyNzSZAItsnLrwoluZ91K9nedx/wX3lnCR/b7+4Ks++lTpVXoDUkzVv1JX4idfHcwb
OtCqT7dVLydVMyu+EJ/lTLG1mLNXrVtNO/GYRFbWj6yAxZwiVhwXQGNCdrf1ZzfUknz2MbGYIhoy
rxFCU/VGPESpo+/4I8/LAtU0pnxed6zi35rGr7HnX9YxzdA0D3APuWlYekjSLQYH7K6Dr+5dvWcT
LZp3v2R++voAq/D94I8xNXfe2JUigscCKntEoYqy2CMh2hwNBrz0DOuHmnIxlSDHn2UJuOEXcHg7
vjkVTqzfk5EKUwLB539JF7g/gA3/q9T4713pZgCZaicQyHdoUpbDy1sW/EeMa+PCaE9AhQ4XBE1q
Rz7xChnbF9b16o2ubxZAYKd4I37j4iYHFcTaEYYbN4zscz/eJ1eRI0s1mkLj3A3tAIzNnsv3DKgE
68/L3X60DY/PzdMEDmGMS9iej8VV41gRQB/UlVkSc+y9IMKL6z/FMYjz3ZxsEqWVkapKMrGEV0Jy
iHrRRbksQO8JA+tTRnkKLIFORYI4665K7QLcZudXUixGoyvDRfNUaxoIxATm075EgizSJ8m8Gn/e
Fg9DIidKo33IZAG3Y4jKSzPLMJyixAoK1PfIJk18wQKirZmIo7vxciCPyFJXdEZ3QF4aqfbmWPMg
5XLlGRjpyQBhVdKmK6YqR3Fw6Jp+SuztBmcB45xdvFCmSivWqflPK5ph5xfoNJHBBcxNNrljp9iu
wYauOGRgN+ynGkwnNAY3Nzi9vjpYznV/M7zMo0ucJtETJ0RkEenMsrvw8j7L6y8l/GgC6Op5IcMY
gY2A84U6097uJX83LS4hZ3d9JZaT+CL1tMrJCZk28qO0JwDVLDX7YWegjeB42xXJnfr7vfk33le2
RMXbELfR+hS02I7roBYZpDbWMAWDz6Ui0zKwysbvWDenaaoXVaBJFpARSfakTA2M/1yUcTEv+XrA
zKQACmvgwidvamME6Ncl6WtEBQY1pb1zmOvTglEX+AUexN+0GWfoB11gDS/xNxhOxA8GmLTJN1z/
IIfuXAm4vbSxCvtqom8NByKaBKF7WHbiOoe+ufZvwbqCueqy+dltdqmM7quJqblVhOvmvQ8+Q9et
FRLiFLuz6hpO1yTyX9uTZ3dcTgZ7h2u+awMopgqQ15bicSnSHgDlwxU/OCOLuKO42n8jynEZnZPZ
rGaYju6B2oqGWzdaUMp/Rg8ue0CoYObKcT6D9q7NEGtjq6kiNFqbSIaFcCei4/YbZuV5Ltn4npBc
he3IMwpmRS8MH/R2FzZYhdn94MkMQX7Dz4NzpXDaCnqknEyymanjbQ4km+Il5rHAwBD/9FyRPqKv
cRFYWKvoeKa5zjpm2qQCH3xxyPbdlDBBmid9SsbwPvihWdNB51GzElP/8FXbX2Viob9ChCDpwdYo
IqSkP47oknCiqgdnn03ogr19i8CTPrTI03DtdCvUxz6rCzcJ8ZetCXVOcsIlXrE64kmFEkBH3AUD
APrEKuc28lFlENYoPulJrd8seF9yRZVc1xWHWt1yZYtPJJPYUjGufwzMJy5rMIrZ0HyOuosNSNUc
2ZhPoyHx0SCm0u26DxgUE/ujMq0Qqzl7UQoAQfQJFWm4gLSHcu0IvMz/pvpY5IqV7ASzF+E4qaFx
K2vjIWEamXWjiGkG1qibRp2wUimp/eRqSEinu/JQv2FcZSwpcB6lUlEbFKuz/eyCY2DnFpBA3OPH
uOzXdmDWyLeoh4EAd0xA87Cqa4ZHzk5vY0JZU2qO4o5BtnloVGq0o68TOHIlkW2Nf9OjMvCzlYAq
wvkiwrrls+GphyBhQJ0/AC3FsskZghzf/1XbLQFtJbnjJxRJmpkYXoFlrFQJ0TVd+XAcrUmGzrIw
JVqL21wKXErv7RzFURAXb3bYtqazOeSWn1U8g+NfoKvQnj3Aem6DQwf8YghlmLX36oXOmZr0fl7d
wzFnOxmo1X+0nmLwkwhBO5b+h+j0rWSHdjnZ9ZMCgraEW5XI9cXyBcZr278I4VqNzVUjPn0RxXy1
A3l+5HHKkfK2tAaVob90koEBFQAN/hNtWe5Ry+Ucy2miEcGBuik9gmoDmUVAUthRHrd8FyncfPvo
eUDlWa756o3dZVY3S2CUJgHhnfUX/njNMtJP5ZvSHAvQHCWjUo6YlybmLJyZ+goWRQs9c2MwrbJU
vugprCOyg83Hd4ZGtqPH4lUlebBn1L8jYG/1Ix4GLQDpCDJRowdr3/4Lf65EkQVunZBJZyBeI7U9
JRNaS3O2VGXcxTYcvJsKfMtHTudqOICs66BbXgjvG6xlUwVpFbuhuAqNGSVHiAqIDwltbddiY10c
m3faSDQ8YtyRaq2cKSCT1pv4z7qupIfIpGW3/m+oDLTYhEGG40DKWiiNPQ5+5GlCI42cRI8rRSzM
Fkvv2S8GRiuIv6q6uz+GsSw63RQUqTG+XRIvwI1SKsCoB9+AjU6gOfZ/tQYeUCAqzoTXAZ1tQpYg
FyhtWJTJGU2X0T4xpxIsDEJ2+SHdpa8Xct/ie+YRGHvPZHRcF6+/4mbNTlUOvUYvYTvFq/U3N8gT
doBFiuo5RRlkrJwcKkBDv/c+BqjCESkiqJRuFvKB+n2A6PItp0hVKm2l24jlLDA51ZnFLlKMwQI+
2Yy41yL6yfdNpFB4tHI+cwKRSIqZgZuSaDMUKXmO7egUvtnSVUuxX1hFPpZmyiutvWhEEI47xGgZ
sziKPLBHwfoNAwt5zSCNPRj1W3s1DfQGZfbkA5eMwn3srL9zPN+2Y38dJN8vvjjwUDusWh8UX24l
nzsUILHcYL+VRsibMmhmdjN9hdLPSCiyFSts0M/BEtV+ei/2zsAhgj6fSF0GSFanScuEblhst0S1
jH60uDPY58K6piUZ4gSkPNf26uI+q1Rpl5r7HcyGschGlrKwjYXKw80HAPzCTpmmkyNokmx5VjUF
bfS0cZDsQF7Wv401sHvoGGcmBOLBVcBzNTKZGR7q3rAtljtpriZGBtaZE010Nwwi5dWfoEVQHafI
XwPGe9iqLjDGB4MFNtI3MqPESJ0sOoFdgwB1M64lSNwnm5cWIPYF90uvxi7aojbNS/VdkGvxfOnJ
GcHsOUQTs+H7gsyQ4gL1r/8u9d8ZKUvh5Z6MRwzwox7oETYszRHvzDjMAc5gIv3ADTh/UkHgVPDF
bCgkMvkj/7zncVoBKYXvlPrOxU1bk8L5gMMOLflTF6GTHK9C2d889bHTCTIhOq6iPu400mOw/3Hz
OxXEUPK/eKtvuz2jEe3M8+e+feOOISSBQ88AtUijYmNv4UKLi7k2G1xtTSDS3BAPGjaxfGjI9q7D
Y73yLvWRCMP7945j2Xw79Kxqij12yC+OJQRemJ7x+LnTXyTzxfbDwcfWavdZVA+ILaEOS1YfbIrV
zrT7J1fLsuw8RAIZn54JruYcnxjr3ySOopjQbbczPs+mhF551rgbGj+MYwrQvPJks6YlPPUevddm
N3AzrH0Q/VryABGRoj/NGGtzmaSa6bDjgtahHo2PZ7U28ZvkvclozefRyYvfLnxyAhZm9YtGqfdt
bVN3t19W2cGe7B34rBoTdocB2oi6nMgPws9dK+RGgtIUFH0NwX6f2WFMFsKpAGumJENRj+ZFhE9p
U7TrMiGyh51Qh+RmMTTUd5/nzphdTM0/pyGjtWvRE4aW6RAt2s3Vzg8gZnh6iUsMMnzsVkeumoUu
xroR7ms17uPOlzn+ZSE2hpEjNqeQf+kTDgil0LABOpaV9if/2uJs9M0kDFjjGELSHpZBaxshUaiV
PT1x9rVua+DSYb67+9Y78wW6uDzzbVyn9s/YUBJHjTpcqMMpQPhZsnYvHxcUemywKVuj0GmSyODM
KkZuy0mOtFfIFehCkT2ZEd2resaa4vAMFqGRTTkXblWnx7VNpHGOVxywQh5MTjRTC/XakHrcNCF3
m0QrCRsniqd/BZ+GgaZpeHdySvC8EPUEwMTjGGNgbDZMbcyy7NmQUCexAoxeXG/8rMXAwSxqW/By
bORpf4hkakNXRFzBORbpjTGJhsyGw1b7kOmn9YIu2QpYi87E1IwlHoCHs4vJeQTyHAu+ksbhlENy
d7PW5xdu3es4/xX4AvPJ/KT5RUlzEnmWuU79lbV2JdrWtEnym1ZEnSd9nbv3vPFfdoDh+atPdBNT
/fFez6AzaxgbIl9+6EIzOV52gvg4211NPDS1kciTeQGHBIvkEMv4emzxaODf2G26lnoY/sNmbNKa
sHRFxayyox16Jtz5JVpcy5729FkrmJrHTpzHhoL51EIfukmprzjCF2lJnuZJELv1Vk8J887nGeE9
q2XMEEf2d4N2ReqOtSvaLqyAJyT7otVW7t+6w36vJZpBgcFd1fKT+gczbaJEGetPxS1ZTtqafXAY
BQA1051tHoMv6PoL6LxQo00ej02efvXMTB6SfJRa6FQ60o1uLrfYwigX/rRmtvHpqmu9DgPvd7Mr
y2FEsRKy9RxkiaNXiZiQJMVTtp6RJUAYO5qMqsauPo/+bO4SNlSy/4t0gJmYV02lKC+a9X4kJZND
ZXn0u0it0kSvtA1Ir95B1M6EdRYGd/ysd/rAVNAAq3uE8A+JwSNj6BNHNYaxMKqrudYVG3hO7iEW
cOL/B2JvTJyx3+KimiT0l5wC5Ry5TJh0Rm/aRkWkxUcc28DXEo3ToxfUiLMVUXN1hBHe75m2PWVl
DTe4OWYfiyalmDg3eADJbBToUztQonmdez06S4XuKpOpkFnfXS8odvPDQQcOPd8BpcnrQXyt8WhL
6faI7aS7hW2NQjYE1H7ZOdoPSTADrfdjEsPHxgkovreAyHi2f1X5hx5HNNJ8Bh+zhYqum8VZt7bD
3u4yTf2QwIo1ii8KIH5j9MLjA0p7BLgZjkZLVRyrRV7e3IULpOZWyU/VPJ2gcjp+eJvDmJwE/nnr
3JtigYtXQPZJac6SuQqSnM8gkSs+/a/NMWsjkdTi/H4keH17krBOUwY0haSG19yyD27i8qKlOOHb
DUIt4DUJA7QMWMopCkrEjRHY++gGCkzfMnMgnL05hClPXQfbGtAFwIE7stQew2HfokMTBLlgFhHT
PBdxMqElP9rNYr0alr9JaVhXsAXINBFYtojNeABwEfXbF2dbvFziM2wXN83YZX09VqZCk2BLYwe3
MeSjCrtazn9VV0O3r1OJp3wsbQ532WHTQCDO1eTejsbsxHFm3l1Kb+bl1qANePc7/olrSOfeRl1m
w8JjBrs3tbNzVLby2weKaQYkJgHM/Mrk6aTnsdWsj1cO1TLgL7lObd90TmcbNy5UnN8WbR+s8JLL
YG4wO1XMtmK7BLXzxf+2r43jV/e7feDqzfURn419kQgr+bb/ckuL5UcZSJKnU7pu+76MTTYSY2SF
+tTwK+xRymQ+l5l8BLF/2w9TCEgaLpbdcQu7WDX7iJxXkn9r6qDEPkHZCq5mdfyHxrsQHUBkwzye
+GiKRqocuVmVQKbATKHnf/rZaqWjCjySYYkGI0Rwg60Em6bfDD3c9d/n/WOtIF6u6vPaCLtkb/9s
HNAJEniBFf8rQiabC05VyPfrlvTDLy/9yvyzTetwlD3a3YLoBi+N9ET1T7CglKvZVobADl7pKkTF
42q0iinq9V4bGQfatK/Ywp7FHuQFnG/IgZ8I+9EkRtUlSSj6QCIiYXTTGmrV3bl3HsmVpqEaj0fL
75oQnnU1EvVI+Cnd3XXER5PlsQLKPNJ5rmCe0kqrOTuFPiYUyN+1JH6NuLOJPhsP7zRj5BSH1UVv
H4nLPFH0zLvM9v9/CicKbXBgV21FerXH9V6fbL1aASZP4G4wQGz/t8obzczSYi0WHfuNKKVCyMvM
MqTbn3cMV8UKxxyf/xCd38zxF92hy9aHMNxzbUqVbOWsfy9yZKGRfs2DiBehLJ6A9SGqnHdjeDFj
ptgKNHlX9vLhHPPxgnK4zHfKTcFv5RXER0klMahgI+dfocuGqiUd1tM62oHPRfU0LjaSEu1Ff8WT
7CxBPk3G+hRSaSzCQ5giMsoFG/t9YO1FNEVMLym+/hnwlL/VFBrhqdStGVah7pId5l9nEvLxiznr
HOePpqKaAmrESADbwwFAyVlDyKGDnvQb+wMyGv1zPsaK1h7t6K19JbXhSmJE4hYXn7sgAGvGN3UH
0Gtc06944t/KM1UvAw4QHqTXcsplttmDlrQ6gMPYXyn8YhBTcvvu/Y6lFPeLV0eaCWh09luhz0yN
HdAdv3O71sQmu3umH7YkpAllETKaGE/2VfUD750SANxmt7ffVautAJ3v9wVvDNmzH5MQYm+YrDXd
7BSykNaBorvn2p4Xh1JI8lPJnifSN3+8dpeof3RW0hgWB86n1iHfUfD4JtKU41f8Y43aZUhb0B/+
v6qYDjLYfiXlzByo1iL59jlW5TBTRO2+si9V8uj4ogQGmZxo98G4JUxhEfA1qtslVxZskVXaJmTB
9Yfs1XC+QhD6+qyM5lRQuOP/8svfZF91mQdQ0KjqTgd50iFypxiHuil/cIGZqrIs4UY/gAIHYXXu
8jRYQRKonqPCbzb+Y/uB3CwiQMmQwxXjQ+GZCyxzMEAeaKO3u0dN7GQUSSekygg0xiiqkY8intnZ
CaizLfPwJqod4YNNXTfxR5VPAHxASwBvzbkBujm+5Gok+V3sKosfQcQewBA17QJB/40ybHNyMVBg
h01kmjuvc0SvrWglVR52SOa2ZmvXjTmt65rtad3vCzyji4TmWa4D5f/72FA6DmUzdFt6fQCmLkRq
FDAqicGBBIXgY1jkgyRfQhGYFjP/4Q7s+ooSAUynMVzxQkTZ/l54oCTa9fDBOEmvStdqMSPBJnti
mpCZ4pNKvvauBDOZEt9iN2bFPq/DvuypYY4FPC8LgcFkEONqXf9/qcfs/W04ziOEVkAoSuXpJiFL
NtB1hOWaGcEGEad94uSm+2O07nSqfKvUNW7T8gbvithKgcfOpkNfgtxuNl0v1XadaihpKw9PmfOI
3/xkErMAitCUWqCRbHs0yF2lplMmkSCN+rp3xnLTo5oWEo65O9ijxPqaIKynXd5Rx7+BejbI+ATK
pVnAfXLXnXFi1LS/RoEkNo49YNBLwR57vK4ol69aj+rMj7Qzqb6RlxS8oHu+BWguRsK99ZdriRki
2S0y4Rl723J5Ey2zSRYe4hvUppBvTuBb+gX+TW0P2yayHneR1RTlJpEwdzWkv9qHyDKbvI4eq3Xo
MQDH8hyvH/UNmzNENNtcTanBMShMtUrs2UgallJgA1h+oP5D0XAANUDJgP7t8tHwX2+9D15UMtUr
VGjuA39tQpIpxhRDVqBBTuOuuWoSGSodrtdNyR9nMXhmAgRFHkRwAw9Keq0Hbqnn2NwKKF0TXaW9
fLxeULhB4SrzWDeXCY0F/QxPymK2MjczPEANCPQMQXicfWREf9IqhVdvYlgUaJsQ30PBuIKlxAxe
F23Qm5HpzkWcO0EACoUVlTAjfLN8GuO70pHhnVT5Z2gTN+HMiwm892BvUG4eriDomQl2lPSO3nJX
opcWD71xKAQJmoQk+ADPJHph180U3IhOoG8iJx40L9EdMTzKjzJ2mMJ3kTgjjI2rJLIKvCP6eP0u
hu9/c+vWN4MOEZWal7znx9DpdT8bOUjKNoSAQ0mATJba0NuGOqYnOxzy3YfbfycGYx+HEzZ3rKgQ
yihewEwPmNUqrIMNdMcsoONdAWH4S7FM+pxkhxUMCBaLW0UKUSKpdugBmBczTaGx4it9XYRk/v/W
yxqnBQNWHYd6FX9kKsg/vmLXvbGESRwIFFbCULI8vaNCVbRczKxer6kn6OMMaWJjNj0VSBu/XDYh
LcmCxYDp1tWD7CUdU9SwT94DekZVc7VTynW0DByZB4hiTRngsru6SgPGmFLABd4i3wsLfX+kEgPN
AIM1l/Jv/xwiuorL/cwM6kvQESRM6RcEndhKYQToXU7zYIHB3YkFQ8asVjZff5Mlcuo1R/CQfrln
sqLPPiv9ygPog7jusy/AfoKK/d1foz/aoAEEvnoXmisSWzY+h11P0444yt/3inTIsxB5qY1Vg6sC
YRy6pYfXouajYCkPXRuq/J18RVBCqz1DbYFvByZl/OHgrrpGpkZIf3keozzLOsO7vMpI7AJgRl50
k1nnbrSRqVPdEH67FvT2MfELbSxGJ0+qHuH23M+OVvFkZXqRtwcBm3ijDYM3Ox9GozxAwKDTpHun
obxNFo9BypHMRn2wtC5/yrl82M/nQSLCoDBYRxSz1sagLOyw35ypMy8+VKtq3j4oHH20QfXsXRmK
tkY/ZX6Cz5HOrUoPURBJCW6Tg3FznLLcm8gTtREMX2s4nuKmTK9+AZqF/UBEwr2O0cAgVAZBQmH9
3gsBtnk7eNzlEvbE5oUBABPygZvzH5+K4Zxi26sMYPh/9jzcenISuU2LWKGhcsqovy1Q1FynbyKC
4HsNzc/h1u1lkv3MPwdWV4ZWt0JmbDSo+yX77nK/o60aYe4pJsN+WLGO9y21LXT74doLETiegeHv
GUNRtg8aFP+LiF7ZrQH1+vlV7THLU/C5m0wORBiXTBe5quX+EQiK6UXJETqZgETec9RzIWK4E7YR
rZapYbjEv4Be4pRAWN+U9Yv+Tp3nPiFG7wmv2Axx5rbd75uE4qMDuytGNUbP7a6qcgb1bFuSvQlF
JrKlYiDFYnM0NCj8qHmg9idDuCNhlcTTJAJAvdKcV6C3kTOew6fNABcEXuNvPIGJ6vlB4cUoCN5t
PRK7pUSdxyBb6tbr1UGIhdK0tjZVkHbCAMPv1vEuqb1HBK1vNvpHlDcGa1TFUsHqhh+wme23NZ0x
rnRjUYvqfl5orCFXVB6+fMj7mzzQsx58mG7gsA3DvfyRzbK2uhQtg5r64voVVTsmgudVJ5d7rlU2
vnOTfxul/RZPTnk9ZjTMaPAFvdtrjCYwuk6m9x50VQv3xscEsWbnAvIFnmtLEc2F6U+bRbM3Avcd
YZjQJX3kmKE9kTQ7W7pSgcu68yk0ONKyjihGVWCk1LZwLU4/Pg5lgkEri+tompigyVRZEW5C1ftc
EiUbsKfpGE5t/qUbxN0Om1MVyvqKP4mn6UuRncPM7bSpmYmOS2tHs2FCWC0oRwJLUCjbaPG8LDZc
p0Ti14b1/eJODlnUm5K2dgzmc0V06WKnMgoJfNJ+Q6yQWpWc2mHnKrAoObc1mxM2RPSdrAtBgbBY
aDPVaVixCXaki8l+JvShZxqNylBzPETzt4R8qFBUuCotWrMYO3L1HuVRdzcukTV0lWfCP1GOXuBD
1dU3I4oRd6jui21Ldw2Xgi+u8w+i3/T7kIyiBX+jKxP7pc94/nHEx3DTZYKE1m1ClP3ZdzAUVgrF
Xqvbfp3Dla2YETWCo79+nCUuHovc6Xt1JQslusX7vHWWXayft1GnVdor9bWgEBljkaSd4InHKEin
IvoP8cpfsY8i0vtR9eCoYsRqY0TF5N9Nyh3FwWFXfAKo+8TXKBYXkR82PEZhNTXZ2RU+xPLo40ak
NWbLPMUWH+BO8W5yRklrYZBcIVlzQJeyXs5Y4O3b3RsnDpVT6Gd+8WfsNaGr4hkq72Ad7gcresRd
UpGiTbLWClqXyTheevBZ9KYPCPjs70syiBkvRG5ehEkDtijCy3ugm/uMBcsXZfENSRRDA4Klj2tC
QD+dd3KLQG5OeB2lWmgrpX79Dw7FZppdMOtSTyaAWTLYgu32Pl3160JiyJ1KGVFchqHRpvLSfy9s
XQtvzGg8ZMfggk2It2WDwGD+f43LL7IV1WLVP2hafsBQN52Hv+FOLfeXbAX/v9iBJFLLKZJzitRd
2vMenMDysBKdB0zbK7CZP2KdS9bCE0DWxEtnsbGj5mkGLS8+mRDkHpHyU29hY1SjUNa8z0hDyAVy
80s8uMLI13VoUK+8J0e8tA4GQvi/svCIp3YDaHe/51FyKikam62FRH/egl3pL7zqQ50HB7QB4Vqm
QCUpSYJ76OP8nG6kZU3R9pEsHGUHqT8AoRBz2FDuw9txusQpKuNPRdMkMEDj+XcS9d3HW15H0KJG
JxaqMk1uzjLYhFedznMdsuWMZNeSnluNbPHoJ2rYEmBN9H9zf0egOTlQuBsw4ZoSe6mUkci1SQlI
Wokn86bzasnHDEAU4P8HoJwQluIT5WI5Q4W8twqfNgC+VPmoWbRRkgbIt+8TaXIs3BTABKIod7FJ
HDXJI4286Cjwlv4rerXmNHKyPvJscqL4dZY0qrqkRo39RvYjFQ37XvYGAF4U3qW4tEGTaRl9Cg0j
g0u9/zGn+o21ZkIXelgiivw7Vem4aKR9ZvD36vX2Sg4c7KyalPToxg4WwWVvEjSIoN5BM0Tib2ro
LsUvBl8jcztC283XKCdwlBvL6zB5MoVAO7QFwgyV8THYFJnBVUxpGhTXNWODRcrWnAbvqSH345t6
BpT7hipSgVlSwEEBzL596r5HwOAOZDD1QAOc/iVVt2WSufCwN3N0+5P+UzanOzYX4B0LOC9Frsbx
jLH3IlPvfoAuSLSfX0d/6AHLfS+FzyqClLjVX6qKn1iwsJcWEwMFUazITqexfiogFJAqy6PV9Yn9
aesDCTqj0OYSj87SVLZY3I3JzwCSBbxAzODHLxjEs9v07n0BSWPJKTu8wCBIGCt9ZC5/6O06q5Pm
dbf72Djua2UGxXAIjqGEsf5GvZ64y1H61APihtMDt9bI8GzWIOPsjfq5wVg1L42Snq9HW9YI5XYW
Sk++loveDQfdrR78gGSY2nt78gWssbY+RsOqBaH6XX2PXeM/WYivtD5QF28EAAZ94hCbHCg+ABAV
rnJG07tlEl5C8LrRtgp/vPsZ+sAvplEnFIJawSXKMpnlN5G0xVNbJnhjFTYfJU4I42e7sgTUqOkO
v3rh52NFqmmhlTpJ1uFyhmKMZj3C5hGJJ3o/ziUZma2c+zZUCyow59ncjHPmV4c8614QTgE2QRzw
/gioOkV785ZAa2dEtl4XfNZG1IVk457IHuzDn5yBnwEyyoRIDl8hGArICHxaxupYKLeBJjcDxR5+
Y/PrT7DvMZw9o4wk+U6sdmQMLhrpI9OXfLWXnC/D54019PyM++BbVZb2beFBMBi5sPtAnF9FqaGz
hkQtluORVww/typNpYV4xpHqTdZkfZOS7c7uc8WnBYxQKtfZiyg8ZfWhGoUTvUX6a/VGELAVDCGN
F1kGGu10G2wL55TnQHODpGzbi9r8lFTwCact5FOjQxIwFcUJbLmN6X2SWjfym4yIwh5JpawJ27Me
bB/IhlVpcxNHgtWWtOOoxyPzPQEyCng4ZWqmFS4X0aPEVjS92IyIZuUFW1DoG+9QqvkNRRepp82j
Sf/lK2QQwotXGEr2kMR6qfEhgCswuYDavZa1BmYqA/+y5sj8/AEdPzBHaH81Qo1u+NgOcAhGb9td
FI9bLQW0RBrADFgF+N84Wtd7swa/N/578c2p2qerIrkzCjF6vuN02v2zx39ZzqnNlcT596nq7oxW
YAlp25JYUvyPe3JVaTWQyqCld/KtTJFgc+H9YvwzvWyLR/4qqN+GdsDBNbyFzzYiVdaDQDQDK7zl
0x3Q+FR1Hav306idHIdKVlaYXnNmr5cWubWxtk/25T+ex/4QEaCzZ/Cgt57KftEFAILP0PX/PH5o
bPgeW6CET/0naWHyVyenfGL5IaVHK573bbYClnuGwnFTX4Xf7ejOOspTzpsuqOxibmEuqV342LFl
CuKQuel1e0lCf4j0azweOG9mDRq7P177ezMFxfOKQ0L95wEt8X863rdMKdm99gBrfcnht1nvSqfL
yAFvjw2P9ExDXblLtRDeOphQkzfKslvgRY38GxbQU5nKeIbHcMMH1OHwQ5hiGVWbAR5dSpheSOS8
tneDUx+fy31wMzodBUgGrQwgZtX4DKiqk0pCe2fqRkpdPQYCEJfMit+RPteZ/b1B1TSBFwLnapY4
oiDxQVfL7YELFiOZ41Rjtbeqsi2LwOPJ2hrVNAOjYTALyphf9cS8y+QoAhiJwMQQIekwMkI2gbdd
oMRDHlIGRvC1Z02B+4T53/oqR43L/4YzziW/CWcN8ySMJtfKxFlI8kkVDx8ml2qiluiGkhByWF6/
AzwvW0gY0jz17RcC2QcqbMps35nJOBOSCAgNLZbBidtZm+QovMnWWIoGgRkx6tNTWT5AAEx87Juj
8YGaU9XDu4MNWhNKV3jB/32dKafeSHKrYH+QF2GuZJJQjcNmIoJqnISfl7Mnj2+Ls8mryW28wgcv
4SA0iYrrUFK7PZeWs8zQSC6sxRjSUzjU48zks4ccVCmvjgKSZ//lE9FTZoBayIqn/LeZu45eHI5V
RYtCJPDI8aHusV8TFeWPIH24uGI/wtwzRST+xzhY8wbIdcEyDz0qsWraTif0Bztpj12efMwA0HBy
aXkRCMqCKM716jBMSXEF/MqgcGOfI99dgUAHlHdNuT2qH0MSzAu6gn/1/mHbKaZFklfEnRxqjPr7
3l9Eag2StLf5nNvKDWd0vMbvMTt8poNoOWaL6TMpncKFIqMbUbrFKCxSd37M+Te4NlkB0wQAqV65
WZy0peTiHb/9mOJMY8LcB6nEyKYYMqSQpo7v1jyq+xSZ10HI8cz8FkR8WVHeGTU5VHz1nwuVUxkh
rEi9/zFE50iV1VWPvgzO7WnEoRpkdGGfnmy/BfIsKNwp9yvZRd4OMky9HRBTdmAYe6i/GQvt8vbJ
wg1aZsY519bVPCQpL4F1OrXv53yJ0TlHNx6HDt9/D+sXOVc412ii7jDzWr004pfLpH3bFOyTPxc6
qLvX0rkjXuxMsIgnGpBRQ0ABIYvesogIwz1intaf00UUoyfpZ+OFNH+GxeUMghXXHAjdioowB9Uf
bvGFaNmYgT0GlbZl8ALB7vnLwRhZQmPmkUCGWv4yPmqix17zIz9aVMfsjShag0DQjyQhh7/EqzPV
H4deVyOjRRCgGLBjUIgFMXEc2Tu/dAJMaS3a5SmWi9A4gdFSn8fUOvXrRAunNNV7fkbD5XWaOfYh
GKIpd4RVcotxed2wBx9bnBt3ZzrIa2TMvWk6pGlTUHjn4peZAWsO6Y9W9B5Qr1wRcZhsyaQ1GIva
eyU6+AkLwoZL+tG+JFURspBxzSOgSNuzVsohTVGVzE1X2LEAr1MLSTnLfptviIovHcbB4750ZDzJ
dP45DRbrrOhMztIvNZAqnFEIuMHexlhBRbWXyMolbYiOKFiRqXc1FKTudeSlSQ7yTsyN1pOH7Uau
sS8dSBj+jTdtsHXw01tsC/3hc+GDCQcoE+cR2Gm4d0NU4lhf7tV+pRGMCv2X+zKkLxbrv/iNTyF3
zRVeefO6YudVKU4vLcnkjRC1qeGA5GmwMEDseVOXGd2epcDojRD5dPaJXHteMSifl5trXdpUKJxt
Gu+lDNWE0MQV1ZTecKXPyaAQR9BJyRW3+58l6pwax8usfyGnwNwJ7wIRJv9+GQOWaP7LbXAWT67t
3QiJlCqTRpw8HlVArRPq9kMBIklc6gQo4Tcg0X0zhVpq5OovMaGY5wUB+n0i0hga/fAFUCUHm+AG
dNf3d8kTixOG89oKKO1x4CI2aYw5UDiXNcf1lsDW8bhfgYixJ5O+Q6LjfXGgKLs9v0wJi8UuTGvv
IUYJvG6mkR/9oQ9hP8rQtqVJ29GIea4cy7Zbfhf9MYG9JicPxlHABkDDO+1O2ikCiqkvaYr5whhY
fHvv0XlnDW9bNWbKUUGg3H1eH5+2UfSUTpy1CxlSWEetcBufK6GsXe5ZbcxuadFrQkmGAxxN6iLD
JCBGf9ioVJIW3d85+8053a/D5gHUuIaCBCu/rLkUouQCITTwrg744GkF4jgVZUBEmP30wUp4scs7
UuwwKa+VzuidithdcYS3ekqy9rTVRBWcPPYudnAWT3ewkRQI4F+SlXScEtR1t5pMGEMI74TS5D4p
vPbMOseGoNqpEdnXBYo0oRCiD6Vg0MnYN/SUuJQkfOGJ23n32MbvtqIr/UqfJGiGZ3Wr1nJFwEeZ
/D3m6ThrmyyAHmQxgTtcl2IL81ifIMMx4w0ZIMQyTygZnFvQEpgtg47E4849iYS9wlxkj6NHbDyJ
uGD6fAyps327pqmddWIS6lq/Lcw+UyHVIadWhAyvF2Ua018Fk3RroO+zaTXcDBd40NlLGegdYAlR
iFwtw0V8qejsfFAI+xI9UxEeqohXJ1uB/oOPwYKAfQvc9Jbw2GGeiooF5/7UjMkINAYWkCymwRhV
Pp49I26gk9SuBWcKVW+ejy2wq25XW3cqTSa/umFnoi4OSPbcUkSgKtXDwCJlv+HGkJXevxo82/10
wEgQ9YEtEjP7GVpBDi98IYuFPGT0OZw1TJMM80FG5vJiGN77cmT3T8i6o+IRnbHKCYxiOMBCtzHC
IfDlMn8eyZcsrG0W6TuOnvOTMdRBxWDwt6piN0olZaPiiYPhxzH2jSQYpDeVBPDWhWwGgjPA6Nnx
5bX/MG7nAcLC1xEQc+EBq62Fhdn34mN0RBBnWrF6/MBVgloA/uIuWIZy6qEk6zsIbA+Ez6lCE3eJ
eqsIA4Ao01s35Y99Aidxg8twYmLfmBuXQl+/sfgFHcXZ7SKUIKEzOVV2iNL6KreShZwv6fMgXvJu
3zwDvK/1GEZ6MfVD0FxSvELkB31jVpn6Gqr4qbfWH4RhqO4F8nHDPlWMHvbgA9s1JKRKtnXtdKmg
JZR9YoB3i+TZdR2K+U3FNAPAK41zTlqy125QnfkKtGl2zgCkJ4KPi3dbFZg0LkPNxBWoZkNbrH9s
xNVhj61CTHZSTt1rbY7w9y8BqlTcdTWqUuKcEKem51UX8OBWy9WD/TwpKWnBlEtt8Xg46MhLKEuF
TmtYVZd7odc/dfRlgp0OAlUtUQNAFsofPUt4L3Fx7tj29LWUWgCRm5n1694wO2Fhp0SeOHxvwMS2
6PMau0ycUnm8fVshhHISTUqFktInoDJXOKWUDdSAY3/lpEeh1vyjvjKPl7daNC4BP5Q9gD5QV/RK
jfVob4TpdKLb8dC1dULeXjezmQ04PiiuHWY1/wMJdCT0FiTvn2jda8so9ksMB3q48VZgHrwHInZL
wbSJA4o8e50YzEChwjEY9WIMGDJJO5qkgONMaUumDm8TwZZksJOY3FZgMT9DPy1D8GFTU+44hTn1
xmtfTkEZasqiwU/YBPqkiwdCTgpwNa+0f/Rzg5VlTaedE7KUQsKtGgX2TBqT41wgC5djXVyRp/7r
BYJva2XaGLfNlzsfWjhcCCv3NWJ3sNPJMLVjt74YQv1P63AI86Feppy1iUWF/ddO5cKeqseH3hxL
NKs46vACc1b+2XmBFQAVAplOtzw8qGl8s4ns2szG1QYFR8aHD/G9a0O6wYonkxowLpgWUE+GeWVw
wWlSABfNRHQuJ69ejuVQRMQ80zU6TgVcf07SUvYNt30AmF2CDdZ4tDK2jtV4t3aPVMk9nqkTT4b5
4Pdu5JHTPXVPVeNb37n/PhLCPNIDq0bPn95e4zNURaSdz+kw1QdDnD1oXwZBeEX5kZscwJ662Bpt
CUU+umZVDJcxSLtAgIV9AWN2JILt9egkp03x3dPsx519JUdwzy5aDiOcYtBRc9vEvl8vEdCj5kUE
Onv55+vFUDPevRuZ7mMW9f61hfza3mingcbre2fX4EUGZ3t0+U3gCzV26mGsUsyUAN+KQOGxE0X1
xvVTN9YuYkQG90kPHl/jdbmBX+7L8M4GOzSM35GCztMdAFs0rbitL5slqKZxe4wZwoT52fO11zFh
w5ijOFPztHknqQnv/E8nOv7PCApph59RJXqrMlIb/8kS1aI7pghvtsglo2EmynTsS8QjydTaqw6+
Hrhc7axaVU/zDzPqwDjD0rTkUPUkXQFxOtAv68iPvPj4pWo16NMa1psyYyRXxqTfc+B2bubrezog
oahB7dKIU7AcGXS5F6VfI720Wg6ZHcMiSfKcMasA9vsqFcbNnTUO+ZMDBgIqLbu+PHq67/HtJ6ym
ezQ06hfrKWcj3QO9+RJM5j4pQ+5+wJC//lZSuW2DPhsxTFA2ccdjxi1xKkRtPLVBjoB2tgiLCJ01
aasVyZDXQ2p4EPpGO0ytNAw1rZ2wOWAspa5aMzaUfvocU/7bISENjAsR11YCoQdQhRsM8xe7sand
bRctvArqX1y0VW+myXLki5/Lp8aN6m79Lb8aD0GI21jJDT/wpBNZTgbFRHJdDYEaWogwyDCg27q3
5xqLMQA5Q71Wvga+N6raE8kRUZk/aDf2BHXIRiaX11XmA07WGMx73QlMJB/n/DewGCgsiR6DJKzx
3lwNJYzi4dGEPwW1a0+2puRa51zv8pRA+G9Yo8sZpdsCGJgtQ8ALTxH1DMXAjuJ3ab4ZY9Utf/4V
VPAW8+n9C8W/rXnyGycABM5qOjQDfv+dX+h1lEGX5dhVgmFmJyeA4FhP8iP3n1eSjSA51NgCOtph
2HnZBO5XzOTPjxTf9DufU7erg/8jGE1rFnsTZOZDkk1Sah2iyQOrALkZzxwgIjEEVJLZMsatz5Ui
QWNk/UFz9LHCC1iPk4EdqGLiGd+z6L0fnANiiGCbCA//x48ZkwGXSjX/lxDUhCGRZbiORU9aUoPn
gJNczB89yRvmlzMMPe8PB5CsMeVJardJ/fCeaxHI4CQDxG6nE4UiDl0Xs2arLWQIqRVHnAxv50tl
z5o0WyOp8EwqxdUUjPtQxh5P62r2ETy+dxmmea6rxoOLKbjKw+DTmyaJvr7n7kuv1JhkduT3rsFp
X+cZfXHihVL7r4ANvMtHpFNpdZ1tQStGWWcGwnXyMRoM6oBDoRQcVi2Gsi9IDJEOXo5lW4nSMXSP
SETfoBxlJ5Sy+pQCa54WB25KkCXAUlPe9H1ZzY3CPuOTDlv/Xj5Nx4nV3xy9sGipUt2wxGmPXSw2
QpOUpIBBfLuI8zFatuPBCokNbuwbvOLPx7CtEXNRK93pCBBDvyV+sUG6DAEF4FgC8ElNKKCvEF2H
gIuodbt2IHEw7NbOsTllncPN0usQZUcXEYPLd0I2dx6NKEN7mafQp33sHyQeM1t9W5zDoNGOdgVt
6ajQFPLtBxcWxMXYE839t82SLtcFLnob7RSAWQoBGlNOLsh7MO28kCi13RamQEbSojQRqREi2Y0I
vusJyExphsywneviRdMEGGMEsKBjVaxHjXFQ7NiqjD1ITfy+azG/m42kZtl0Igz0Xrtw0dUaTWoq
XPqEFFzRv4a7JWYzk0oj2V9UtAcuciEx4UCITBxcGxadw2T1JSCzr0tLEpBvWIO+d5FK8m7GRtkZ
Gbmw7PsuqJt4B8bJ7yVY6rYJSJGImu0ebgO3xRQ3bEz4chbPoUbLVm+h5zv1j0jS/DuUk2+ijW/K
shWV2aQbF/DgXoRrtEofEzijgkVgiT1VE77XYtbh9pK4piRlUWkIpXnP3dhjoCNa0eWsIgCwygmO
gY5f9zyzEBuE2pRfrXQfXnEFiItUt4ENQNAue0guNyXVabFWOevPk5p91/VY4y8ZT6XjgHPoFwBG
9Jk1hMUEsGxl51bZQbyDuqtHL53ACtcdvaMaThsSLjSUPFSJKqf5zYyV1DuTJ5dg1ka2jahDyjPp
LaKyMocE9YPYY1mj5pUI0Q+WaI+mZ7ZPr16LtKZx7EQCYlIzLSdMjcqMAcd/IuzgoKhkl51jJzxc
J6GNFUB6SQR4XrnFtF5YGZoUV/vEl8brfD6R7veU/qE4umducriedd3OlmjicwMJWsKRTOY+5r4G
2HSVjT58sSMlSuM2s98i4Dty+CtAveKOXObFfmhnUx2KxhlZaXyZE2PL0iuOMlgHLcQfp8PYWAuG
TP6QARUahamGnLqWMDPatlSAlMeim0+K0SgjX3xmzrCmaqcXB5FHQZGcIaiQuVT/DYbZkkJ4QiLQ
3Bi7J+eAqzWopHAeETO3iXY2D7aHoSuZN4VuaVjJqaUEVXE36XxIRjhAPEF2EIkjNo3DdAmlyHqx
ob4BmAJtdJpX4hjvhbv6nF6uBQMoxjXUicKOmqsVoeRgWhauO3au4p8edZxGa91cYsryV2WFtLLV
KRdt7xBOcUS6hKezJo2h7iSFmZnrZzy/Wq+5k98+8HL+9Q2EasxTH+MD63rsEwrInDp3eLJwhReP
DiIbRErCboiFvK3VbqWZwIXQnlJJeAzLunq4ideyM8tM7LJ+gzFBSfWB4w4arHOOdjPe1aYoPnKe
bhxApLg4XoN1zb4ZLB2SSrrbQ5pixRwW6BEGDOjX5KUfruyGP8K4S/zj2ieUlRysNda8U0RYRllq
q9JwvF1LzMAkQeTE3654vfsnC8KJqnRrhuXKMTQlam6mV3Wxns+R/rjmB+SstyBCBUlr5HbqUiO6
QmZsDBsEYe5d6J+3iPnbU8QEnl1/pnQjUyns/dMdqwYBp8q9SJCJxzaQi5QA3DEVBwMwCLgaMPBz
COiSafC4WsrFYfuND1I4X8d3o24X8QdpLAjn21Cn+69HXpMoIo7JoSYIn2vlBqH6N9LuiLhK/QpB
CrjrH09EXKdnuWkyJ6aQ1SOSnrWI/HaS3DzZ/F1cuDaH5abCt8qojNN6bHFGsLrJtJol/ASEw1Rc
KK7rH9oeRbIKCyBc6JXPQd+r/3m4e8wgDFdC6nYDGXi/tkSqEKJ/X3ATzQqNjAiOpQzXMxajnY97
07q5M1mJXqxOtzTBZOmaPHaRsDh+amFLJsUI+VANuu6fbKf53UTGx1JSsmxVWSrPzzdky/eR3NZj
5bd3fTdnPVAu/eBWnF56rHI6pbgnmV6NhpMH7PrJOs+EMRLJKPguoXN2hhcmfPTQQo4T+ZQbf0/a
u66QtUyRItBHHZekH+/HxvOBRPkaZRBPkTwBEkKGF64YRjXe8A+ucPoNmFOU/AI4AaUNECzJc4j1
6nzUcGex4+WfCN6qPB5+rhdIScxOCZKQcUdDJ7DNabtYV61AWkObh5k8Jcmu5RXOMrlP9vYaSn4c
BZEecSiZ6YeP/FfiX2ZRrc7T+/0hllrlnuJXYyJgxaBYpd8P3FHUnJjm4dqqb1Y2FmaKy9j1NEya
o7cvqu6tEADx1bjvs+1bvLxiycxtGL40a4gpVLz9/3miCI/109KdRhhMptvgyJjMcqzN6hSdtKNn
sEMOHpsWsgOuk5cyck80Ja630+VxmYP7IF24uBIPKmRNM59vNt7FEBfI1Kv6vX6gxIgiePvWlj0M
p1aiPY0Bm9w86fypXSYu12QWEnPaLpIyCtm3kjO7R6Gq+1pEc4K/+OnUKmIAYk2kaH9aL2mArQU8
vt/sY865scGjKPAqz2VSkrLGKjHEFLrZ0uYFAt73/sdXIsdX3GU0g5B9Nd/GgGJsXOV+iAqZCLmp
qVs+9UswLwCjpXKdRfJPm2CZeLHO3ACC+6rKfwYP8kS34dxUUUMyC2+ksoMoFBR3jj2z1b0DLA6I
vyxXgXTlNSNloabT9zV31ywbeZqdVLEaCqcHqzMGdede8MXfHMbTnKUuhV2AcI0Pe8DV75k8+tUn
jGMKTZ3mGC/Ar6fAGpWRFFHuVmFaRcTrFiuJdFuSX5CAIMqI39iPKFkhF718pax8xEW56UnifViB
X1OP7whshyPI5X140r25+vYaqJGKCh0V9zI95gXzdTwv0nj/I34MbVJaaIR6XpPQbb4ub6P6m+/j
B8BUss07deYRKwbtc17nn4PHSCj3k5wj6hLe7d4IkXTuPblf44sNzm8AgQcqQnzLYi4Nm6qOZZy0
uUFyC730/8WamxBlU0k8x4Pq1cAVEb4qKaHytZ+diJ47CWPrOEKL1dmuQ05JadgO9nUB5fUXRFN5
r6WhEHhuseMCM3W67t5l+T6i/nTNww3gRS9vTjy6f5QLBDairgrM+c64FA+ekFhOEf4saOr83S/R
PuYK2Fjz/XOyskDnGM/0NhtG9Rul0Qav09DWyMwzaYsSOecACOwv0JSWn4I9KUwzKadNWOAYuMlk
A6C8cJi8WfyBlw8XPLthvj/pYFH735rM4Qj77ChvX2CoVyUxSb7mnbqLgv/c4G2E1RVIuvV2sd6k
1rw405m/64ywBC07r0Cn7cP+jF6TxVZtKIV/1J0wJHNsP0c0R85t6H7SRMkUccjtJvK0HzviDA9E
RoJ32DZcX0J/7/8dr+ltmrFTOyB4gZxRUIzJRfB2+ggR12NZy9jNW3XicA3Oz3EY+gtWr977zxDD
JElNXU+a9kb2kKoTCpkdmfAQVhvXoXRq/s/YhciFle0yyYk4wcPb0pe54a8okqJ5272YJCTIiFGH
mhzhDbD9+MrLLERnZ2j2qX4Fik729e9j0VETLPGyqEXosUI7XL+X5FHvqW+xpb6DekPDJGmzWsz7
Jpq5uq8NUQcSN6xW7Ayi4BUiiLYyH6Oo3ctYGmXk9wWTfMOKEMbonZ8VKG9H6oIOmo/Z9M3oNWIp
haNYjGyjAfB66RQ8tyyVbzErCq9DoZkl/9sCtwzjg9MIZNK5cZ4HdEpcIwS3/ZkbHzXQH4cRdKNA
3YzXKPg05Dl8I9rfp6SUciT3Fbd2DOP/SqlfeqtVmDpsW7ibWIK3lNMska5OX2/ZAzeqht/TOHsh
P2ZLwDruEXZg/L6YZCCKJDY5JoKS89TJ3OtaJvAojJlaXbvFVfgp17VN2DvfbJSjTDGOZPBcxQ7e
MupB3WZGxwl3rgW/+zo98dY2MHW9HQ0T86R77XnuTtEIL7SwU0ykr92EbfiVKQilDL31MdTh8gvU
CG+6Y4hMChzZycuWBxQkUchUiE6Etm+bzRjlIiqvjmIhlQ90m+lOfhUkEhMcRyCrjic/Fbg5j7gw
h55pNlNDUnDDuG2lyFnuDFRU0xqJuksPg4Uywy58x9Ss7FMQoPFwb1eRiw+AkHYRzL/me1mRbQOi
OcmVUZ83lKyowVBVc7gW1fnKjPJwSoscm75pZfp2AyuQhgrZTyT3fftPZC69rsN2s4lDaZn610xs
NruDw9i4VwkhCy1k2ZrrB9CFYrN5oxm8Fk1da4OaEYQt9MmbLWlOWoFp4gA4KKDuUi5ChXIT0QI9
FBLIcOrnDFNF5RBg5W2itB3YXRr59dEz1emQzwoELZ3qK9c1S7IigaVpqm1iZBWVpZ/Q8chAokWb
pw1vFssbpKxtUadjIQtT9Qr2aPEh2rDCVsCy8kSgdL4gWOp8hf8+AH7/9D0AhYMV+D0FNzj6O7Y0
wnGKdY1Mx816sbhWUZIHErZqja5E5SGX3JwGABH0jWSeH/cWneEUzhn0+MQcZWFIUArfeNayH7ug
OBhsTNiADWXCy1tXvtqwUKbnWzOa0DCWCGew7umyzLZAFTn0KMDG/LM1lJDWQmm786Y3YFh92rlS
qXUYMed5pMKYeSELxTHX6OlmlliByOZjz0/YQ3f8JGI1Cfd9CZDxXloDnL1bVb2rdoa2s3/VsLn4
aTXT1NOkBClqw4WLrERdD27CwCWyVI6LAqjjRrAmV76I9CbO+Aacvn5X0yUn42CXMYMA75X7n0tx
rWszXkKHpJG6tfiFiD/v4gtoqNWiuy0vzElDyEYJZxpiDypM1FEsg5af4EzqCv40U8VfoILjzJWl
F+jOkr61y3nQ3IpPG48+CsPByggoiOJ2g4/IRFxhlFdJxjqlUjzqRD9brMMzvK73cdZmSPycj7bN
qHf+VvpDlKxjOI0hnTKFM714FCDC+kbt022ViVzn3hyvS6o2YPSZauWjBvU0HmivFi3gJGw81dCE
wjgcxoXNRvGNQRIe8srHLBCT2xqvTWSrV/REwIUEhNmd2vb2L5TscNYwmS2elis6ekT+eV7epiM2
siric+n4k42tWgQAkUzP8gnSg6a/eTPTKeMntkZ7noWrviEumgPAeE+d07atrD/wHOwPhsAzo4La
hpG8/ZysXP7m0Y9EK3gFGB/Yizu1eEpsxaPt/l66XxJh/cfBcOJm5yopCShPorjr9BQu6wmfF7f8
ZnNb8LOBkMJsW4hIIhXWxAo4rXrZapA3GJtxvCfIi1Sw18rMBQLzY3eWL18kbHK7sC0uA1BLPPWm
8BXG7mg/DwPEz9lxoo4RuiX7mxynZPe6pKZ5COJGciKdCtDkzOiNeKokhFrL33rJNCQnq6apEV/B
Fr72ZmmMuMaQgwakoxZtbiCR0WN9gzkAwePskYwQqtmttDshIZuvkSXFwSFT8iJ+JIe5B8aDtUok
WEr7PkT1hMuZarzohLP8enBgTAnHLFXcR6dTxEIU/sIPPly2veJJoVokj16fV2j3ea61hiVnP1sS
miw37EmZw/UNBhghf3gE2QFrdQQlte1GwsNia7OZRZuD5r5EFTwVLo8dkT2c88Mpz6MUi06ugeyp
wqClennb99un9ypEAtFWNm9zjEokwyFi8NdzVKksL8X7zuYMWS2AmZP8L8IUhuTEVebnmK0Cxksh
2EHNaoCGnnTLSLawesYSC5YM5w7FQJBN7oMKWtZPpMRA5RycPOESyT4U+0yxJ/jOARt47Q2NgdfE
SBoZV745MoHMGLrP6bbbzHHskB3IO/S5PsOzvIogcC0xujtTZ5ymPlI7RyPntNMsMBrXeBXM0YDQ
N5sMiqeRTGVxiRbSND1mLK2a9DVgDuldVf574NgjyOGIsNlJxYrLdT60qdQ1pjxrjxaEnk+MUUKI
/XnkawioFIzL4FWQVpRfud6a3jx2m/pIgBbxlQ/jNTqG35TB0Th0GU3AxlcDJ2xxBrZGkHjwrczt
Ee46FP//DMPMN+/bGkTn5S661vzMoXg18nu5w32r18WorfNXg15PUuwOeSwyCdFYnBaK7R+6mulb
UVFUdcwkXbZrEDhczg48iMII/kdJZkh2Ci8kk5OS2J07idOb+qqFpQsK+53KXUjdi+3T8quSWfqX
wD/PAgZk3zQ8gAvaZ8yEeEOGy+PcfgKcol5tL28vIFNcZtPnK9tzB1Vps4gOh5Te5vJ9HPkZ6E+f
B6tN52p4gKA7dC6KE0baSRTQQnU+HimmY2iXs2t0NN89M8bbfgHj3FcPfDqjvMYzNCP1O2FsbfwJ
kLWoPTy/02/A7Ljjsjghnb4t4iOhIizveDjnTa8mLdfrUAV0JW1y8f+YBIVb/v3mgLrF6jGU6U7m
LBFB3CDpw8DLmrZeA9UZbJY5gyjBN8SHQuvgxoxBCu4cCZusQv1wpxEK95/v2aNNyg6j2QC4G+wu
gpIuXZqOXtOdRSH+8xxBhaQ9Pbcelvyc8CMZGv1Ybr0BQOW4EqLK+eFgxki5pCmlGRGG0/4KyECV
SzLdzfun0sATK9UwmNsqVMIb25NDl6ShfGvJxVVML72dikTGAkO36EgNHJsx9QoCFMuAYbbGeGcC
XJBIqDAFX+re7NZw20DfrxDB1gLESe+mWTun3rKstpQEGIZ5ukrkaYZypgQSkG16hQR05FKJITsS
zSvHdNggLvFiudmC0aKwco8d/zcQZVqAaSHIeVSGtRuaxflyjlGavTAd1dV4nys+08pAaiocfghD
0HfGQUOPMSRpuasO36RLTuLRhYiaL7L+m/munyilf3aWDCfuzNGAeYaciNG0QYfyAdLLnsGvk7rq
neLJGVAHxUSyCafxkNqNXB7OtAkxVPC1K+eRo8NdkK/SeYlpV/6fX+4zEdeDYcOKM39vbwQtB5Hl
pzaiKNu9PF4McJG1/Mkh3+M/Pzf6YrleEwWMw+wKhNQTSytrGcvudTgmIlnBgPAKsrPE75VRzNe4
AoNdjAMqVS0qYY2CMdVPLzY61nOzuENkWa27RDcFCLL4Hrps/yF0jIFrCoxlZ8iPO6+e7lDSnNIe
LTFwUR8L/QGF8biQFdwG/OyALk9FCAkN4FalOvfgaXScrZ9Em36K5ExiepiZSCyH+13pX0pt8A3S
Jgb56Pk7+rLFN0/KRczxmWxPtodK9Wmn6TB/rHG4DunWuaoTQt05XZmIA8eJDiXt7CErp4HQq8Hp
grmcd+FhSBlcVggrWHB0mQHim7VTqe/NBrRS7nhvxKXtQ9X1UdCmR2pC6DQgqizUAFPchpFML1Vn
IYmUZTDHOWGywbduq/5f/zq+isPk7NaDt+uidb+qyAKyvl5lCqq9b9cRuwGWRtrcIYeRFtnMeBya
U7Gi1Th/DyEJEZ3daslNHiLSkluVMrwQ3HAh1ouD0dhdO6bjqTDw6lUxK53Uml4Kwfal5EQIAh7+
ONfVIxCvNnMKcf4X0UPGNNDE0GX5HPZkIjcU9FEXwE9KG7TB/pMVHo8c64p4rPtlZl0hiocinwjZ
18ZXW+dSig8PRPMmKGNqrrM/ScpPSFMKob9QeU5m69x4r4R/36h9ES1x6xYraPO5kKsjUG/K/tsc
dubu3iE1W4MvNSLzP7uRI+3B2MTou+0WrGG/djCoc5k5qn+Wol4AGXqUtXfb2zsSyunqemczUgLc
mXqGo6GXJPfhPZtIiRPtCKHP1xG9nakMTn+DUnjJEEmpDiCHhnG96k3zIdppYr1It+MlSkpTLjqY
DJ5tva07/ke6mHDN0vPrTD1/xuuQeCJWI5fJ8aXFYumwaHIqKugx795IyodSu4mTC+PAa6G8jwZo
zYwH58KzEiIoRhTPKcSGNDznzRoQKgjWISalHKwZDPPYGoRmNcxzF1T+ezY2vschi9LLTWhavIoj
IoeQNSMRlvswNAMNatbGvsf/7J/FHVUIXXFkXfql3rNGgD04V/K5K5pyFa0UxI3bIiZC1J7nONuy
uXnd3BjIEohoW3KFGh5/W4HVm61buf/XnRbdIsSO+67RoZQCd+iV2iTbt6Sm79IneQFu01Fjif4k
W0FJSPKjSrOCVB9sZ1PK4EGfh8bz7jWWoUTuXJvNOR00D8rViPurwvoQObdPsIR81RLXI/ws2FnQ
qtbx0WKEZqNnytWXenUOOvQo9yBmwLk025nQz4HD7bjZG6TP59ZnUXoETtMjkPKrSt+80nTs6/Tf
GIFOZkbkdW/VeU65UNpWu+tq5JJ4N/iTMKkVeJrk/DyakCTWGpKqYuDvfQAtOwz9zNIsAsnbs8Zb
LuYtEVRxbfDHjf5MNDALZod5u2nRgf+y785vzxBDfxfa0I05IrZIWvsqs7oHFpiFILGU0EloyD7d
jlLRca5a98hTc46NHdo973bhKq8E7iopkvjpkW9eJEcOAwYqB6teSzitQJeXCb5BVVFdaW2fKPiP
9m33lZ1I0e3uUEplkCi6iefqi33pk3PIbnABYybCe64yNVY5ajo49tHHl2qY+L9b84xvXqxuWi/A
JG6NWnRhdl/cWWz0AmMpN4UWB4VNbc+o/6sCVOmCynREko5agfB58YIhX6rgy3dMVtahEySULs5j
fhsdqGFtxlP7cJsvgIvvUmAQPd2zBX3efsnJvYLTR1U97PeiGKOtX0HbStVb2vNAClTvqJoBWxnJ
PQrE5BGJXt0Qjt/rKG7JQWGWghBpUTxwV1G1wbGAN5hJlgg1al2IQTFRXjae5p7mg5K0q9LSmjII
gII5XL2a+7vYZVd4lJ16NihW2AYFdSqiSOYbpan8w44zW16FaLWmDQce5Bf60AdWIFRT4dQYm2cI
s2I3claaN9GOUZK3u5yq7RpBThUu8xm/IczO/DfIf8qweU17ogxfjqoLIwj6h/pigoM4yBDQwD/d
k6+VwLkQyi9P8y+n4XURmfksKWBA4Oh8e6tsybUSy2MmCfANZuUqbcvI3gEpVJYAPwo/SbHMegvc
RhhelmVhnxrP69hTf3vaJjSJI8ImePdXBeR+iF73dTOLWtVqkbupiUNoTpRGF/i5aDTmx2ztcL4J
11dwRskm5RRT5i4BmRTDB8BlVPZvfzgvCy+qUjvAEJOVt92SKoeaKqAaZIYHdiXVqKoH2gU7eJWR
gviC5Q49Zl1cOKVUgC2+63B0dGFJTIlDqvwFBZ4xzFcOJO/ClL8ycoUBwx1pVEtc0wpfc2Gl1aZ8
N296Fi+eqEylk4hJBFTtuBsyVPvqd6pFTyPuLZu9Z8sObr3lwiXxOnx6t1qV/1S7OcQPNYg3jFdC
62RiJaIaNT7e5KuyG51yBnCpoMUImmiFG9+1/ZrEIDTsv0SCv9SU+Al9rF1SayeBS4AxtB6IwP5B
4yDSIKlrmDbCYyCoV40R5RcALOdL6ihJr85phjOfJ5OPMCa8liDJFe9K57IE5ysouUMGKy2bQA1B
0BY740zg0OM/UXhSXlMmAzof1EhHS//gxEeCd6Sy1bZx7zwWi+6Kc7RPNoRuvSj28+C2fmi/qK+0
vHrlN4TalnhdnbIZsFFp1aIw+TX/JcKM4VCVRc1uTjbL7rur8Z9xFKuoinoe357E5Hl6uckJvRhi
zEx0dVbvvkno/O8i0VFu8EpLd0pq/s5yel5oGsuK5nq8K8WrdLD+XhT9CmCkAXOS/hZSQ7Uk23Fi
7vO1vFQpBPNp7zUJS9ZGlFpsrax6/oTo7rEKJQj+KBdwNLkXwXEkJeGPO5N257mI/NMFD3RISotf
f0D9bnuRpphWVKNj1O1Iw23aOJrzkFkDhVEtXetUWYKPYe7HpZRy/NwDYuejl88969qkeXhPtPW7
kLkmw18rRIZxV4ucyq5lu57/Fy0XNJPb0VewIP26Ih1Sys1r9oz5JLOYV9/pDELYpo3tK/j6/RqH
Z2mB+cv9nGTwY7Aql0kqn5txlpMqevyn2zXQPvnkmOUPfuWv01PoHjhFXdOh2R2ywhr41rB84Klg
67g08nE4ea4/mWbOPFhKAbfamziVIfsTmCrp74kLbdQrV1xn47yTwg3QwbPkwyeQLLAALb2vO/R5
de6JKKgkDtkljjMECQJkFvkGmIBVeIbK5MVz2R1z0orSyCYDs8h+TEwVnTU45C9/h66aPbm1mC7g
vtVFEbdXUYflG6cakP0vEx/viPNT0y9JUb647JHlbn1QldRaIoiDIBsZmgt3eKgkGibkLAFnmGjY
QARu1P3MFwbgTNldmk5RBEE1rZvgI4ACGXTBczdSbGBQJWxVTtoddAbPCBv+vO4h4UvBqmIGsimu
h21EK5WNDOhZYaB0/Gpauo4Gaoy7AGdtRZSV2Hgwhj1NLJixp76jGUiDiPr9cf44bYvDIa7Ug8VJ
TjlVlBB0pW+mKuvTJ5soJ3S5X8CH6rcQXh0shqwDveZGxaSiF0oTzh65gczHGsUPE32WgtboUYV7
iprNPlvlsZbJib2YAy7TS05rAacR2Kw3e8ZbygfPhR3W+Vy6Sum+uCerpAs2dQKSvKmEH2+pcsNo
ySud4NQT65rX8NLTFcLlXX/HtqgCR+3VIiJEfktO9P7VbxrunsPAuOZT5cbN1iz9MmLKWvUIABv1
Je/tPIB+y4++jEEi/VoRsANA7NhBQ0KzImt3eaAcFa4X3PlBC3Tw2cEPt86n3pesVk38+pYD5Cwx
xxC+TDZ4ay7e/eeHP+xXjsTHsFM6nJv2um7H41veq6khSXN/VhLQPlR0EYYUeKFkYJqnFCwkehLZ
CdgOWFtKY3NDxRE7dbS8JgaqwPHJc6naXyyLoQ6Zzf3LTDGkjLk7xOUIRyvc+TGHfrblexfn/7KE
1iv4C23coXAVQ1oV9nN4OZLo40q/yZXVc2M26E9Ow+azMJLHBcSSM8mhZ2P1c7ggvjmag5Cyr75N
w6b94KNszUVCnkYpEGVU1vCT7JzzBKmSm1jjOD91Qh1jkIwB6XQdfVZqaE4+jxazszWS8yAwOvUg
BJHhDHp/mKaOTaec96QgRGpJOLWfwLFU6n6mSmParX8tz2UGhaOzFdYhy5Mou4HcLX1Aj8bQzw58
cGFnq/zdhq9ahq8ZUuxruM2DMsumGfKj/ZEhteddqvGXkG+rPYrB12A1OH9Yg5X7Zy6wvs0KjztA
AsQl/hZNe2bIEqqZ1S84O0FL11jMT1ufd8kqPC2GaZkHMGaJ4PEehicTqqjfqgpNipmNUaLSQQGk
0qye3MiM9rC/rThY5f55gK4uBvGgA4eL3H2F7Wfgh6vrZNs3cx0wbE8ZzrXRuZVAxk434VORutkV
8JFieTIKIia7VE1wClbDAT88LHi36mCOm06uywj2WMgG9z2b90Nz7jTbJdKUxs96wnZbqZyMMk56
A8mZxIDGi0TiBddHG3g9PT878AILmNegih9a2cBLC6LKJMLxA1HxJuMdTC4QYvZ2rZHI7Amw6PBD
XcgqJDPtvkO14QFaV+FsvqccQZgjM12UpOvfBa43ROD9Oj3a8DcVIKRKzYujDe1vKQel+hWOeFN4
33W0vxUBDz5WbdrlCurAAZh9YGCY1KTfJwGhVpo/p8CuR79lcRzkYNc9qWMbDjZw3zHidZB9nNCO
kIi6eFcsZ/Psn/c6tv9996ueFa+kik6OZI1jACU9ySFYyVDXxSpSlcaMG/Ojnb5rCa0DSDLF2pKQ
IIVIgmcfNi/RG9niiui3YVQJ4eSHBX/3/NQWxueKTrdAN+1buETQiJtcWc8LKXQe2bOd0OnMY53U
4pyvPabny8B6UXuFq2M0XVgSxNWmOfAUvUJNijSt07u+54GIUHJO2IQqgZ3VlXNT9R/lESCqudn6
5EqzmTti2wDP2AHgGDUGwpC5AhCOXbOHqr8zDzT8dkR15pFZXLLUg9qkwj2+qdKHjPP67vRLB1He
OPFZSwMH0Qmf7z1sO6ScsNZW4HzOxrpZWYs6b1AKrdLBKQAuYRYzyuknRKHV2X/jdIae9w2MPiLL
C52Mp3jjcF3PXQBpf2CPc3l1EC9wbeuqLR/j/xwFUTib37LTsx2OJw42dHNYusZTfVaEDzyYkQRl
uTSUaAdf3a/p+9TecTmYqj6YvPJ+80QXk/UdwDvCy23qJi/fov9StoGwLWGYtHLeTH7896xRA0eF
RgRk/eiaLG2WEYWEG/jYCSA2YdbmWaNgcOhi/6shI86njQNfPeAh3OeWaY2bQuqEgY879EiNIRSF
bIPZzr+3gx8WNs9uFLbbL/WOLpWcAwxAgGLfvgaizc8vYBIkH0230h9270p6MzZ7rnaduIPNvvzm
qKqAU+HI2uI8VJeNjj0YEl/eBjWi0BnMPkQXxIvbKrZKktmQxw0KIc4JbA6LcDDi8HEJRJhvTody
q7SVYOEr9eFPTUzDVCY8McGCKAL10f31T/IeKWD+QFTMgjHDC75Q9pqtlfnPEheYP/RdDjOdBMdO
AK/Q8zPPavE0y7QctwzvQyRZm4fECyJeLcXlS6hvQIwM0+mBGvU2c2upPdodTvRw13JhbjMpqZLC
iaEFEe9fZvOs3DR0ljRsiQbIUyBcVL8iyWdd1sfRlOZg2W2dVcFGxZNviUVhqmUk1n9Q4xTmXYa5
O2OQSvT/ia6NRGvwAQ03RUWYcykHcZcIdhnD16DDWLRC43Dt0MzXDf5uBLbUjK7W8XMkr3lguIAr
y1Kr/eB6EljVceAYR+gmjzU158sX8qDukavy3T0o2ys1EWVCuVpj3NYQAgdWC1bgiTFABKfwRxlu
P1GZAJQ7teocmulhho9hiYdAAkwFJUgsG924dEq8JZxA1UP3iQt8eLL9MNrjEkBDU6r0/MPYs2H3
sWCsHSO+bd3HJDDxEgB6b1o0WS3rqPP6jbChQO3/RQc4kwq8zNlvYTQkw5p59ReVZ06rzYdw8ims
K9f+RS1dQakGpb9RXunotEx5LBesxjOh/BrPlj/g6QmR3dZdzhr8l+OWJPqZ/GznWhMWrvl0qvzE
Dwe1wSdkVatNxfdR3qmTbjDak1NBATNfMP/a0NAcFbhm1GIJ11dhBdeQFwW561ZeSjPayFDOLmBQ
m05i8XkULjHyZVbLMMjPeYvInPEz9vzFeYmy5DjkEJzJlv0E98VzVmE3HZfcpWaT3uMNeBTAw5gt
glNUSTjW1FCEPgspuLeoRdi21p9QIRA6mUMe8mx1fHPw5ktwYKcmXNgFalPY6HQGU/P46/EmsHqX
Ac0SfQiAv/exQGl6oCgOLZiWgRCxpjAXcucvJ9j6n8emtoh8WMoGF2DWsEIcaM2sIaOBA+sofy+u
f0Bc27Wjz+UVdfBdPj2VbbZrFlM5wh2bPOBX1Nvet+6U4U1VtH/wnJGMLB/p4/icHdlXDB+3EGYG
3qk1HGnCCQ2ZN26gZosR/fcLTfGC+VHp+B+YViAv3g9L8t9oUvBNlqR54MXQsivNBoWz26zioNAq
hPfwIqFo2fBU3akL4tZamW0HGNXH6cYKP/ydSzI2DrLw7RwVyWsFpu2DedvuQ1RciQTKWNGjn4DR
Z3WDgTmFY+UMjbtirieh2p2VcfmlTYDUcWOm4ooUptz9g2i7/RNTc++WNSUjdhL7984N0wIXS27j
WXyo1i+qqd68WkovFaS9xcG996os4tfZaaOs1yg5tSsiqdfRu8QBSJwUzupy02bJwclzGn4wVKTi
zkyE22cnq3on80P6GgmdZCpmoviTDFCj3LmKZeZU2e23XtKLuqexaMZqEkaDejkVnKmHSg5nxKQ9
NmrD/8RGZdwATD+TSBhaqVW3kWUyzOTGbmlLUyykgWbZT993Mj4THPSrAkNDwGTKLJqYsZl18tCA
F36nEcIiRaqkgpaq0CWfegrlRI3A5dloFKkGfLRlEt+NMZ3uY99sKL2g1Nt2hql47/umGSnaMVw6
QE48kgcdXrelkw+MWEK4SKXMNPtQ6KqXwtj6pSyev7VUGNO3zOhSppHg0INIEZSov4qMLcG6Wu5t
RbM3W1Vj94N+mjUHqJ+o12BL3/ESql1D16klzc2odVDLCVaE1fP8V/fhlDVX8TX9KNflhQy0Dafj
q6QTqg+U0+ugF1uiG7HQmptuPJ9kOuhpdtoCm8CHBx0F1u/rMPvwvnoJCDznXiUNVheiTpqzck0R
g31k9yzS0v8+iBUFyHF2Fhw03Bhh7LPyTDLKe3K8DVkdSrcb7e3xGf/1qNkCNTZOPUBEncYTHncK
PpXfJbNsYCjfVCJ9wXP2mlOI1m0e3lBjUIP22uSUA0I8o40j2n3BzsFCM50TZXhqtGwcayBIoTl6
olPqI3lMUlcL3F2YV8bIfdq0YNmRfdxAA6918/uhnBXNTtyKJrGAhCscBrSmHpmlRR0FgeRgkNzm
uE2tJbUZ/Vrx9Lf/Eskm0TPQyaytxsjvZkJys4QIoVh3+4xwN9bCyG4FW4mP29Ou35YiB/hjP560
mRmTlhetRVUgO852VpbNZeabGtNbIVnaZvzlunV8x6ts0KicN8QryCAXMmEG6rc4M0YX6vTJfhGp
KsynJb94TAg658q/13cZwaiFub+iYXw0HwFPoHgLVSwqI/uy5SKG16V1xJ+9wJyiPQS9GSOjeDgr
qcLsE7aaR8Y2xroyDuRuvIYuNhjEyloBIGGV5CnZV/KAjbo9udcC3IA/KE86VXIBcXByVulYXS4p
nQXBP0M4Zwe/qUwwWVdLWPh12F8xX9P48LhIUFCK7glcN9zYQp0q3juJiQ5MN0I3PYale8RgKaV2
Hs+Ws4vfq/Wd3uy2FUM2xZQsV+jc+19qUd//gBTom6L5zUNjhnsFp758x4IWXuG3zjAQXLQIljbF
SlWSMoahuOyIp5pApxtDk9m80XgOgOEhF9ox+oU4jm0ej3hKL8ikIjtfJAgwD0voJJMa3CFfXTMo
he1f8oYZabg4DgrGBn4V5MOCby5qeID/U3cshKia3Q51DI4ziC66PvnctfSphhKdhfNCkgV8ptfT
QW+yiJXnNLAh3ITdYdLoiP0yPEWZFwIcuPS6reX5qoJXuokGpKaqMS/mPY743/nIwK2AROn4lQji
izhvLTKka2EpazUKft4VLuVOPH7jTKGG78Dr8HBo2WSe9iBeKYI/PsTPNefGcK5gG8+f7D19ZFrk
ngF4/GiUPzVBaSyqbfk8YD75j3U1fwDeWR1kheB+OBJBcqfBsRnHUvazPlrYXhwxTuWhQsWI1786
vKOlQbxC806tAycJY9F4zBXGYjSLFh2gRl73UgUpPofeDopQc0k+Ljv7S7yJ7tG7yKwQxNxYcRra
P0+JMYDhH/fm1pCvalokk0QXY+VGTrqkDqDirHCWKo/4zynm3kM7fvjcIbHT3umBOrcw1yKuO72I
XoxoJa9wEcJQSbm1BJi2Y6ajyddF2wVcAq7Cx9I/fD3jLqwvcFQ1wHHGDsDuRFmkXu4R9moMeKl5
0/HBtliyMus/sXRbfNADJcyNmJRdTnGn7DgsLCi7RhenOIbp1rTTazILSnnLPNDAWiKZ6sT+zmEZ
3Y3MAV1LprDWSmbOrcwduAUgdvWUVL9jQYNJh4iRKx5C+r+I5RtiRAG1izoPt1q21bOTVFxL6jne
hJwQmPaC2myeGwTrR+VLC+UYxJ5N/GWgrkWPJCtiYwKu1fAc4qpp3dWad4CDFM1VBvU6f3y5osbu
A7LiOJfFmK494oHzJnR22HGAiedLf9oyXkhIoMfO0B4e8XPGKhkm/BofEJ1/l6Yzdjj4hYFP5odp
DfzrmlKXR4StWCEF/2iq6uz/tdsqkhkIsH0g6W73NXhpdF2sXlpeMtCbe62Cp0BiSDv0097ih+b4
JoFzeLNBLkrESRH1zolRHHb/6LsZ8GfyYia/qkn/JOXUHOsQvDGRBm0S7T/Sl9t9U41WugWQXILp
mujUymYBR+leCEFMYNMo9PLGW820hLPOVfIxM5or2dZuI/vtvZwfqn80HMiBjuEfZaeNNtmf12Kp
p57kzF+mYglXg0/ydQMMS/GSpVKjs6cwxxlM+XQvCC1+a4AjdVbPFEaUBFNCFz6LbPBWQEsnk3cj
ziykQWJCN9yVYVSswA1H+ueZOILRhOHEzqL/BbxGeFCXJkxsq6nPbYjE5QzrOG2q6FownWDCVbAe
q5ZxM8ydJYqxXOom4n3fbhkf/oskRr/yu+kg+O7q4ujigXrUyXftVWMKs6VzKPT4bKn+v+0tDy57
U/KJSwRlQKvbZfLuCRS23iPeEf7QAidmqmmW4kG3rIX/etyGku+CWwPDbKHxact2iS6WIZX5f/TC
rawXEMOqN04IMDKdB5bQwnoQ/Ws7tU27FyxLedMEuU1yTMsMBOBigAhKguPvhUlye95R9BaSOeHZ
wqOJONEGIz/33f6VNkNLPdUxHkPBv9bEzsHPO3lgasjLAdKe7K1mVapy1ED78x/Fa53QxLMgkd9t
B6LZaj5ch/YxTZBSo+d5AmLWi1ctyBTKs/1P7UdvkVxN4oHog6T69coVJpEjK0dTZ7UAZ/GLua7r
MVKWIM9fdw7/mGWj89TbHzTQwB0OHFvDzW5O7TKZoawOIuWej12CtZaWRH1g2kdifuWze6ccIC4i
DUm/SGuA6gImXRyC0fdt/KxftvwMElZYArS/aRlMSyXTXhdsmMxUxYitXRHeQj9tgg4BVcewKS27
a39ZZAb+VrQP4qt3cTqDMnEAomOCkVskAF/ItPlSUk1zbXj034eas6copBoPC85pAhtiMDRWW4HH
t0kSGY7G+09SeUBOXPJ8cjqLyp7cBAqbBYtVn5Y9AKtsyQEVcoL8X3MmOYN3T8WsqT1CyGEzW2B3
wpObLzSaxGn0wlBhKcu7CT5hWn7d4JUpsm5X1bKvpl7bXIeZd3tpsLGhd2Gygm5igmZS6C3AjDPH
6ZMLwLWCJbDb6jXsV4IhV2Mzdfc2IsmrfsQjQ0CWunXr1IkMZA+pHhz6E3UD33vPct0BxiD6hV5Z
YuYu6aV07eDB/v43cWArVSq5JZvnxocL2OASRyrg6DdJ+zkucXvIEzOyU3q+oGfaclf7+wxe0S0Q
Z2SIk86ywXNQhCa4+umceWSdUQ2+nwkSIv1TupEdJTWMDvVShAkdo2KOHviY3dU+kIaB8QOkq1Tt
0rutCRYzWlzHiF13qw0dWFl1ze3CABnYBAW+yqOlVhhluDaW7VSPNqtbwTfO+ur8gS4XJ8EALS1E
lFia5jbY7+KJ+sE94CtS+cXitiO6Tdhs8ESjzXYOptqaVSnkgTxxTRO6gYVduhYVDbPUgZq173j3
r7afwGQVAOm9wZtYS0UsCbzFiJUQeOIx3vHxHYEO4ga2FVPnblVHiM5mo1QeOOUYTmR+s/gi5Ym3
o8RxmfwZD9VVBDFsKPTqCzPVQvT87HV17WEeTGNxWqzh3qKfgzTNrU7Z48yrQE4mrbBifjd+8W6W
hlAW5f7iFteC/ESOvAgCZAbb/hpxNnUQKZdhwE75q6RgBm+8ySLYlrSvKvNP1MB9+8FBBi04iBor
HVjh5ahAcatr6dB2unWjhjoE7Vc9V4Ys++T/HKqTysRolISEDtlIt9RTJgvQpUJQrgs0L8Q6Gjrv
WZ8FxJHryhy2SgHUObEFH+l8SwxIMoDke5KB5jiBZ1fGVi+hVGc6UhKWYDlyOTHJvzx8X7a8YeI6
yV8FDKeoQbG/K7CjWTstqJg4GefkKfzdS5VBhAzuAYRAmv9dSm1NNlXuMb4zWz7LLHQTD61Sy2CH
Ky/9B8b30OZyg4eHDubCly6P4FXi0K0APbTjwgeRfzceaZFyYYcjo8dAJl39vqUqUUfPyt8XVRuy
SV5URP205stRmlXJDJzw7AQIy2/ixGugGTdBHzoQigGFz3FvRgcx+wiAO/rX3d1rKbGsH/Opuki3
cPoW+8w3/puyg9qg9BaPFfOcLHauY6NiLsnEy41OnIneFGPxivENlO3nt+PccPAp0kh3wKdydBmC
4aTo9tCmAXsYzU6Yo9fX7wadG0KLyEAw+wWGlq4XUmWWlGWjRsEHqrcvbTHNu/8PcrRWnqb3zbC1
EnW6LbCtfvARBEVMI5K4AkiSx+kXI5DVnwpWEL5A3sejoMyhf2bcepmXA1rnRUjG0CBdLuiZ1TCd
7xwxew/5Ra6b5NBVBaOzSjEl3+dPvyHlHltjMjajDz4drfe/FpHaxif1IpShF5FkcBMO1ihFBd+g
pLX4Vt5hmccEpNQ7GIyZhAhHli9G08QmV+PN51FXEZD9UCoQwQajhKVBNpRpExFlBSD6FuOp8tdp
pQ9hSuZoSukL7WkbhhLY73Mj/qaFJiJh7CjGd1QO6dkPQQ8rAECSisx8XqNwW1Odv8BoiiK+Nimh
iZNEAoGhefFGPMnTsYvZpk1WnT4zyB6/UDMEuFh8SyUNuHYUXfEYCvsGol0U6I9ggO+NHVohWVbd
4r6m7LTpjARIqzWw3f67AEH57dvWJtlMzGtpJ2IIi7apPml+Fr1yE9BYkjzYlBLuoas+lNlrBv+N
OifYxOKZkGLY22GtL7sRDe2m5qfChk9CJNTsGbWckGYMp2qtHg7BS/Mdo7jSYAB7XGg5Hzsq7xDk
Ne0SJRu0jPJt1zrlpeb7+FPwuBzBrDKFRIlhMEySeOplJdSjHzermlpT4vC2ZDpSsvXPDWFyTSoC
3DHGi5MpXCJ+xlntcnHJkcbw4URfODH5E1B6b0Kb+iHyoYqT64gqdSLHdzUt57oqUY4arsMLVEEm
TC0LlbeAImo2z1Fez+vGREHI31Cbtyj35DMeLajhXRIVv95DLZJ7H/yi/rwCZeX6ZSmK3JjYWdES
3ajR6o2X+kaZbwvVQpt+1buLc1HCub4YB+4rB0+JbW+bYJ5fMkpHk3bFC0oWXr+5+9JLqV/3gg/2
umUnDqHu++IcIo9xJhGbXa/sAwsMdAy14R1BbCpy4PnoHh6r+DU9ys7SOK0G/gDGKmlg84HJuWXw
1cz6wLQ06o0Co31OmBQmfvXQYL/reNLCYHHGO8OgRk3iqNOnY1cRDxkOMEdbMofL6T5Hw01yzuaY
wLqf23k/7AaiR405VCvRrzhOM8+qDvW7XBRivoZg0HUUC1FCuRpVvsQljY2IEQjCV77TdL/3T8Cp
h3z6NgTMZ9XSD160nrCPua8ZdHW+PYT7ETclTpF/y7ZqmzyyTHEsZX08pIlftHjtpnHgh7UnF35U
8Fq/ZYEEq5waNlHFRQbj/MLgGvprgYnljNWw+6PfnS8mWTRDqSCp2CJKwqtPeK4xTNoaz60OyeYG
8Ek2/I7qSlwDU+L1hRgyILFRRE88MqFRpM/XQaUBAHdateSZiFFTorlY4FVj65E9is7/AydUEhvr
BvirAlBf8yBE/nJJvO9meEu5aFgFnt/FiXPpkyY974v5WYDdwPnN5MdybHuHNp3wkllef5bGZEbY
hMwOKhja7AXawsVyWigZoPGCcxwFYuCfRBdiFQIqP0NZWwoaib7KdL/8TvmHKHhjz+1A5fLcnYg4
wPHO6a7PYSYSOs0Ut15xEAJwA0xrhZu5Xt81Kr+KoOLBq5nt/1tNxxZshlqzo3Rp7nus+5+0JxGa
5OOxDuNjZEfcxdgs/aKozuwyYyZN8deRrkyyPGph0AwwHQKvtS0tA9srmxUxlyuiLQAYFWBk/HaQ
LYk4S1wTzv5z2KQ0TP+Yo4OSFh18Q+fKe1M43Ex6YGSUmcjySfSDfp93WeRP4VcflnsuASdbNTaP
DLJrUKtrHQI5OwiCqsnPjCgbcpWGGcjgVi1kNDu00YrE2WzEIBC177PFucKCVYpCwrsLTmhSuGk6
emzQ6TyLbBfCDWVoxz0Bsbx0PKX/rBi2aVd+xesoZi6k9+An8mXs7E0fjlxd9wRhNg0uFFc24qgf
qnJN6Is64dW1TBt+iAD0OOBiSfZ2yQwG9ofXjBql20tlBE9zbcOa6QBEr00PBw1YOzjvXqq0Z8D1
yMeppogE18hpgPjjevhGhudOuaaPU/JKScnCY7KHDo1MV82Cx9iJ89xn72OuJ2No4qSb9Vtr0dk8
9TJUavieGa8tJrJKblKoOkhLpyKWISLy9einXH1P3cI3MwKXniVcDto6TvX5zXo6eS7tEQFW0eAj
jlAC7l6nxMCsgJQhGjrEDHyq+CLXDZId75fy5z87pfkIzIRSFflx205ZzjbgbBOnRvWz54MHxmD+
bEUxGLRxFX2vjerQjJkGdDaoIMteYd5x2m3iBh6Wj95fuTvjkWPK0CMrp93MiSKUD8Dzuqmm8Wl4
Q250GnHauLE5RcNBgtOuJn63cTNYdJ+RVjp3UktpUEvLG4v438LOk3R/Kd5kJH3AjgBRtkP1CvZu
Hh/THGIYb0Kuf6SDOZoX7vvMQvXU6mA/AuoYKTV9geR7c/K1NYXYoXF+a10r8u5XGd88yBCCJ9ck
IF8/14Oh2EViBRWzCm5uzO4UJjPHqY6Bb4FXznNj0mjoqwUBtUCJcOfBK13aDwkVErx8KspE/lJ/
Hka5ri30HJoaCkIABgPCZKDI1V9dAiph2xGfuTRM1Lv14gdMFiYAlTXR7QEq3OP49yapDELI/KrL
RNh2LrzXLYLGkWDH5DTLqFU9KPQggoyL6+SztkaCimPwCEOpzg2ckl8hxyV8PJeXvUpafw+g8Irh
GXevXMl66kv9AKbVWt0Y3TospDV6dHqBnOnh2Ome41GQCZ7p6FqTPntL3Uph+jgDalEGXo/4mXnY
IHGkbftXQN6slQyLVpmftKV8JYrRaElfmJAFZtG1cgTY/BJPJVOUOgZS2oOFr7ywUhc4Ifu7zQXm
TSQ8pJcU11kLIxnL6FrVguMED6TxXUUNiFg6HGPZmJvhCLiqFbxkgjEDpK/ot3uozX+Ubm8obZDq
4f5lix9Gh2u39VJ7EExhzGB3JLgnabUKXXXm2ymm/AcA2jlbpEAwJ5PJ0mBZ5Ig/nAX8xb7FqBmM
qJqXc9Uqg6r/ktIh9DIKFNZjKavTsuKxj1TDp4GSegEvHuzb1VGz+iZHkHs4QhhKMvTuhKm9kDv2
ELXNbQ0CnzeMvyoVE16ehBNQYupS1Jrm6OwNiLfBY+Esz9Rz5rm4FchP+RzoNM+qEpzqbLViTJcj
Bu/ncXusRYRTfa/bardYsA1/vKQIGrWyAs4Kij/RLaoGtML9GNqSipAapwGEYQ8qXqfT0v9V1Y91
mspE4RVZqmVjTRGGk3x9ygfWRfkHdU1tCN9EIt2dnqq+TLH2JP4RVYhSOf+JeZZtG2hEVGjq8T73
9KYL8sJ0FDFuJCnM6TKN/ng8ylIDOkuljYxI6JzzXh6dTvrc/lOdPESp/fKyCqcGobA3Leo+ahRQ
x4z2Fw4dMt2QIURhCULpOjpBk7FsP0NQk3cICAytpadBnCq+r1JxokRGXVwLghppACkxjYduqNb1
euwEQ81M1zIUiUYXQiPDWLVNYQu9ep9OZdKZdPNpz+PDAA+ga5xunPlhiPD+igdDmeMr2RvpByKJ
j5b3E/YPmPMgxLKtQcqIzdWluStAJ9WmW2srycqbYR1BeMUNNNdfPFzxupHPRDrNVBGdXhKgXpj3
nDaI4POHx0sXKkZX831XMqZzLgG7y7cqckbDs3fguIVciSgw7r1uVzpwKbCs/FLZ+SmaEPyXPB2p
I14WsRdt11iNsQUBmVUtHwchK0WM6wHH29vhbMC+oouqS0/0gsj2gHGESBYywplKTyYL2qpgMTgR
gcCsEvuCZAvp0YXkidSvUfZA4CO0vngnHYQ1/9AYe3frMjguhUGu65f5T7TINb9vA61iEeOTGaay
0SrW+P5pdCK2I2fO8TV9qvP+gpGSd/vaLH2uhKpwB+5qM3h1NNTNAsVKI9C6G1VFZ9jLwCUUNKb4
0HkjsTektX7CjP/DDSokTpx+FIyfN0js0R93rut4AhNSf/lfjg6E5CIrJ/wCEoHIKjzIYaDAAXVJ
YxUz5QR6n7uHDUFV/uy2WXqBFEcJ41UMcnjuN8DD/3Ald9bZS3yTaMPbwErv8OBqU8VdB+fE+PKu
in3PhQsx/Y7+5qu1UE/2iKijRvbHgGz/Q4T0zXwwYArM8cCZlqJr9Sty80a/H1ERRWKDMmfi5TCU
79HZ/eeSVTPySKfaL+El4tA1GsvZ+DFMvxYGUDHR0DbcVEpL8zkFpQFctzQI9p6Qbqo6GU5Yk87i
kZ3YC0HJQjkPZqCs9n/VI+WfPCJVOCVjHmk/ZEoh0KW8Z3WT4s2S69F7sZKUXRYsxDqboVnPGSOj
Zqbt9wBrnAoFJ0vkoIw9p1L3VrGMxpbw4DtvS08jXcbaV0NVblsT1oqQ7cQv3twmHWfIf+4q6T3S
yZ6JF8tQMwXywT310GLz0HSwGxwnO14fDQFPddWLy1PZ6PtUamIUZCxAMXYxDjkcoP647jjv+0uA
iOqDjwzpgM9nE+S8bzgJwBY+0yZ30GH+/eQizPKWT5DcyaINZ3dnzWaox8uduRxEBZ0HENl964V9
HFqkKGDUIn2WV+TWlg4qvvzFG8bK4tGCYZ91d3G8NXUV3xRWI9XmWeYfApTv00YTxjELuRZyT7Ns
jX3+nIhX0Yw4koP8Kt+eIcRoTFb4UaHBxM2hliQcV4H7GUw3d5+7NAyZOGZuaGBNZYXbfws6/qG6
D0D0kC63bhEaOiD9xSQcJJVpLfRVrYzpUwjzGZptCLhm2p7XQ55VJbyRpZli5QSJmv5W2+2S4ulV
5TDF5H6exYajJ6bAok5P5V361jEdT3/bxn1GvHHjWuYdDyjC03rFwtIFPr8p/QlGFN716iwakh82
7fN3L3+IGexPEdtRt+ZDyPQu8x2K446XlUWiz4If3R5ZlJXe5Fy7UER5f7kGFyVEP2Cz3ovlrqQc
1u/x9xs0+CNSDJNEBDRTYg9kdMcdp8iiON5LbFl5R542n8tfUgnz3Nf0GuOg/gPNThtDw4vu3evv
JLCmEeuT7cu9VjwiPIW9kyWfUUuAbqe649a9DigdrjBt6i+em4uRKx8ld9ZrseeHIe1g5oWN7kwg
rYhQ1c1hI18GhxjtmdJQyNT1RJ0r0gbDs8OQg9qwCIwj7pHZZae6qNjbJIEdTGDmAMqGX2IY3Rjg
RZkMeXBnyang8Fc1nPSLIOUIfnaokKjIbCJCmikC41s6/VG475DgcM/GstMHjolPBMuDWJ0C/8nb
Ck6qbA1TkmkePyDPHxwEDF9xLrZyLHBa0pdMai3z7rAhs5cKvDJfNpbkrumw4WKA4Aazy0Xl5t+0
8Vdn9WOFI8sqeo05EHq0kiRDaoe0GgbWLzs6DIW7HMBi+AksA3i9u0uLIM1N/zGT/W2MESV4cJvG
uivuSB+G6YPN7kOsk+Wjs183Rg/qY9ONqMZ5FEFkq4lgNlsraZyVsALuRmSfN0nxi+dZo+wty06O
BbDSDsMYmZzDpQ5xF6mb8+Qxy5jywZG6U5TIbCBk1ufp9w1vGIiGhJgsC7PV3r1QD684EjZdZcM8
oY49nxewLATm4ZNR8432dXqUrgAmTrg2euVv4ZncHNLXnaZvMjokg27llRh+ybRi8dh4HBpdkSf8
b++/YXGpLxPQSblgk6C3WE+Sd/N4t68EOUUX0Bo8pbe3l8YI2BWGYk1dT7DlAZLIqwIhaSsLLoDf
JhUhmkqMeaSUxZmUNEacqA3RdsEeSW5ZBfecRrK6FO0FB71bYPvxHYBbTsu8XtJmMeFkWqHuiFjw
Ak3mkFnmvPbNSB8GrerQRbKZATFMWnc/ZzSU0HIrh/Sk5g/d8nvOUxnQqj2kv2uTvknDbEMVLvGi
KxDBab+fpxRybDBO+CReiJB+9GLNanZeJ5divPKOMXDqo9p8SOV8VM8VSwH4pP3U2onVMW3q0VFS
oTNsfMgDAU7hqdARcg/zh+KTQdwA81BzbN7sagYTu8qMPampCvAxL0gI59gNpv3lk4fgq7xBRwK1
WOCD9te0CiYJjddUCMb6sZNkB1nctEpM3CFPZBcy4cxRuPUecTbq7Rr1VgtPvJYqUA7Pmxq8Kri9
pZwKnNv0FECF++tmHbQ6z+YHxyCRP8Hxh6EGDZ7k3h0nbTj1XK33o7WnvQhZS8KyV2jVfmPBDN+O
RqpqGkqnYPwBnFd4KuG7D5brHxOmNITntjpoFgIYXtmZkqfPMhlTqnIrBLRKPu6IBu13pEDE0rBo
Pyhbv2dk8ahMCGISRM6ORhu6wzmgSH31keTlMy20ua+nxZHRagWtKESy2s3dY/Ic13t/hDPfDgHj
LArVB5kH3tUYdgzv3qpSKJVPhl3X+pXzMpQOUbfKykf7SCjway+FOnHb5pXLthNS7yPIq+iIw1+W
f2dCHN8A7O3EGU1/jgx66Z3VQx6TS5Dx4gAO2BAjYJSO4NQzqd89Yj3N3RRrszFeG/X8GDrM9K/I
cJfSEP+9K4wRRqcvU/XIOiDJFkkgG1F4I9jshcH17dzbgdzse8Ga+hFddBgIGOvI/8/XO9XsUsTV
vCYLgzeLe8K0tGxc75VkJtjE9ojmgjgh13/ZBu+VVEhW8WjrRamKLKrzMuav8EIHXML6cptudlez
JkCqZwuSj6hh932OmcwYp0lJuOT0aGVEo31doWE0+sQaugSCtHbq2lwJOgf+S/gSRjF6jrxdvgA7
F4fuMq4xPQq1gcG25rrHC9p4umJCpKrebjXzVDyEJE0WEdTDeo6k5jzH75QoZbtmGR90zSRumiKu
R8CpZnuQdFzE7G/7KsktiBnnNdesO4SEj2vw1sdTWUzXWGxHuwI0+cQjx8V/KQDEElwuLpVxqTp3
mey9523jpWEI3X/mGJph3uOcWllYbMNMiUf0HPzNpAy6TRfahwYNHbGwf+V+jOdrecJjIYyByzO3
YpCwAAMo/ohk3q4OS7S1ghQcwG9JZEKbT1zAxcyV5GichPFfP4IZ6rGaOLF5GOPpVXnc0FmtbEQi
ffUDokBb97K/m4UuBXQc3xVkra2FGLX6DGSV/SJ9/5ISCkPIL/cGXMPP8EWop2cTVS9wXJJS86dC
ch0w9dF0RwqTgWcWSSyAYyqr+nmmKUAlN6/k9OVxrK6aM31DwUvJYpWRp/4EByAyH6EBNDX7k/7g
p0wokZAcULfzhr6KyngxRzrLA3NIlC1wFe3j4skgJVEbxKlLjw6FuiQpgj30DoG8OZH4FGcwYGxP
Q8U2iQ00ss9D8b11C4/DPkYB7JSB5wdEjlfrZz2qLh0JN22NEZMOoxJbu9Gb7AXexBW2v2T4Sg/l
Tv6MT5FOPfSO7yA3EwXOwOrpe3JyJurrSZxKoL7eHgA6cnceHFe8CWy7bIVf7fmCOKKKndgpU8sZ
g0ocHLdAz+zNumjNFf+WJEea+s3Pfv0iAuFocHPMnWB14zMXY9RSKT67+ZeTSzNlMj/kHcjhssol
qot8Nuxa9hqrrsm46U/LZp3LdpOzFMqeaSHwNE3YAfhGfB5UWO5EwhS02IF54xu2bhok2sxoCtMX
rYEl6Adevc61DklzIu3Lntq3CzIeAZCXpYyjlvYnW5LpYygEvQGrCLfY+Fu1GIygl9cjIDmdJX7w
JZpEzZ/WYTMhr0cOm1T6Kg/IUPLO2Pyl8k7a8xVC32V718gNz4iixCH8FYm7K9wLRUFOHhaF03BJ
RMNFM2IBQ9AbJHd7UydIoNEScZJkynB2q9WSz2BLopVfFE2WARrvtBkC9KikjGd+dGNaLAiBvueL
lOwGIxCEx5gZdzUx702wER8I80m0QjFVLzMUL80ZMw3W9G05CXw+0W09+QkZiC9Y/5Gnp0bGaE+q
1iJJgfV7b7DcwlAbo5UgGr1WCLhws6sio4YXXL3/ShoroPCzL6a0Ngz2jG3bMtOTfRqwxaYgOHU6
f8JH0LmSt6V6uX3RKDWwncHGqkEVJ2eVnqaGBGewDw4Myj2DP4jTjIAgZ795xWND0nNinYVpaKbE
RQd+Ji6bouLUo5Gt6XISDHwNA4y6CB9w2ZYobMKgNBwAw72iTetyheACeEm1Bf72r3sN1WJE8hMf
3orXmIO/pJIYTyvl98AyFxedkBQ72Q3fBLgwfvjiyxt31YShw7K7PBXuYX5kT22LXmct6wWwwtQE
VQ8QM5qZr4HIZ2Ywux2zyB3SCVgsanfxBX7rrpnNuFJRrkodaC4h5xPIJZzmYb4U1K+Hu+CBAnWv
lUkadQzVHXFwFv3gQbjl6D6wYewhO0tdT2sQP1jdxrPo0Clf3+Ak645pmIHdNI0/2mkQ9pnJlY7Z
zFzrOYiPWqSRjvwpWG/rMjJcru+Ns0bd+zB6j4Qzldko8VMLCufjywzmT3lNcqxUo/k6DYWOBidX
pXoAIlku0SiIbVqZf2FJUp5ijve6oZR8+gyE54w2CLsb/0ZZqf47SwyonvY32PT1jMIWdt2JRUgt
tOIx/zu5yLlfnGqR+x/sJZrjxobdXB+rnHP/9jM8x66agz7iqaLRmVeBy29oipV0bt4vtgFNqgLO
AhI8ROHLgcf+Yfcm86nVgGeAqGjxBDMF30aHbixmi8bZWclKfp1PY5kfddLkawjGYkgUG2kUGgrl
1RMihFMC5zaDtwObrOzXcs4Yg2uBdAlLhYNZF+9a8F2CIXB4onf7+vvubz23b7n7HOYLav84nXeU
Z1T+e8N7epve9Exkxgj4qXhNKmVTZVrdkzV0ftgWF8/uGp9as/Fpe9kf4JU8ygPJT6pgFOun7n5B
PASttEdm4JVW9vUdDiT7Au749OwGpd3xLSkjnPXxouHTPc8wC0dKhmazSrXp9FvVdborEljn5sXf
60Y0GZ5yK9GSQqmUBFQntCtQ1zzI5TxdJnpj4t6nMiQeuxY7HyADL5kK8ohMWDqaHKuejADwdmu3
EsorqUGTD8lor4WQ/ix3IzO3TC1LnU+OfOsw5rN7DPtkKzzpmZ0CQKKCSoS+la8mQm61w2134Se8
dPCiO4yTvQahfNRuOxbi2ydiHjar078Kwm0ZDa028r/8wHPbZH0ufGvlLoaWqdUhttggy8GgDMB3
17MD41VknNlMFOyrSyn0/4w50LKrTEcj3qyC3omF/ReyvEysm6L1wyg1/wo0kMGyqcLU4yvFUG7f
3ozDg8reFhzDKmfQE98XirQi/QDmobk5/RSp5/hUI/ZZKgGdOMX858hiESzkMY9kwjurs2/MAufS
TSrZlq6qGOdiG+l8hE515WmElPmJsDVZoOg9k7mIIJy7fLShzoOM95bNM2OlVbf1FDPb0dMRDDwn
vEZLtqlmYxeGemY1P4a5JD/qRWsalT33BwIoDFvDezW6ZmruQJNADkxq5jw0vuis1mz9ix7sBwMM
duUNLVzc89NTaMccXGWJeEsn/V4HJwQWK/7QqtXMAJOI85CAPmRaTULKRyX2APNZTQxY/F5UIVat
HEoFXThyVmVlufD8I+6xjnq/vPU1NVPEWDChUFwO+O/lNY5H1204R/LTSYyRRWpT1YWGPT97F1YM
l22Qghfr0EaXHvsUvXjeSvJr8ro8TXDpvmPzlOI6/KriR6vjcGRAo+E5vyVip4IGHJnt01k4MzoO
UUKV42v9fJX8Ybx6OAtqS/Wx/aymaw44BPDMT/60cBOD+J9N5msH67EXNYUE+ho76Yoye8XduRQL
nMtbDoI60jq3JTPkJKZUWo/6LE++46YK4Sr8rHcuiI4m9yPESplcNPpfpme3OpQZ0hbJSRTpiC6T
QnHOknJT2NvDbQWDOr+J/zr25hirdbV+8bwLbjWVwoG3EtXHxwWtEc8T2KVcIskDvefeOckOpIvR
1giigPgVl8HJsp1JJHEwVdPflbxe6WA9cXHjTZOREONxFwheLBxizkEyyduDy+qloMu0MyK2YwVd
yZdEK4uGtFPH5qN0uSTd/3lSI+v/UbZudrtbPT2u1IW5qs225sl0974Kfm0bLMfveYygegnd7+IB
Y+pL2k+LG4UiYvqJRXy6M3A3SdiaU545LCL1dFi7CC7snGmq1d3AbSUp6Ohvoz7i8TT1kfcjgxm2
ec9JfP9+/aDIwYrMzotkSgi+JU8scF6xIPn2NPiGN1Lpf+bo0zVRdTBFs+WziRd7jmfyXekrTT3y
r8EJDzwxUK2UA3tD/xrsSosQw3bvFPSLqd7GfWrsnNn6yLxa/AZUt+aMj+IrEK4JE+TqqPmBocjp
nnvyeMZjpkzJ/PFLMosSb+60GU4ZaXiSz2R9aAxQDVWcu+KF/9UJlYIHrOmFi0A8cGLuef/BIizj
w4qxYL21wvdHRepS777zsZgIgJq3U+XILVbsXi2XGE5etmC/p/1V9aBeImbzsGlY5DscQ/mzafhV
SJ/p4LMi65ZSbN+p//un7LheGBfnXkAMIJE/jtxqSmQVaTo8l9aJKjl0NDPGD9yFBqrFHCzfjmXo
ebeSZwKWoDAHfgBwc3FmOFqwjwSD65vjVs5ToSy4PaRxvmznScbi5iLjzA/XWR9vK3b3D+P27tFh
YzNDu81fGLoSold+W5CUSUbl1Zs1hLst2PwvN10DqmavqiLv0WWKiIFqWadhCzg9ZpcuoI7DUR4v
+zPmpmzyoOIPzE9TUah9RHJSwM7iyI7xAsbBbXtiVXUbfCkChnhuvMrgyoWImksZc+zrvrEGqg4w
Tji4/VOhoKq9KW9nqEz3+9P9lexudiVnHIz74b5Je9tfNRxhZaRAsbHrTzfpouzy6r3SpEBo/2MX
98AqiDTTo08elN1A6fIqKehUhLpEU186Fu8U8DigfyXl3ZWYR6LDK82ofXjaYuqg13tjXbSyZFXj
joEm13KdLNhE75uB/xUYnIejVopPH6cNvJmMuWkuIa1vVzbXSPoGRmMt/XX5rQF26XGfkXfWFfBS
AfSLA7UInqtQ9fhdwGdtC6kITvLmlkMhlHN1E+Og/660sbIW38la/bfq159qzaZwP9KCPQerXau/
BA57aAgNAuTq/rKSgchIUCYeldzuxaA5n2T+lYuc6tb9rwMCV6ia/rH5eR5IVJOqEyAtQDS8FY+R
vsz0CiORE+q/2YSXRkWG7eoxKh3nRlAIsasDhNOaWsKQTs4XbTcnG5cGBj+5q/CfSzj3cIWhyCMy
njKySZP0nkBK8YrPgQKfHamrrGEmf+KqebgTDnIN+83MjVT+NDtShkXhkG1JENVw2mSKFXNAYfqn
ryI22FEa/We/o6sCp4hzeZYnw8OkhYuvmcNxpXESZdHVNFL/fKMJ8TEJ1z8pcMxFASdBO7jg461k
ZUCFsxxBUc9eX2mXFk8ZnykSx6DKcHi0/TJQMb/19KrXT7lO39pcpv6k53BuOOWQfZrAPgB/Uznb
n33c1/wg5M9TqtVdgs+u6xzrwaMEIjJ3ULkeNCi2LHPEy3RwT2xN8o1E4KUDxrAIJq7edBOm0pLO
1SwnQIezbcvZT4NxGvPPWnI3ysvxwDwZgstp/I07mMtiFQccXTMXPiBd/DxzEdVWuuie9HfR/frV
ypmxD+ov+VMX8V3WCwFhoSRoCj5G72D2TGmyN3kBc8uHSStRxrGceDa2KWJXUQQpy/KmEsbaasVl
kX0RktVEtNEeVi5bivZ/eTs3eHRHnOA0ZKGVWt4GEvPgz6u20z+qaIdS2DcqKlcPr1WtW3PAXBsf
rKH+bsDKYN4wLmbHRGx9YM8782Cswt4DJue4mmESmODlis976Muta/BnXxNgz30TFMRIgesELkI6
zB7ckpZ26TWVa8pOmW8JHfLrMAQEjTuxA+QYczxZvKODWhe58kfaY5z9043YTxJ8MX/W1I+4k2bL
XIV+ZtAWc24Vy0Ee7t8RktGvFvhRuBdt/Nvg4QUMGwsrZj0tb7Hhn2b/Cdm3nLfmSeb0xjEfR/Gp
mwJVj9J43kz21uyWf3OrdMegbPlZp9QWJYhE7pfu5ixNOWBfk4WYy49EIEDGJQODiE5xCTwNQrge
Qk1oqnxBXHd9Ioh8JL3SPJT2JrpREWHScuopxNpqO+g7U/LIPPU2zP4hEPNvvNTfS3icFHPCbwAg
TQSngXpCp8XYy4bMPETEJBweoEtQqtJMedY2JLlcKQ/+aiblNH14uOjHI7iuVivEGtrwVWzx+0We
qszvOQApZ0OOyHzfd4eh3DoIOqLw0F2n6HWhHMPO9b5qGoBM1fsiL1KyTEZf2Cy2hSlnU11oyDmm
iii0HRP5TdIoQnPJGgDINb3AUdFXpxSxq7frhSgA0DQlCTZsrRQbegEtVz3Fy/V+QYRy368ogVJB
IA6PSSk65RIccSR0YCA6yROkE/C72SpwJXKJWJWYvBnGAIVxvFNEkJrsOPnUx3FSWrBeI6BPMpvX
dWDj4z7Dpk2owt/HaA7CahW9DQ/ik3Ix+7tcPlV2c2PELwbxDv2YmYtzJHhtfp2UL8cXeLb82BQk
RuXayqhtjTWlGfzN/Np/yzTzX9A2NcqngyOjGvM/3QR9qnh1raS5RlAalZWtio9q3OcAsIuRNZpS
TNFfusQk2XQCrubSnks4QSH8fj9NYLHFjGB/PrZzq3/jXAdLrKSbu+FUDNU+4YBDobGqrE/aBlEQ
OpjIXiM48nLtUyH0mbLfxMVhwE2TBxwKfwrC985J71oOnCN15JPusCh/lz6kSRvGH+4vMMuNmSj+
FYU5zSsy0H9C0UQkrXwfIv/wCa2s+MnRoCOOLjSCg292tUkiRguJgXXCvyn04seTOaftKG/N9THB
NG2wANetCg3Hawctq2QknWFpXI64PHb0vkZHW8hmop+PeiZ4A5h79oGvkpseccfIb5DJNNZ0NsIl
mE97UN6Z7VbvYNtu7OquuVYHwhc4Cf6fSQmO2UHziux2XrOUykXglrcsFp5mU8EAd6TcRfq1bLvH
UfPnzTv8QHJ7/NaUPcnU4Kqfpw6jLRJuHrneKxKVHsXdCA5lmUT5kgUQnWNEkRF9ZoInoaj0YDd8
KaSdKvXyMNlj0HNpPEpuxDtec+lWjtk4IhcjMBJX85F2tZHwW2sArO8z67m3RNNCodxgAkPRVFYN
6+CxJVK0Ck8vb/DMgtoX5GEvhvwqKh2jwm1oDfqqryr1AlQQFrOjfspURWcI5WMY59r2i3SZPbLD
lE70y8Va/1EHyxSrhOJpz9FQFY697aRpt22TMP9JVhmczIPEuc4IL0oLx3UOeWNRzTfgMyjI9pud
S6Z84xRD3pV6OSOcLim5PeQyMPnjDAMT4+QVuJHqzidf703OTtwL5rspmJN6oYRtMRuMW3xAJYpE
eOR4SsENMOIKPX7GVXOfF9T//jBeAfcMiYhfFoxNrWw4gIXGyicQ76PFVoBUZDwmN+edHcFDnFlR
bD6N1VHW9YvN2qwA/otO1bzzt8ZpVtSZA9RvFuv1D3auFiyy3+U9VZzr5wRNORE5qkUFW65429lq
7eJAni6BOz/Fxsp0xsu7ji/mmaulR0tPRcoE8v4qdXEpyideW237wO8ZUa9jjr20QeK6hDir8ivv
kNrySGg4ROL3dnjaKIPDblAqlc9JFdTkLS5Cj/oHLomvmusgc4uUZ5twYEsVrNt5o1kf1hqhaDwp
+c31Td84VpJV3Z2VXxgQhxsvj1zrkpMrLmzGdG2wM2CjWcHtKfMYC0J5kpaD3wLe9UXsLHHMZU80
+rtwIHZ/CMt4R135nXeQFR71KyMNyk6Z2XVDq0reFiFvpIBKGznnzM+Nm2ZQYYPJKHX106UcikH7
HgTV+5dIrLX6UYT6mtVgNSiPYazEd3xa+QFXC4lIwR6NmPYxmHrkze7tjIkx5+1bPyenOXNeSAtY
+GsM/5mMFE3edPR7CBxtRDpickoI9r0E+AEpbZyGifNacOHk+pp6r7MZouq9uRvD5JiYDkqOtmtt
x9WTfT4N093cmapI0jvuMZQnk0AD/banO1XOYSoGBvCyrwmQwX7yIvTnVaiwKkNcor0g1+KSCGyO
BAlLVp33x+KFNUFvr5VnrJK5Jj9vumz48Nt8M7dDKcGjh47C772BXMME9JLB0yS2TFpz5F7PKP81
OgbjAwVYV1kDLjoR9/dtV7qlpACkSOq68RX8TQCH/QvWExNWJOpuWCGT4XQQF7Mhb1DFLU+EJT1p
FqbTzlZtDo/EXjoHJoJ46n1xcMPJfkOHqBDfuEb8IbsT3iDE2zruHk3jh/lIOm59cRgjuZUPouUs
iwgcGyYjmXiW0vAoVk9bPOpDm0T9844vl3eKh2dpTDX+o+Nymcn+cgXO6Si2riEwhxGl/vUs8zG0
ZxvEepIC2oFChzuKwGQ2H/TVJecdG9ULVY5H5ZDm9P8yFVtRmHubLAXi3se8eSWk+ny6aArepimf
OjsbluaRbowkWqv/xrP+Ozsrr7Sn1zDKQcdokUpKkG+3i/LR0V5AHFzihs93F3h9uVHJoT0JAilo
dlcjMvGqu7u8BrB7yYtw2CkExK4lWFnaM8wX75UnB7ITOGhgH+B1+NS6IjrA/XpjIs10jOn4IgM3
Pet3SDzEePsUDCOhpdSEoFh8ZzCmv9xJO62Po6Jqu5gov+CNwJuA1/AFuSSkiTDo8hEvybOIVI1s
tB2fpbo5GR3BaekbZVI5HmujdZLHNkvhRKpySEBEztj1TmEFS3s0tdvYbCVwAk2B9b7VgMpQrxiC
9YNhLSXXef38B7Wg+ICMOYaLikbveOnp3m8g4YrI5LiE4AWB0KCGuxdYLkID+Fr3dODuwWj3lPw0
f9kZQ5+gcdqPkxljG68ds2oJscO1k/PZhb0Gfap1OC79KamqDudmeWkggihascxEJu/Xisc4BP0Q
8FTIkIWPL4dLwbuuHFjRaxG0pLMrtBAZhA5i2VfzxmQSPSZm7y7fpSG7ITb7vOReg80574ySVdEu
90nQIFt8nNHb9q+BvZnFYCDYVVWeB0AywNZUhkOUOyfzb+cADrTXmRl0Bv/FFT5Y0dZtRbkfqwgX
PkdZBJVPwflvn1+Z1+WBw2qrtBEcjgAaLq4AGHbnJlnppNxuSsFRbrNUuE3SgRiFYSTfHVvgU4yz
fr3JgvxNBtkzwyFDRzNTjzIWRrr3jTXRQzo3WvRhJzDwsLSPvY10ZCnWT5Yz6AD0mX4fxrrJDk6j
pjUblcYO0WziUh0Z/ISHflT6DO07bhzPGpZQ/ht8ciVqWva8wu5qyHV01PPpr2qtJNI9kB45tBbi
dNaPrDx0ykADu9D+pz+zgoxBK/Uat7aRchRXyfkbZJTVRbln9cpU0e89VLgWBOLhffT3o3P2zlxr
djsXVYeAWnBT4dIGYVQao4Fqz9U980iN1gxy6taQWWDFXUy8grIKFBAW98/PH69abDTUUAQ46z1f
CKEcxkWmb5E8jT5WplDo9gH1oRgdYVpIbRiizbPJvhfUHL6tE5J+uIN7WMr/JK/S2sMOBvec9AtI
6IG8/p9EpyNQk3RPUHHvmJoWWnB0MCZnF0simWdSn/XGZE3X8GfdmmK/l+m7NoRnxpBZFHRVS2ka
8cNKfNQ5OM3Z7cqkrpTIdZpITNX5ljzIOCPaa8JIul7bou3kS/EDqSSkbpHiOJDtWFLQU/qhJsBM
IiJMBjGJZacZqJElsuedPeShNkMCbUuN8WiVwwUrkw5j8T8zTFntvdvO9589vnqdTKUzcnEIEDwQ
HX0L7adNo9ySvp+LmDq92AH5HU0mec3doArxmpU91Io91Y3Aq39LSi5TZE/9PjGHpkNK4Y18PYSl
fj4oIvYNWVYp554onBbXN80rIF2CxMiIYZ7yUgjaCoOp9d+aFi2t/92H7SmooRUxX3P1SHNaz33x
8gGg0D9rX4y9AUJcPGYF7OmXHDS5M2TzyHRHvUhPmTChJ3SzCsLlmaU7tAjWGWQU/axDNs+ZMhVs
dOc4pAFU2GHZAe/O06UySEW90gJU1Qfs4p3M4xkWzCLc/zT0F4SzfTG8h9F6nrlBNkHV7heXYAIi
gO1AgREbAlRXYbpWkc/WU0APZ4pDbDK9iDUy4YT6JbRot3hrXvyu6hQl00u7wMQ079UAEtZl5qK4
7XAo0GSG0ilshwx62LYSQBSzjO8iJWIUkwLLXEbgjwlwxUXUEjrZi1+pM2pIXIhOJkVm645hP5tg
tSpxw1hWivPweSjrp5tHmviYPEFKsQFYjv0neWcXcNekRwxO6Zh/OILWr9HwBK5c922oquc3NiAe
zX6Mdh9Ly2FZ2LQw/LNmFnPm1KhTBGeDLHW8zshGSyDSNMRyEdliNEjGpqPGvYOVcOKa4cJeri/z
8MXW3Op8ZpPe9fFV3RMamx5RbMgS3eIZS+rKzgYQCRDEoLPq9Llm90yrUXscP67Il5Q3SFroIBj8
+2FJJ5Jg7HK/HZ4lmkC5kfAD1XCvvdpoSf5dqN9qT9lyxHkkvo/k25G3zJomLJHRays4G6EHEHjT
oMZMcqGvNM55jVuHpE44biiXn4FFPsNd6FB71Wfzpzc5R0w81B99is5PDVY1LN/StOcv805X13dE
0wh1KEQ1S3/OzFi70hp9SZ1+yLKpN/0pBdVwmpmrxAgnvQ1TtWDFAwv497siAXB7VmkPcu1+7jkv
GwK7sELKSoJlbDI9wAT7Wjq0inF2+lLEnBlv2eujEvZlHVwi0KEZGe01mLztWXS0YA8xCatgdkse
mjuTrqmpCl5VUatiPBtm+1wKUncoZXh9Miqm6g73VwO67vy9X9ePqTYvz1yzkrDwZ6dH1Lne/ERD
q8Bs+wiCNzNnTOFKxDNrs1x357srh3ZsPsX6fGw0upIw05ETEoMNGbxBvKViqLGTTd7hlrNA+GYC
YFmk3FkFVUxgNUxXE28brb8q7yOes5u3+ViUzBNvecPAJwA2T0fKgDzw/XqWuuWiTB2VNBzOcPUF
yHQAb5glrRihAwF1J/elNTV49gP2hV6HFYIAyDJCI600oAoT3O8kvarEmZhMRALqY20WL3lM+EzT
4g8wZIPWiUKE4CZY6penGdtbKQIdFdCJBIWGohNyQdNVaj/4m0O22r1dCDiDolgzFlF2cbBKcyNk
G89vEpj7jdkC22dBodpW7fgkugfPmigwnvV/VNgGh/08gmVEMgYpadc6MCpsgrZNTHKTOMP4WrGw
UEg+xpZh8zqXslkuvaLGuAD4+vI3BopW/QkpD2t1FCZrg1EDupLYBI1Bh7s4FJgCiY2ePlOR6XIW
mz4taj1Jln2DxAEf+IsrhpuE7e3oiGSqUXD5hA0aiPG+8XVu1A5o/W1/LQXskxzaKAPC9i2nGCVI
Co1QztLr+i0r4Dk+u7/keL9835FePs0phIQAa+MTwISu/1YI099PqcQ1JigHhMHT8PwETkcw7RS0
i7FXAXbhC+7Od9vIcmem/Z6bErWNAOFmQ7Oh+qkRpQo6qTFqBNepq7JySbI3KLR0gcL0uW1cWtDn
SEwGDMuzXUQgFSX+7mhGYX6RCIhpBeuEvy45cZ5Xz4G9B2GyA2TpvrYgmT++5Bx92/rIk4lmDbbg
rYCvDNxGQ4p7gNKOWsJvXFj9YCCf7ryIf1sOzqt6Pl1sbAm5CSqDV4ki9Y4CqBLgfaO8mElwm5DI
qEaCoKOArwhs086XmFYk67iekw9IojAA9yzhGrgL4kKJ+Q9hOhSDY0v1pBigQSyZdovCSxbysvzj
NIDd9B7FdKzpVeLXLpvl2NztaHGJdFuVd1PvSx4dV7lXQrGi9Pi9xp/wJbfDaz/rtXrLWGNGQs1p
E82KG/oPVMxV01oWNSBo6bJQu/XzN9wyZAwJkCvTI1p8fqX4HaC7vkXE/LbCW1KaMrh8bNU9K0EI
OrmOBckxCbwgwQkt/dM+534kXzH7RbZS2X1ReS9UhNhJLdkoKKYsGSzEjkpyeGqrW+yPYn2V2mda
NPl2GGb1GsnT7exQaB8VyQ9sQCu72yHqfq1/0iKPcVsbyXPT+WcVJxyiLTmJkysywNH70U+4yEO8
Ncb5knyYZ6qNaFqkdj7b3QsBUOQxOqW2kL3VoNYlLdPZtn2ZI3XlW4KRkr9t0f7oEAD5Hv89l0Ow
UzAP6QBNWMrlYIUMr61UdZEJY74Eg8ho+2aKam2O4ciwNY8+6PjssLFcVLnmVcR4JbVxicK4hM1S
jeJyna14WGRycFI/vUaWZ1hdtgvzomTbUrnBhxjeTOrp/gHPkgb4oaxlRvhpNq6WbSy/CfiLkdzS
iYrwtjbAuFCx76ppmy7PLIVLzQxOZmx8tQ5VvSt8d9vN25/g+/ley+ffGqVQcp7WpzruE00LiNFC
A41ix4fF+IR6RY0BXPiiMzCervDGW8QvKkrH+9sIf9OHDbz/CMi//CnQ3S9ShMjfSJ/yyBHa+/h7
xEiMddmw5rIi1yndHuWhQ2hdSZ6gKWQmDpAHWP/HS9ekOajDaodNlhJ7FrylAh89oB8jesAHmuwm
Z3l4cMjwMYtViEtcXbZgbLqT2Fi5AAZ+WF4+SlZdYV11g4gqh9/bOQYMqI8/5YDl7cl7bv/hvYrv
zFDiiAeinwRXlq8XwklTk8hrUH+v9aSsdQbhtz2QdJG+KqLMB4vqhGtlfcS2aiVgEx+fze6jxnhx
SGZduV/h2j0ODjcFpZIP9EbnBP/omHPrfDpll5OqA6hz/l88Wca7NG04c6dd3UPGRS0lqLAp7AtG
0CCINks4QzYiDP6DQjkHAkHKmjoN5tAfaHN5tVTI4Lcj/SKQXNBgx8Wfa7S8poAfhpI48AyvNdC9
09d7gNBcOsmsNahN1rD/jIJWLjLIOTrm1QwWMSXeLN9GUtJXe3I0n7KyW3dpFL7zMOf0qTdDCts4
RyBCrZozQKj/V5jLRGmFkyOdEVQmiyrnsawQeC6Wzoguj4iIntm5Pp4T/GM33cBp6uiK7vz5+ZGz
6AQjcYYKiMJ7/bLf9ZmAhubm7TMFKND9g05XPE1Gn8zy9nAS5QJZhdQs0YPHuMGngS5NEgkfjJMG
nJ6tyAhPYvB/TJ2G67x1Z3ien6WKCVJg2++xMQnCrTFFOBrES6NPAq4dV4mFBO24Ics/zHQDsFhs
GnpIiannRAEAegDsBYBkX5gzQ4LxL/0PD2ttzbMdO/kwRF4q0nkTvTGxd/AOB8Sy4r16RZ5TazR5
LpPEYmJjGpk8E6P+cA1MGl/4Xfxp9esfDDibWyTdagQJ1CmhVsC/AeUrJjnMDBcqh5jlRC8y6Fmh
690mnDdatzZwVbBnLkGbTwwlxnPkhPZtjFVLplkpGev2WTtWlQ3N7n8C9HY9Gk2kIlAqUwsnm0EV
W5z54Lik6jzEf6jzVrrZBa06phGn3wcoEcD56w8BU7pdSEqq9Y2HVHLEgLWQR/pYpju7oNhNituA
Fgz1rU2ZzFshRQ9AHQtT1AthEZ+XxtraEm86phy4IpbiVKKE6ku3Ye2OT8d1bUXVSvMgkmuz41ao
QlvbGoNT9YMWnKCpV3eIeDzCYTKOOEZK8k1/sKoGyxUzT48nV4Xhp1H56uia01Auo7OSClTkGpvL
tUixUjmJuUVezO9+Ymlz8Enebsc2KOKS8kw5iacLXKIGDEdlQubGwMs93+mgV2IdhN43v6ow6eWD
+P2OHeBZlmapIiWhBkRGwNqgwIyrJ2jrNLwlkl64/EkEmkm1WvXedMkFcwF8Pl227BcbVhEzQCSx
nGQZmXAq1i3p4Ixp1ykKMSj4NLpaChKx4a2bm8Lwx4vKMrrlCbG8L5vBSQ28gzQ0pOK8Y89t+nIh
X0uxw9+i8HyrgWFWkKUwUC49m8GFYg+qt/YBXfpu+wBdo4yPDxTpC4P2lmyjgayfilvtU/dClPzo
XAPShnLdqLyyMJFmdyjbJYikqV7/kL/+bh767ZB0i7mTS83EcN6ftVQcR9Xhd7i/IT2LHoKxfWJN
ThcLQFc0jeZqE6EZSZ1+RLdnlgbxLrdDu17dBcoZuEMvqApD/f4kKz1ntpoW1BDZBuTlrp35pEEv
l2K0AVkLVeaf/hNU2dE1XnsEsWeWomzNZ2N8KccsRLqA5qbequY9EX6kHNgMj0xHyo6QLLCtjymM
gVbM64jtsF0+75CNJQCdGKELmzmYb6Gb/Ip/ys1BiE3HfThkIYssLNW3dr32/RW7AWh9D9Dt3V+W
rONLcWgc4FXJBq7ogl1cTlfPsnTU6o4ounvDKF4onzwtxxFrsT20YAyxP/7w7LNrve0G49qhe2er
dxdJ71mgoJl8gMt9jbPc/rClC1WxT8frolv3QMe45mL64Hqw8PhuiAIYym/oOq9cZ840iOF/b2As
tsLL9I0tGPNYDoZVnrpePMRewl3wGS1Deohx59idFOrTqz3XzMm4Zkh2saYec4otN+uiwPoNYyZf
AOAwwDxykBUdWg76ta4gT+lCyS5HGnbRNqwJnbDWZQOeCRYT58lIW0tcZn8d6eGIj/rAbw9wv+7Q
Ny0ukgM2UJuz9K7bQ6Ey9YBWGxJuw2VHItE1jf29jVGCj1hPodu0dV0H9mW0iit9A5da6k6fMzT0
yZmAKCXKo3lm44NHGFSDiiPtB36twkEToMP8Qfha/7WfyBXJcs/JjQ0mncrtEpMpHOELSfZJ2NRZ
j6rzTXSebBT6GukBxq8AklqAONgIiWN3QKLKcEgb0b/r+pnxwMjSaH4rxnsxgyw2IQi5HgsJOQTW
gmVWHfErKwrg5qQS0qMPcKwm/hkPctn7Pv1VYqSOb+GYnvAkxKKG3sl8Wdj4ojJf/hQoxNsTQWZg
NUMIoawUKZXWg4hhGSVtnR2NpoG36fxIVRbACMDONiyIAnTniZmDOZrJb0iiwDP1aS4SJx5gvT9M
sqPQKebNRPosUum3OJxC8BqpSsuYji4b5A6DjpOgpMQsqBNUVW5Rzm8304g+BkOhjUhftLDSTl6W
zNFnqh9NRxmK3Kda1ZCwzmpfJTpAwK9SokQBYk7SptQ7oVVzIly/yZr7iQNaOjukZ/d054Vl5jgJ
PCw33pR1Ih055rj7LWhK9fZXKphtmhqPYgnjuITL9PO91RTmLmIoSFR2TihrjdqZRYYUAjUl7RQg
+d2U6uD29yBY6xlkc4HMkvi39kdrqIwzP2lGkU+SwxMKYfThOl7/EWCo5f4+bB9v/d4nY2nIyq9D
Y8no6/sl47WtFnHg2FvVHppD+8DeHhFo5Z3Q+dLdNOYe4S5hjNLS+4V+V3iMm/to8lMuK7zL32GS
AXm4Q80GwEGlWD8pCE/eki325V07ALi3rGQ8LpIpOnRLHOwzUAXLap+kp86ZgpAIpOM2IWgkmi5m
T9HDdoYN/VwUovj+qC7Vga9XHi3wPI5WBzKooXFErOYflrzsY5gSWqeE2dLlJpa+8/dnNDXtn55e
5ZHKRVMRx2GLDMCJjoSioIGvqYuGTTlP0DgaIvW3tgrtQqw2Tin4JqCyIKOFQkgMt8xO3w4YlXfn
TI6wtaRtHKPOQsV2yJJIxgFURCiDLwZ3AHVZyG9JMaKqV4tww/gh83aWCgyNCmB5ThiG3FWQNWSB
SCNW3vQ3/J7WS9g0npXqiuSlNLjLTN+2lAQK48WtRDWogdUhqgd2hjcUVDCN/UF0KxAmVJ/5bxzQ
L0txTUmpUD/8RBtv9KErCKyvY3DtK6U/MuWYDrybb6fqseOBuaiR9nLdzg+4LF2iI8yTl+b1Hi5J
mUBGgEjWXq5UNKFRbQYpfV5zRHW1iiDnXiQoGVE264OG8/Taj7qSJkJossdDQ+c88gRP7VBzDHUz
nRQdviqKqNchnPV1o2X7dS7NcGZXwEkQpcDEUixNpSQ4XyDyPGKLErM5RIboN+vKJhGiuHgAMpoH
etARPXX5yHuF4s4pVwZyCn7CrcJi+RSZCSatzA2WegLHWD6GhoPbW0hsJti3UzEsp8BpYSp9VkQP
a50SZ//GbKbllhd1cfk3PiXLNh289HY/73o7wMn5B8YzdE+plLmMxCr07g132kMYazB7ggTZqgLK
0rWTI4ui9IlctOiXMUTZ/45ax529Swl6kdooT32w9SsL2ENL/dEYlScpoaHkySJhbuF3oUbyrgSm
C35NbdO/vGo7iOsmxc4QpcUYFTnRhsfdjvQxU6WEwo5VaNWUHsnnIVTJbJ7LTfHaCg6Xxl73EPWI
vV2C5m1J0I/x7oRd5ARfZ/jD1NvULejKJ2r9KmF3kBi9/s1cqDcqa8G/5mM65mxPVNPbCtX/P6IF
Gffxec/6bJlVNhwGme9KsIy4Di7gdSE7EOTsOrPfVhBig9enUAM6eDBW+Gm3QeFNZ9JQdwc0JLz4
NrEvmbTaguSafy3mFu7rR0xQsbQ3bzTjw/Rwosq88IMbZkRnu1exziiNkUBX9gpsgZeOQhVk6c5d
kj00CUYDyVBaw2nBexcUiFkxmbkzPPX9g3FpPA+Rv4TE19pGUdZyyXSbKXhbvC1s2/fC646ODUSJ
0B3bPDEhOpCIdCoJW7JL3pYsHYYMUOv5y/oSAGwZuX2+M0wTOkBY9azNoD5tPE9Ub71H69WT49i5
gvZuL2vFG8kAm5m8Pci7jFFdwoqqQZg1o5JOGLrQ3RP/6/Iju9M59/hIRvK4wn3CKK3RuEs/r78D
o/uwuVkSV+Anek9Sdusp+eB0pouR3onLpfhmSrV16VixaM+Huz2J416/buEXGiFx9Vor3ckI/vX2
GAHiR8plBzjn0QzpIYcSHsrRuptYxgI5Wq3wVMc7IZKK15JPaZ8Sb3PcY2+UxkHqWl6zORr/nDyb
BugVLk4WG9VGAqJ2kUQ4qxl+Z3od73ytMSfyPq9XuOzoU2ncdw/Wf/e8r8qptYJHwy1gEQ7E2/Dx
lXy2ltPowtKLNYx1VyVMntFzCvkpiG+PVQWLzEbM2CtH1lsNJebk1L9E/1itSqAZljlF9zbEZQcU
nEHumUP9mSTZOht6YBJg4L5RXuLQKJmnYU7eveqfWcC0Iy/X4b66KhwHUMAPSwALGuX3qTC4A4lD
52hoIhS34sq3D9T9CKRi1v9bsFoIBJnQ0CrdfzaOixU6cU1T4J8vcoAzrLYt7P/lGhQt9t1pvIiF
rzDifDRBu1FQeaLxLlMwG1N3F8L1SbWIK5rc9dPtxhZDCMsWcvMKWJ9g9yJqxkrgJ1qAoe5v35ot
wdfqATkd0OhR6k1vN2OFhau6Nomj/YNRlafGbU7hSf8rwd6x1So/MdZTGNkHpQJ3107fDXOHPvrh
BTB40fkOIgytll7bHWdty+6Cmh1GBWJV5DkPSIAcWs4qnvksvZ8tnSpAdIsfw2jheL9NaYv+SDdt
NIdLXGFegJJSJH/jKcGAuLmbFkyu21F+9k/8caerCsR0ECcWLcEvZIlShxFp0NSfbQqKKwpc9N0S
j/n0nXgomP972wLOCsZ7on0U5qmBAmFIP+u073OpSJxR3cdTDSvUjuA0u3jezg3Y5fIPOaGWoKq+
xQaKqB850VJZyYwIT9xjL5jJsm3z+/t/7LJ9HGEVSaSmr2XQSROXXzUWscaSU9Zoxnb7zECKoM8Y
1VwE7wlOKprAaA7ToHofEGM1zELoQ2Zjug5q63LT0fnLlhNaPHjI3cwOYL+0WQnQpgGbD8/0v5lZ
Y6zNZDSxUy7uxcv7IMZaYtmoyULIY0RGZHo0h3gD9H1jFxaWPI3JHIaODbaP+YyuEc8h4/KIp4hN
9AQ1lScrQKnuryBJqL9Qmt/7unQRLMiI5+L0J1L+xko3ZR+Dz1xtHBQwqLffAnQTD/Ya5aoaSlo7
UsSNRNdwn5biMOF/xIMJ8sV59CXL0OS47Brn7PmL63YUYvxNl8A+2f7xw+0j0RyUo7HztZigzz0k
PqgmKzOsK+cEecRSeQsGUNf0wGPed6lo9MJmDgtS5XCtlPydCe9TeGa+aE/1a4JVpjxhT1GZw02x
0VC30Nw+4S9lPep22BudxoRBh05fIYLwLPHNTeGK5W3gzQroaTCsQu7s6vJnAWcMNroyVjvJ2xEn
4LS/D4mBsjRa/bs4lrXm6FznlSohBEwH3Bps5eSrRjkepyG/VMFKkE8IdQPJo6Ti4g0Xpbkm4Fhv
OT7SHsXI4HsR+GGAbdK33yjrqt44+x+Zbw7vrKdYCVOMpbFgelgA35iJHnsD2Qpkhe+jGoKdpAAS
qKw/iEwbtJrsaXXuQUpaoiY6xZQHsYDPBiTW3f1Y9z0sd7ZYNP7xHgaL9b/7kcgXue3pCX7O2CsX
VZEOvozfiOqrWwcekjjuZX4NhazM6AlQqslPqP2vhN0igCTPPHp4KWGhn5JUZIkLyU68Zd3MIa5A
EZ/BOVJz5YcAnn2WSb6/2kbowvA6uzMyzdg3bI7ZjVP/a8FbfTGqd8cky8BAfytsTjuj8K5XAKnI
1Tt6F2sqLPjM5d+XfidgwRGzhRLpiN24yp3MeXe6X4yBbmkV9IxMFmaEJ228pPjvto27bxH6bPhR
wqM7oS1cNyMulIyb4J4reYZx2rLDXD21YDPpcXBgSV1O+jUR5z1Sv1xezX+2UNTQfUQ86hMvgN/7
/p9+AWsMGkvLEIgiFgfE1F3emfJuUCpxK4vXWueTvXmH5JyydrOj3OITGvIidqoTDWu6uEC1IkKQ
PMA++rxhf1qROklzmNySHpnUN1tNfKS6/tdSRBox8gREwG6L9hfgqyACtX6DBzABP74z4VwpwSm0
MJ4u84hqTpBNXstGN5rdelNZwsTyYUeSW2n+wTetoJYSZlrOsMjvXM7zm3EDwuyjZTNEMRb12xgr
vreVOGkw9HbRLtyGIF8ZwXm61YzEkBK0Bu5FmnsA8Lduo1+OBbfpByXc31C2/00VL3XqPrC1IQIg
dqMcVulZwrRXGEo0AHvEXvgFMEq1Z5bkGoLeyDNfufZ+a3J4vubnUXHyBbEvb7hHDtwdTTM0FC8b
fMNK8/InLD3CKok1PIJwuO63eflSgAaOtYTOMhixWY2w8n2WFFxT5u0Hkjrz+eXG1DKNX+9oWtDp
kU8rcDriDNGmKYwwl7CB0UyBAOPJB0N0TiinXvJ5GgC6mKKqt2OBLVCZJSLljkZSFKtKhAQkQJKG
T+h2d7HseESB6mlXnB6iN0nRTLajefRz+m213Ovu0nxJz2JaIGyegk6T/1llui6nA36eTsS/CeEj
+aNGaeU37XL0BgfDqdUyDHhZoREDNJEMbCmLP7jozs76dTY1FZPrdIpkIJn9wmEdSYTUeS8cuXuF
hpuUq4/RPEZ/a0HsfzMgN1B42EZqwjMhPafLyEYzu2u+40KAOd6UF1N0Fz5vNouP0jYhbGl8C8rP
vghglEaMYhBvDuCmDVsmdjsBLnSHtJpU/ngvkxfVLaj0p3qVycLSb9k3kWlh5Ow5s1lZ4DK3aT82
FNdCU/7nExzexjR+xGbESDVbHgjAT9eyGoxAgMIcF8wMnwi+fvEGpi8f+Mfle8mYM7wfb/+BVx5Z
QiEG+QynF2C5wyk8P2JkRsIAJG/awQs9eJ7KO8AMHnWpBa1tRnoyjd4xvf9lOXFq6l5f2+yMg8/9
kYTMLsKyMx/MOpv/VKr7wbv0/b8vrOjQPsmqzHctxFMPn1MV/PTkGoDiMSAVtAySLEi7PgZ9koJz
houwPmKMCPC/xhVDGWfkTDJaBpI1GZG620eOVmOR8suZNwYWBTU7C3I0kYCPcMgnwLShKtrb7RPb
NsVtzfQRfm+8j9raa8hZU/zbeKgFEEbmaVdB8exbJm2KoDqY5kpQgs+EEXdInMy0w0S1qNKV2qfY
gIB1JqTljTtY3z1xJVxhVzzX80satRMMKmaN/XnkDwYORH4qkmDhHg0tdG9Ggvsqk58Jca9oon3k
CELIGaDk5J00fb1pGzsGnX6SW56662Ry3ivf3irw+rxi0IcMBfPuoPwvQlB+QcDy6+/ISCYoOXtS
tSSQiByxLSz9uYxyn0QKJuDgHrAgX7v4aSX5awU3e25jg2fQBlHzMT0r1ei2ZXVSuBvbGd6g4Vd/
qF6OONI0hfn29SsJcRwAI+H5zfki1/BzlHstggQsiYSEpqgKzIQy3f2owjFhDf3Y0iRet0mFRXXL
Se0IvdLLUvUyG+73l8NmbmbIZCnGEandZ+mOQD6bgRm3Sqa45xt2wefsFKAquvvI0413Atk9OYkw
Zcyswy2SMZ2c3Er/Blfaab29kWOF+DtmM0fMn9IjnNHy6L8o2SN2YpbrFGblxXutF2AmaFjLY06R
kt07trl6aMQls5cOZVebaEDqifpg8nr5kAPR5EoIi4JFwrQclOmSqP/ny8FqiAJEB1V29CsAcf1y
LTu5VXm03pB/nwXBP6WgonBN3STIUThjEDrYQYTBOdLwaaarDghcvb1UtruHEPfee8gNQygZFs+k
ct0xtg6tWWzTEnICAaEZkHBH45UaiG/X4frlihGMhNPrXIPAW1/NuBgW45oJuAdPwx6fG3IWQ54O
fDBqO+oyVynW9lBs9i9Jo8Vy0dVOyHQGdWc7L2B9BwDMAqSYu5i05gds/uIlW30gPKj2orxjTQt0
WrCeYHKkvtFFu80n/M9TE1gppMv+u6ybtmwyyVWwaUl5CO36xKTGPAFsyzHTz5SgNL/BGabwdJzE
3jOjJ0emJHcf4kCW6OZMBRl0WCIP2Mm8LtoEuIReMu6+NpLSHRCgkAB3hFD6Rq8w+Bz9pglID3ok
CR5D8LZWU09O2n9S08+2RixhS/DQRfqzN2qNxjyoku6hWtg+R/X/W1uJF+Z1VX9L8QKf4r5KX82c
5Y5RpEQ9RwNgZRWVR3ft83UF0seGcQQ2CVfimMXupfDffz0XgNNgDNUT7EPkZ1Re9NhBfclg2Pp2
qz8PWWzxm7YAHhhpbyhm93ARL8tyt5dNCnzdqdKMcui6i1XEFUMphMBpUG5wZnD9gMPiDxLiI8Mb
5C6kuG+T7rNcOiSa8uIOFdXOoJnNa84Yvv2pO08XiMH5b4Ir0bcrslhykD8idZTRblRtsACz+Kne
rf0PPPXOH1pKBiOeD9BReyhKPV0GhDRy9QpUIjWR5wxkwOnQ1yMRQ/Yn5D+6FJI2KuXTsPcvIysg
AAxAFQZmPgvZx/TKE3uzqQNSHXHb2/r281rl7QUTKzkkwwqFQ0rl9TV7NL5N0+PxD/6gChTOD3SC
dIzWWTXbTulhF/lhFQYBE2sahpJf8npoqWlYqWu08vXmjkFLwibrKupFlhpnjj2yeon2qb56f/I2
PotTLJQGEUCBXTEka9e2FfQPJHZ3KKibtgmSIbIGAAcuhyrKTsEakp2Qnhxibhv7kcW9s6Nq3Pby
VJVPk/rJh+iHskdzQVlMwOwLrJT8/Vz0Ur22wN6NB4AWV5DCaD8de38zoCtyXsjMnEwPXdNJRqOX
e1By85lpeIKSgWc0uAyf5AVRefD/KqZiklwG6hczDfI4zmma0QQQVOtWna+JDfDKmIG5y7f7f1PG
Z+vQrHTS92HZ5wvlHG2MP/8hCzcleQjd3dS5J+KvIny+tz8TwRlPDEn/JMWD/7uXWxACOaDJ903W
AdOqPvdJUaLHoi10V9uVFNeeX3Sjjwqkic0t09fJnfES77B6+ALaIBKE8HfoX8OBL3XZlDhEuJ7u
YtE2Ckgn9YVKLJrS1Pt3690YuDknAh9ZUNsSfrNQVAMiQdhrdi9B7Xe2gjBAc9e1WqtdQB9LJCSj
P1Zjhz8TmIBlyyxor3wVvCpS1C6C/DOqJEj2qXGqS2nOzRxqjwT4B8nlkVX+W3zioy8/HSCi5URa
nrM2JJ8O5oKP1XOb9bXCwmaOXlpvMMEOX/36NrYPMMglwHfubC7AAxWqqaQqWNR6n5kce6EdkJNX
6UEZX2WOn5TFJAaI5ccQwNaTNy5iShowpIePOOX+92nUyl16iAYiz1ve4THYrj3gFobP2r0bT5k7
OQXzTPHxj+DyrOdvHvBGtBjBN0aUv4g3k6cK8wnmqALVtTZe5/8e4gJHC7rizy1bwffSKyt05i5A
hrUCRiCd2PtjgwzLN4kSqx/pfR9zEC3xx3r1DnUrnA85ih5C3DTdonC6hNF+m88UeFgaMOUSChEb
EEzzgITljftNa/AfcbffwipDoWK3N/LV77ecXXLY7Slg6tMPD7YQHENPYRb8hCe1P4EunKjsN1C/
Hn7wXMsJcj0O6R7Tdqqqri5Bf9qZp+nIMWagRBYwWRwZDFDrVfVC4/uaR3y+qO1dNDTzbuUyoQD5
1kBw9XXs6Od0A4RriPIk4wzBBmRukm3q2e20Zr/MlbINLhy072v8r+KVwKg/5YNxE8cxEsrjJuVB
YK1rcLcBouJD4HHIxf9ZZlir8Z9V2rx4MhJSHq4uW6I+Y+WChALB7rk6i5BXzggUqZoIChF6zjtc
uV+lIo6m8JqmWLnv1KV0V8MPzhMRqKP+a8c3vwAGAVkdch28nUonzzcPUTG1LrwYhwfqp58XOyEB
/xfZT4jDuiOpX143LpQay0oA1vwvRajeJX0VUId6qunVy3jM8we3wWSWBXEnqowx0wwV3uoUXN8l
MALgI8SgX08R36Y7eh9H71TGHInc8Vux/yfvCZXWuMLfiq/5IuZ65NqOHZ6fMyy3A4O2ezJ/XRLq
fGCwOLvhljGEq0ZzMHGW9cUoTBlG9KejxJfdD4iqLAtXLZo4Ah1+bqT87iD9UVGtqme80Dvyx6nA
NQ/nIhhb/wWpCLDtFWX6MF24flgFqAwhg8cADFj6f+mu5tUvyfOkKKx8SIEim6PxrjAwZfo+mtWU
T200DvjPMJ7pUmxUG4HSX2wcia38m2R/kaHEqZUmROYwL7p4hqjE44SIa3SyXlX6XU4eJkHbLuju
tvmoExgB1MxNVJ3h8M0wJVp5YwiuM1ROzQVj99jJeihxQvVUK6cM2q0CnweKikceG8oUaHYrkEzP
gKfTfjKEpw7KYFezv4+F+K7AXSk6ddvpcOhgZlEXJbCkMUf+1gLpF2Ix4o5tt6MXHourOhQOSjlE
mYmjaJEDu1X53fKiWXwLSHdLZ+hapghUDfnoq0H+5k34+rrHGwwjWaDxZDq32w59HeVyfE4gEqim
P/ysLh0IUJ5g9fV7yTXgXE81wGPXW5vkqGAnSNEjq51J2FNe+5ueANlIBUMVamRWJYKuPEEQ2F/u
NQNzDRq8/Nrt0sDbY3OWHpTxDNtVPuoo5BXwRXk/WsXMxxiTeVASUfbwdhd5aaBdz5OUyeycY5FQ
gR2ylH83bYhEclCseIDnIRyOLh3sJ5sp2ICL/DWv3CxLjB6Q9ck1RWtb5oL8v18ZEHIMQUqbMVGs
hzFWKHtVNKNdZ1NDBSZ+wvBSGbHwZFqng+FxEdZWIG+myD+p9O+Kp8Blg5NfIR5TEKpCR3tmUIye
YRJ/pZD6iAGZA2MgbeLQ/Asjl0jlvtg85oQ+YMjgq4wBB4Yg/d7n30z8+jx/y/etzQT/+nIc6nNH
6CzxXWfFNpVOun2q+GztXkhEO+GsypMiyDAvpcWbGKpvxF98b4UGUs0nyq7DFPTcUydIrC84/kz7
0OWvai9YTeyy27PeiAasDUfjGD+CciIBuT0Zr5aymSvMhdxbjuBRuKgghlTPBcvcZfEc/WcEq+St
6oG3LLRqz0rwHvVzQtJyOAl/xuJOBcJzonXY7TXgvPYlM7eESLdESYuAcxSsbYOn6D4GxrWbaHkp
vnRKK27G/gSPVJsjtOpE8faKbekUWuGqan036593bCOXU7/jJjyDiALWzesmkxes3xcASJgI88US
U1tkAnXUkdC/FckwW+VujAexErwWp8gl7wVx6z5A11R/FrA31bpOof8PzLOmzKo5UyVeHfIvO9E3
VYIIKeJ/dtk9HOCpnJVMAChls/vJ0u9PJEFduNYKlCzb4FWgK006lBMZfPHQP+L3AiZxAIE94OeZ
cg6rZ3Lql2I43eYcRZrvXJC6xZPBN9L1s/hQoGsVyHUm+Lu6ougyh/5c7uJjK6PLchaVyGyXVObX
nal8SKJl/lP3v7UQdg7SL28l9DGmbCgvq6SOBlETPwWsNx3HnQ0AfA/HOhXgwIXOr7WApYjx8lVT
ZjW+SFmXW65Tu7JQZu92vXcFHb9oDDi6BzTjXk11anNuCvWhLf+DmWMoCckyKkAz+FQg3kxcrO0t
t4tTQumTyUjCpFSomE90mnAxnzVZ3DRcQWrfGyeg26QP9Z/hqnUOhXjBnh44np+Rp1bOCOslyyGu
8RUgdCnacn9O02kFZM8zQDAH/l1GWE1nvFp2RW/kii+Bgk93rhUHP7Hb9m+IFZhTh7YpGYKTdDL7
I6+OoLj2KLeiF9FAT9eC7HRrD2D0k7MCKc2NnUPhHeo1tQqICY4n2cL/tUsPR9vlhdNgNhqF1GEa
OQSXvg305r2u4G7VWjvHzxk+00q35aeB6szgjz2mY9DVj2CZBzm3sIm0EDVBvdyOopItVIipWG3H
4aCmFEsEUODL1XHtuJZazY4ILtGIzVZuafPf6Z4VJ2ClWvFSCdrnAj9N0PGfIRBNrbEqpmIunq/r
zAc08JTSf1CnUbUsFy95XlfueD1nhbBxgPxUtOM1iZrgsY0m3qclXbCP9W8gf0AUHZipCGDO6nSt
+sDIDXbqTK+t6eeWjo3obonGv7SQFllEvw6GN+lwJ+8XJTynPami5bMk16UULhzKM8inibDwfBJh
NYUTOvuwuXL1W6r1xiBVAsn5yrjMhZf5gFgbwIALSYkmfec9+z0CLPfnVzhnOlU24798QooMX903
AKpsec8mUt4rImoUpTrw9lZBEbBYpXN3UHhhQlsJrP90oQolHDq983qoq/T08NXSMyYLWB09o6ix
cnIVT5o3dImM/7PklXEiusySvqdjOjZAQbViaw4Rczd1KCvamBSjUa2TOOreGrMLpt48ng98j7nI
MddQwkVWSlpUVPSOrtpvPEgU5zQGXeCL654D4zcpUAAf6mtwEzZQB3E1Y6ffB/s1Xj5AoYwbfkiG
nmiOY/WxsJEisOSErOQrtPS+C5I0lT6xlExI95JBpPPpkBWzowE/MLilYuthHPua2LFZhL1A66CA
ZG+AfaopyKbMRc1wcpjihVXO+A+UVgAvpXwZdKsP7wxWXO8B7qViWa2wUwc88G+AP8TOr6GVU8wv
zlvtTWUFwmd7U0D789tW1frj0Be+Kh5P0uQtdwDtc96H1G61mbt3tf3RW34XBRZZdYw9ksb14+Jd
fQ0zWssGAtwuGsitJrKXySaEsHXYWw0HxErzn6BRkxaFrpsSOqWwP+rI/fTCta6Q5MqD9Ep5Cu69
6qpSYdgW9eF+2Lmi0y3c3tGblkKhHKb/W1kK/cZTEnIPd6E51qZtmZP8+zY75T9tGqzrh9FXCm8a
532ip1vyhdWmZiIcJfeXE0RewOkk3iiy1Sjxgae/EGxeffGftEEUbEgA//1IQEe+lw5xVx9SSCQ+
jR2mqMdMa3Upoop3jyVju1ITQ14J8D2qLSYlpK2ZhyQI+OC9uivM6akJkiGKJrW8mPXiHb5OQ4aE
+Zd3t/MCnGaSY4jEMJty2bhfKT+qR5UjOnQQP95ciaOw9UyQm6L3bui8uwIaoIIPUXE8Iz6meC+A
XIXDTZ56XIC4bzfbCvso15SkWpIkRouI2bfOKtKn4jgTfReLJdGiBymDlQ4MUGR7MucWsOA+Hboq
R2mBHBU3YvBbK/HYXwHE7fIGsRYAiVzOHd6MT/PIMKbEDVR1o5uUsPk/5BR1h0wzl1yxYVJDY16U
nN3fThJ0H7FBESL3M2DeoZMco+ZzI628Qv2+pYf80dGB5oWkxEXg0aKaT39IO05jEeCui08E1RQq
Zo7autKsr5hTyw5YxMoHTdRbctLTTyyaxa/uOP2c/2dQvCzYL6PyFejUDaI/8GiU2zx42fkjEyk4
D56KKg6f6rL3871cpkQOO6EP+t2p5Xy2xqIJtwlYaMCvtjpEP4nvVF5hq6sGqvSJxopyL5AEAfy6
v54FpjSo3yJTjEERT082tOd+7Lon9B0iQAdqVSpZlB4G4VtJu5x7T3OlXkMi31WkvqkSsttlu4B5
N8nhPBLN2CQ2BKdS5md1vj9GzfWUKsDmjJBI5wJ2eNEZdljaYs6qM6/yT9BlQ9iDcTGPlMbRnmBP
DVMd6o2yMzAB0nVmlw4MFuOoGXtvsmQoPa20XWUIq/9MBo0pm1iKAWzwNfzxsgopw5J9hAiThtkJ
h6Nv3EegSh4SHjD5oUuJ8DnJnT7RgVLvKuLIasdYpkzz89VEqTUhAC4yUj8bk1eMDlwjv1eCgBTe
+XhAFcYkm8uWt6M49TjSYx/dwPwbHGPxxp3yBCZigjW170RhEB1sTMHB16BW/0zbjj4FNYs073wP
ICu6+B1KljRLtAbTMuAzGkyEtTSrNvy3TpXyzLTmXXBf5ojse6gjTS307KRtBqf1226wcuBnGITe
E8mhp5gcNLp/jfkmp2NiKoVFAX/awZHwr06ZanSb8HCMxOrhg404zDV7eIDWNvbq/j1I5v8k1PaK
xJsPlpISKhOZJCkhdMDk+ciw5sfEH29W2FunPvmAwGpCtnKNXsa6Pil4mzx3O5cskbrFuRPx/bWo
ZTwck7CZo8e3k3ZSS1OuPtJPtr8NKy3OTHEenZtuZAmzTTPOGBKRwJEfmokhi2bNLbbalKXbpIzJ
tUnpw2XWsU9TlLVQQw8+iZUk6seMzAcbd3m3v4abMFNmklW1bvNHVAPd0KvJru5U3CNsa9mSlwqq
gtFfFEds0ikMn4O/BEHR6jSPHlFTtw9JLCwZA7wJ9vYtHWsIsFvsh0ocMNbnSkTTA4DNlJokbYbP
chNI1K1TajRHyzvEteDoon08SWO+O8kkFKL0rxXch3Vo5ydqC9HRQtpIahKAO4h1xhgj529/txQf
jceaJxEXftz11yOGoVA6n0Cr2KE9z6KZJr2tPcra4+ODDp3KkEF8TeJ+5p6ClLiMiyQaNaB1XlWJ
/YDoe45mVOP7KSZGls/0j/rA40TXdaJ9d3sDc5YRGtIDtOoTVW7KZ7jPc5FotPgl/o4livHnep7d
6Xp7egYqGvHmLQwfNwfQfWauLAnQSasr9h+ikAV+Ipz3SY1upZxshD1CV5a8FEVlLL0lrvFxNeO3
Gsz9TbaWlTgZfpoCHM7/6bFC0B+aJhIKeK03YJlvVqcIjX/a51D6dmH58xGC9T39+vERf0274X/D
AAt7/k+BIQXcJiw21x5NXXOxwKzJQJ0lWNbzrHuE2/a9JVoQTZBKikSgn5gO5FM/GOhTSXtWTqWb
lJALYOOsAOjHsA/wiADv9bqwKUFR3uyT2giI7Vt+yRwthJXDjY/42kuVDtIIskXnnGFEVN65i+dG
snpZ6SXs/eObzMA0jW/oY9kg8LhKuqX0RKtY251k31p5ccTW/8FD/+QKJBKOXPhNrhvpmuDGIt3E
cSsxLf42vqB8OHVdLg3ly+dPTcVqGsIoj4c++mWlAD4Q3wJBHWzejq7i3RqquUnKLaOlOUYZVTFh
W3SL5zJ6SGBqLXyRbDVcSbYFGfhgiRIL0vopn9blQP2xiTMU3sz4xqTZQND+rIRjcKPJ63yR9lbP
jw+uLdgDAkUi5bMPUhdqdtjF3fyuJdvRGBs0X26e37/4qPqni7UbgSNel7UEPPBA+lkqlY17mGKO
L4MPzYP1z0upYFSRNnJdJDtGK85Nwy7Cdda54RkZiO6mjz6Z5c6uRuBR2+3g3VpPvamE0L7lGxCF
LvDzGFxExJU3Xlp9rBMllhdiWQCibLT2wpYOjKCHCgJUF6HDW2XEBJXodJiiifclPBKnKfmeGWra
rpySNK2Il2b3mRvNionRtZGB6VuWGIouDINVIjbk78KP5jlzbzS4TIf8+pW5CnoYw+pU19WR3WKK
O9sgb5mohBeePOO9jKeF8DDK1Mimd5XlJ0H5SCDqM1X8DQghMrjjHIqTGcjXp2v1k32TJwnym6+P
cbQE5nM6kjCr0fwNYd1EfS6MTVzytKleuenDzDtUVV4beDrldZSq6dtYr2Nf80eAHdyleD2Z+5RH
e5XZYvScaIZ5gN+k6h/T5F7btDqL6PTH4EGCAjhXYXo2LT/wi5gU5vXEqUZTx9KoJnR2EUk405UB
44Nt/kvjNBaRXwdIHdnzTlJfP69BHOVQJZ2OHgp51OctHt6wVUF/i01Vz+YxkreVMhfrQCn9uKax
TCmjsM62rqDTS25PTOEtmLgfzsnsFyReLiNzXE8Asppbg/EyB9FSShDmkajhwwUdc9hLljZKh4GC
P/ahUM6TAQMkkzUxR0aegiJVacJZa2PvpZuma7PuGbpt81+4gRQMZFwxWz5deQMJYrJsahlMef42
9qVhKXcwOzppNhAPJjdzHvjlGr9WfjNLy10CqY7vo3f4fYKTviuieTzmPu8/juAgMR+MDci9AWHo
hSSJ1CZDtHYlghDxgMu2GskAhRue3nRWRpfyUl7OKamq2kvN2zHl5miTqNltZN/CSlRSyi6N/XZ5
QYzBEluV+blLur1BKo9VPuMpWxX6aVfh2znHch6jnuiYB82I1gpPh7k+egW0LAPxg2dfEV8qtExs
PqaHY7rT7oLg+tMfjYnqTJl8NYyyJI6jQjSuUT6GxPppfwayxR7IVlWyjlTw3LdAScGHYu3SnNtu
S039Tob9XIfGG3rknx0GFOlmqIstw3DARhFfnXQfIwHvIec34sQMnDDyScBPXTsKg6uQFYi3wdct
1QCzd7ZqePgWRs7x/5nQBbosOuEkIW3eJ3zr8R6JfpO6TTaPUVOKBFGEVR2GVkD3JrRiP4A1sdu2
QnYnX7Phhizq4RkcGeU0duMyLIt4u5OaeeXmgaI6cOUF8RsMNEmN/Vhe+LEZFLYeU9WLHP+17AFe
FORBJQnoo5U8l5+tkMBkUzFg3Cvc7GIGnOp+itQ0MHkaLsTrRGJHG5nOMgv2QW3G0OAkvKIUZnT6
q31vAdG34Xy20vnRHL+qtOIuT0tqvus3WNh7kHqu3D/CFZm/39rt+yKftfnvy/N26Zu1WHDy2sev
WD0BXTNk4wFzl9gNqKBHbRfnYzghFu10Ic4bloDkUKtuejg4F1wz14G6pnyDZfVASZDZ+6LZJpri
ta7ThJHnqeYmFV/fe0KhB4EguyIaYpGNEi4ysjzpWlU3mrdv+tbYVquJoHiUjCmk1Z3s4BNZkepm
hDGhEkp+fUWFo4q8pxnpbVmTiu2L1wkLnt25WI1s6MJ+wxBea5zadp0E04mF+ZpjX7mmcAvfoUhE
talVzW/vOmWupBMJcJ3P8ZczKbl/v5ofruBlP9GMWUktKvaRrOMHVQP39htt038Nv92AmYpKcDrN
tU17bpvqvkYGoWUPMYd8zBmn/cjM2EdmKYFdviz9CNCgsw7H3pD1z5qfqCQIwHMm3xtNSleb4/Dv
8t5GmuaUpxEgq9tWyalkJVPbIxN+HNpbRXnLOoxH5X8YB76DwVZpu2Lq7/8UtstgTTQC7v/oIGr6
1Bi8fYeX3il3yM9ef9kTbyBC3fvi/47XBtaFVaTdfWU2wUzceoNbQI3knRcVJlnTLFLI4AWn2khz
Z7z0wujlvXliFRxoL03x/jYd6uDiaILoerlbPveqFRdkhZAQ8gqQoT4L6SSYhbomvN41TfGKdGoG
UoPwLrrL+ZgPyyj5ojMWdRycSdr9KhbvB/DpzzAGE7cdQSV49y46aH1Eh8jmHd70HMeYiun+XRog
Zhhuypl8ri0YuLIPyHkTfPnEKH98amf01QlTxS3McYYRgWR+uN+2nxop3E0B+cSJ4/IuHVyrR2kp
2ATtUwY3I9TtIbrGaxPuUW9V8BRbh3HirWtis3j4xCDOtcyyCcbqlfRGoLs0DyOuDrb+tjARMk/I
x4fkIuh/3EHHwG/3UStXK2zeNNlbHeiB2N8+XSyv0HwHIbGwT4i5s4OVEtPXpUj1t1q/NuUSQyg1
aqP+yEqnG0fTU1LC3nFW4N3UGSAjlKnU5f4OJCAdKK34ajCY+efYXFTmZ5g9GdoURv8UHOvuiNV6
bqD9vLdJEIV5fNwzNpEyxtVRD3HRccpaVRsuRBtdHrqJYFEnxX5TnPEGxkK/jIxwjnchiqQQfXNz
zYwe7d+juGDAKbXXkJcJR76t28U2gcDrwQ8ex/z3foFE62wtxQTnJameSjt/tIlQmJBPzu+HvKLz
+TtcYEWpl2K8VMRYbjNWQydl6j7bmYWgIVXHvsksdoHSTPizaF9v5c7hxpLmN5uQE0R1kst42ceo
Ti/ys6S6DrwvWUvelC5FwjDYzxVtFPIBn7XrSiQOvtbglmzNyO8AV/EE5pcu87BhL5+L5kROI8CE
fn8GG8L9SYYKcvCBS/44P+QVGA7ku0KANtFoAfQnTGaDD6olshLYculSQyIYJoGk1JYFy3HOZ15d
YhSoY3QeTR+BprUuT8kDFErmoy+ufwC1BBx827obWs3f5sQI2w1cKimmRDQ4tP9XjVldbFQjR1zp
8J/BTpNrQnzy4BuZjkbcN4gg7qrW8EeiG1Px6REybfdFB8ps+SAy0VQuVuzXJFdXz6tZogWImwmB
AWCqWqM5UwyxwGBxhcf9V5OJCMYfb8T8Rs2iwlCvpyxR3TuZ2+24+I8WMM3RZNNlafGCa+1gxOZ8
Vib1c5aWf4wCyP9b05kjk1R/BjB6bsI1fxivdGWOjhgFkxosmynJekTqks1r1sIIcfdu7w9pS2aG
XR+LAmq5RJAEAp9snTiJJGmdk39oXT1gHMj6MLXfDSy0JisyiN4ILb9fu7YgfUYon//8f79n1/R/
YzN8TbU9Xbn0xPozsM7CyIXP3tFLwnBK1Kp3s4RSwXslSpjWnzyBZSb1eEEOgHur6eSt5tKrussH
z78fRjucS/Tn/O0ChXuZzJ97+LwcYTJ0C7i6YThf/aHkhyQpJftkF2i/1S7QU3t8Pgan2JRTysDF
Si0CAPCV892YvkiiQqfJEW0JzEMTLkjF6Vkr+deO8ewKvhTup2IN4XpdCJV6KVqDvbZ221ZKwUZy
M5GMy5WZnKWmAK/XQG/E5fc2gTcMAjanlm1zMT4rr+G/TNmGRZDc2bajsDJNOpR/bTxDJryAmXIZ
zmMjd71GqDL/gkn9og2QUUNCyiIPYMqojmj2xe9ze3XZrBEjVqur8wFeJ59zJzQKxgI1M05H5E3c
YoG4tWxqs+1gHhzZtsRoXXiRrTcJpN/02QHgPDhEhw95tEUlKJUTpWP+HEYZYBLWjq31DUeh18gm
OtCXWFQcpRv2msHpl+jH+TV6xqEyK/tFNAIPE17Wf2amDGGoWMem775L2EFh+/4HT7eXFgqmXIDq
Kut3aRHIwjpD1wNRlzVz2e52eIjamjjoxpLMN3Qft6YPCuc813wAqUFVFIgU+kIRMb0KUCiQbKcE
5Ku/L3DqeSml6b4vsG7LDJTbHMfuMnhiQMDUV/B63W7uWXT9r8u18QKAnyrB95BBYL8WcA4uprkr
P2E8dJ5PchxoSH73XAsAz+s4SU8Ajr311c+rF7vFPMsXIvSl2yI1wbOAD45ynA1LWlXYXWx2M9ik
QfwWmDL4ou4//8spQqGzoveRPKP3MUph8UPIvy2oWtVe/d0tEpS8o/fh9T08NpUMihpLAFofq9q0
eVmiGciXkrQXg+/V9XEAk3vPZ5PbX1mUTfFrYgPG8OCveKYdsc9GCZVkUQbn6moPMossXtZ9U6Hv
AmJ2WVWQm3RLI0dqi2T7v6LrBIMoOC4Btt6BiOBoeuPtzupjrSK+PW8UkQw+o3Qy/VeKBv3QnDW7
K1C2RxYGzxNQ/Ls+q7ZJaZ9ABgDI3OXuK44tM6AggHOhz0txY9V2i01rDnE0Zn7ol4OkCl/LhLNt
SDgZCmdzCPE74HuvLDwVDmGG409/Ck0YRSjM3YDCbDSx+Rg+8tw0ixVPbslamlAd6szOaJmlwpfC
aLva3L+NBoAwW4DATkeYUbaNT58U3e5NuFAwM9mrI/kci83uO07D1B5EXCDYrFjrouVrA6my1+ZQ
XP63l0aNc3FqT+kTXXAKTkRg8owd/tm7u04AppiXIq9LVO5Gtft1Lgfcg98Is0YgbubLw3Ltb5MV
jeZGJ92f/S1wts9sxDX8sGyz8DTjx6/1WN3neEUmsWq1eHoapqQKATI5vgNZTbfA75Z5Lp/yK3Cr
GfyGNTyh4MeSFYWLdM+G29eZqaaBOUdeLcHfbVQptGCutn8XKcfRsi/BF0+rSaFytzfFsq1cQFc+
AwGgjBbVVPiNNJF9lC9SlWIACdAEZmy3KVs8AYBgkRNcl3IwsE1b6E9bqt/tiZ2T7GoqnoKzcwYR
y6e3bnvtrAe+BUjnAdRilIu3gR02D41zX7HxFRYTb7TusjzDlBGx4Ld7dsGUw9ZYTqPPtfeECJfg
+SK5hHA3wTImmWwY5Nt022Pu2hh+62bzz/MVqPCN18koVPiMPCxhQ7n1xGtvptPvyltZP5fZ7sLa
o8ZRYqo8IFiS5LwnyzQ7Xs3Fq00N9HemflXU89HvXv+0wxBBtqSduPASYw8BTnbKj43M/TuNhU0n
l1JqFgornFt1oC0tH0g1hJfVJta0+G7gLzWda6BS41q8q6MOg8he/aAXTO9wA28qwnGJW7B0z7HR
+pF8neFy7ZNq5PIZ3FktLLj4gpLHxItGIv9pkB/YXHEpkTNoHWtFvYSAf6tM81zksZG991byjtVN
aKWuwTqRRcYMKs+ag0P/4wOGWgfnF9G7mOpQOtGp5KDRWQhfJoTBFVPQexY8BIwXQWUXkthBtoIk
lAoisLAIHKWo4CTZmSAy/ouLqVji7BTWt1lUgNNOvF/mliUKsZOGUbiJTPJ02RqNHuN5mhfP8E5V
bjuSsFx/9YWtW3/bCgZletIZSNmFu5putlWM3UUtO2rHQuXOKCcwBMhlX1VUEmi6GsFmkRJjE4rl
DlULroFcJh+2/Lsx47zWia54TdrU94KT0jP1HS4zzuAF+1H0JqX81/4Jgfi4g1U1Cxnyja66DUnU
WEULZU3QUgT52U60WMvtBq/Db/lYgYh55/+xwrEbCkLgsbUGTuqfK9h5PtVyOyZ9GdDGXawZF4pI
nPyIT0ygXRwlaXPCgU7AaKX2i69iSv78YKexgTW5zqFHRoEDM6DzsGEOiZaukRe6PLAzBsZA2EQU
KIObfLRBpk1+NYFglnZMV0oO3qbYmX9Gcir2B+F6vgFhVyMtFLYZM0/WA4FvuS17pxX/eK6YOE5b
H9D+heNQudj1FtFLrDHCuRkZ7PKVP+90GCN2y93kMsjGjTCQxwjwY0E0pzUxrBCIBC0zJ6z6LGB3
4XIKbO64p3BLR39ii1Gx0swDPlkbyGkxJs3/SW+JbgG3G51srgyQQW4uptgmpKh2Et70TtlxOHxb
en5+1YUVWXhGJ/ev7oa3U25z074iEfqqvPyv6I93cmKp3EAOmwQUfmpXkGYxbF+hssuF4arbsA2N
/gaTXm+oRzMNYHkF5TR4gvkVwl+EB5mEkvFK2MiklLIkkd3vWR1cwbPLT/OOLW8EQ5c7IqkFrGbe
5ggL4kBsCMFWdpIQNuP9Ag1j6/Qzk/ygvk8YSjQIKGp4aLBHa3yfweAiaCBqkGPRIKymxsxcG7Td
IgLOent9Nex95GPcKEYSdOqxx4EPLiXmt/VVOU6RDrouHcb7z2vuO9jCcAYIvFnoFq58O/dOpvKf
OT8drVQkR+jW/iI1O/uwdeh2y9WwjvrQyG3XklSXUSF+3na/ItgorDFowT/ZvSC3wkfPWSPqf6ZW
hGYQU/CQWkUUsC7jYQhxBpN/UJsPSRL722raLb1cIwz6KQJ76hmKRcBgilSxYzc1d2f2SHaj53Du
21lkOsmRT7zUHUp+FIsuRBPvL23c4PbsToRd9ynTs2Qt9cMyiSyNk4YYFpJehZ3TcdAG1BqiuBo4
uo3ynokktjfjYoYNGGP4+cLBA00XQTTv5mFjTVgMXRIEbYi3bAJ0PQ68T+U5mGvI9x5HrwcQ5J/d
Sgre1Pl3A7fQ7nhOTQ8RxY4ajU4qOVmhXYEC9vUq9Kr90Am7+ej3MMw3pqzLZ+sfbGF5/Td66FlK
1Zx4mQEIpzSWm81Bhi8ZznFrCf4wJNQ45WOSXrSzdaj6ErCofhnJ//CdZgVQTJH1JtE5NMyZtrj1
GBWdTizepqFK9NhmHU4QrH25Hb1+4I9gaoB0vX0U2FH6qAhaR9TLt0SAK1VHzdpJIcDPinejjNTx
NOyg6MUd+4j3Whu1g8PjH5hMWFEpTtPB8kW2hGQOrmhKgHus0k5M5ra2BddjOn9u3q3U+73+yaDP
je2VFOvtmlhDgeIbvumXxvyUf8RQW6elRjgQRJ73+iuD6KhY1/xKluBYF+DH0/uis2OX9BuNVk8K
I75FGFRSmoVrlwzgzv4M6sb5yZPjlyKBbkMWZrjErqd4+ro33E9cYPxeVSZjZTuoYUjsGcD7mEwb
aCXAelEDB9t9mSHOKBiu+PKAEROMl4ms5op34mra23lsFyHxpvBX9Aj+/Vg172ZPHDDPjeIk2xtX
GTYM0h6HjTBXBXnOQYfYZqx9Ekr/9uCvTgzKmmBLjFROIIKfUGE91bA1EfLNo4XAJSWGzGf1Azg9
3vMDvWRTo7vX4UYprBWq1sBI7UeRDq3dmmsfdiEBx56cp0nKAqHALzK6jGQrICSpXK4SADqi9WgH
mxJ3WTKutENTrdbGKlCztbc43/i3wMeupm2FYfGxn2u6mRGYBJvV0zryoAIK5GUN2k+UUxQC3mMf
c3jDYj39DHoAn5gnOldKgB6L3AvcU6eOpIFx8iFyKl8okt6b+7IewkxMu2I7X3pqtsQGAEgqem9E
V1PZjYmGkn+gx0Uju5s92si3YAC08Wm1S4PbuHQZIcTsuDdsfTN7n7WRFJGHoUHQoHCRZEqZ+1cn
Oq9cbl2aOIRiM7GYxqmAiL6LqgqFTeWFF3dBeyzUckFgTQHjTrh8egEm0aQLOusta+MaN18OvScy
iO9Q1K/0K1O8K+FhtMgLE9/M104U+xYAHu0mtDqx162kkFcfTXQUl77wHrhQNPlNnHORSKTeJeAh
N1xTNyiOW2l/xFQ4xIZJ5gzM8RE7m6aECIu8p0mkZ6SeL4yRxypnelArOZCszyynmon2ZuC98cUc
qv/me4kGJcMuPsZaWxJaJETLYSdERp/gDpN8sjVmg9xy364gm5OONl3oNJP95GT80iRUPMKJH3+t
D8J4vcfWuztgMm+ZrpNjl/t2uc4F8/f82+AA6WxNRslHEiCG9e8u2TO29p1G+kRb865fy8UMw0eQ
E7rE/+XLpjypjsBv7rNmlW3ztdin1yU/MP/hccj9PRQxq4YoM50vHTFa1HRYewPnmJ6jKOLVZbeP
Bcnp6roph/RAzikjAuogJjo3lPTUAgLkaKn5+lUjKS5COu2HeNH5lAdp0rZq/GtC17zE0obIQLpp
KOcug/wCSzhbR+IardNLXWn2MA85PjdqTr66Z7OOyTL77pSVwGAOgqwABrj+vsenbAK3NKGZRFnt
2qOkxwaIJ43O/1heSivAwalFG1F9LQDR0k51TBbH/RgBAu7dJqR4i40AbuI6I/4hjExash6CxQD/
SzhEvUXmdpem3HEalUs+yHRM/GMceXuPldNJX8TVHkQU0AfD/B2NXAVgeUHxo+3W6575z4v4EZLo
I3dD9vGiEyE7ECSChLkH85Pcki0zwxqg6nmrtEwlliVQZ1URpQCrOi+4F9bWN3GRK3esgC+L1wa3
Ncg+nwvOEhA117KAMjQqdmLPrrGKbGQdo9Q01keYvKAA9odanzDGrd4mxIhFEtoxwGCz7Hj2uzd5
Iy6vySdni3nleeAP1Ptj4/ErZ5+P01OKjjvXqTUeJFtfMrHLwYlqiPBBIa/xM5Y1vhdpl2cT/VnT
VUBExdu+7VFYNQCX+GHdGDXTAL9kacUmBm4vFN1qzDuzyIpAgA+VMdVGJDrcueUPEar5euh/ic0M
O/VEM9EASFzbGUGQgw5kZo6LY5asY+LSIGt7I/FnZFSKntBIYEK/US6NZoNitcZtTGfiUCR0Xfc2
kHt3bfPafew5drlZvk6BlcM3HYW907r/AgFt8CQIRQBXIV/VYXyK/3jYwjlDTBUr0C9nd0NoOKEQ
/E6Ox9KWqm9xPJgMP32FH/jZasX0AkgT03U+b8GYSgvmkSg+JZg/88LKdb3JD1+BzCkE+iYmoRnU
AThks34Pt9A8dzuNNvpHN2a11+Oh43qkfks52hVg0nX10/4rEZtoM85Gu5CUdUfAekcSO0yfYQYM
eFuTYjAaLLi4PjvlfLWK0pgKjW7ifZHM/I47H1tz9/EWDYNwrhIpa8QQFzBaf0DxHCgdNPK0OtJU
8vrzqfhwvQjbEfljA4f8nxzQ+oxYtR3qwlHkcw6u8oq7d8Bz1/wzESIQfJ+YirVkxo6YwlQMH3hD
iynGbNCesGJsKOGjXILg0b04bIHBWtopp5Pz8GO3swFhyn7s5Wlztf3g6HgPjVw60bWA2lAYDUc+
QOb5Gmu52cgKN0Cqjyfd/hDSsEOeaWXDwe0QnIAJqhi5EpmiX3r4u29dmGJg+s9yTV/U0Dv0+CTo
ddBKVvk42vSXBhU2/6WUt8UEopCIcBEH4ebE96mTGUVO3EMizmC4BC5+yeX0ohIakXI/Z85zMids
kC+yyy+SAxp9mxEptqWZS74qU4t/OO9qv3fosFXdxE7Jy/FVJw6rz/hw6hSLc/7NaZblfJN3oSRG
aKNqIxCN2+Gpr3nEhfFrdahyNAQG/cvH2seATKtbbGcj4O9j6A2qywfDHKdpOdqzsI36KMsWfiCo
7ifi6YNqZIrAOOPwFMNiMJ3PjqnsmgF+rdRlpa4pY4s0pxTZhW3i543v8xBPidwMPP/R074XAQ/2
nKbr/v+smhDGrZHTXRfafzvahouSD5A/G6QhhZ9vk1NGgcx7Rc62W4uMWkcWPXIZqi6BL3TpLlCn
44STUt2RWq4iJ3eJDXeFL07oZ2aQPdafV41zTqOuwLn0q05HBzsl50YqeOnQ4zqle/SdPKRBfbke
nQDDzzstu3errJX0qEuao5Rzb6ECM6dsN37f44oYHBgW7YqzCqQ1gUIJLLTm68UqtY/CZcTYrPUX
GyUa0AHeUAl8v2Fgu2Z51dyINtaON4SUWHFHVQNYbmUgOMbSFJw+z1QzbaEXGDfwR9D0szTjbm2O
s3SJKa5jQHuBiCg1D3UPONLT8zlipt10ZCCY6g8JLINU25CSsVJFfiskiDUEo+bRqLz+z9dr6iBz
/7gKCbshRYOYLIbbObJSYLbOLi3gWFTj16DVwHM0Q5cYXsOUroUKK0LK4gVDnU9QBdunKXJkjlU8
4vsa4gYHMbwXOtECLAbCDtPgb2/yjk0EGas4CBliFCEoJc1ykiRVzk9xIq7QvS/vH2/RfCYa4Mlx
APkPtrPmJvspmuGs+NJEX+5vRKJZmD+GqVWkQug4IiMvhTzOBEJQ+DhXDN51RbwvvyTjtjGEPbhl
KhlsI1hhfy05ed565l+PtloOjxEq9i5ddSnvcqebtws3gamBHVg5LxO4IuBhWsLFI9lhXW/OXY51
p2l/92/Hsr+ceEvVgipL6wnWxF8/af8tR9CMMsJhjSrhJsoS7ou6YKZ5iF5Ar4q2w6CpF8V5E/aa
BU21752Vg4U8hKVQlfxT0uULEhBOPqgMrz/rWTa+njnCm//2RlRvgxYUeRCMj3TdhGMANjj+eXtV
acVlg3EVs4DQErUAPuMfBtHXtouY9LQJUHOePGfqX5SvxbRecvL+Q/MDaolpnSyVuHBgFjYzrbWi
qYTcRxSyzi++RbbBAwtf5EmRi7FeONq57sxV/Uzgj7oS1AbzKrH6ful9+9Bf5iIODvGKfDpYWnrv
eIRgG1L2lL4BQEyzlfwn0TJqdk7MFAsy04hhA1PsvUo6uX0daGlVpVCw5CafWsBDYxZXHReoiLIY
MShAg2XlX3XZre+lGh8wiw3W24FRzq34xor3vIFrhwhhX7dUDgNqiIDkp9dllUd2V6jlI7BRdsg8
y+PQjNIXMT4k+XfB2v9AdEhin5yiRvYUg541PMpnLV+SmeFBKpLkKQZ2CYGnuK5WORSmYNFrTgPJ
ruvMRwXOeYxhnFZ+Ma4Y2m7M6W3DcGcN5X50GUiefYjxZW9dqluo4EgUb1dKqz8cESls+TI30RJB
TTtWN9HyHt9CTKpPjV9uUahErIjkm5QTorf+idhWmA5ZEpHdhCDUBOPwC1bDOFTbmrnvuVVIK0OA
f3jaBIXBvWmh+7946cWdThNgtbjzmNSmYT14epivVt4rAZzVYxzjbId1jVHwKbGpQGxyLL3Sn9TY
8MwoFQpDdB6U9mvWCvnsjkM4TyGxZQBpGp062xQ5HBxrBsXNM9QrZY0pEUjAy0E0t2Vrpr3dTQGW
Inx1pJQ7pANLIjw74nCbS2CQqRoSbduPPJwcTQGNVvPTg94t8MQxhCpJTGGhfrDn7qp0Rl+Zfsl1
PU5EjG8AGzg0IQkxAyHIC6e7VEleXDvAwQsQ5KLKq7ejC67zm2QJ2IZrjcZ3w1E/ZopNUekMouYs
2pqp5l2kkQDbLx/A1jQQfN2DZeX6yS9X+y+tz68YMMLiqb1EmLrQ1M9+aYNFmj7ZkN6iO/Y0KzL1
zp7rNvC5shl8k5RATVirwZNEnkl2quUWn3aRngtK9O/FVtW+ggyHPDFLdCGXp11tvogTDaaZ/FZS
DTtu46B6DHJNwMNQwZOIVY/VxyGI9rHh7uOP42jUb+f4KOX0l31NgFuCxNIFpfO/t/OETag+0X/k
2M3JxBz3ayqOrQuP6b1nE+Zwv1t/43snuVnKP+riByeaUt+XfTeV9kHcDZfLjUUip3uQ5V94zv6E
Kmo4JQNHiQB5k4sja+bPLOkSCSGdESFIQimU4sMXzYJiD02LQ5hCQQ/i9rJk23H21k0dEkBcoAkk
Nry2WmamGkmOl93bSC8xbbBNJ7IHxJRy/fahzu8BhGpy3zIs5Sw+RpYMOXrhsvk7T3eYfyA2M2d1
GBgAqCHobYZp6zNEpvGPCeI1HZh5hG6LibYx1DHKnT5IlbkCKXye22IIti8Gl25NhzA3D9f20CNA
X3JEsLRz0+TekyG1KVKooAuLe/pkDlD7+2l1KyU8SzxGObcPPq11cAk9+p1eVZJyYrOLZCu/uqt2
hj8glRa8SyBU2uWj/XKLj0+YjueLApGC5CrTnkHbeF6C0X3o+ltW0yXFVsARJJMoRQB+hWOsJ5t7
B4hzrd7hCjNl3cp/hFArj3mq32SmrZ+UHCJAjgzXSUv1JCBMm3HLvUQMtNO8YwnERTgssn9uqDl6
cMSZlOTbsln36D3Gho/9+P3FAaHTOZwtbE39Vw3wh8/ETtk3cfPX1mq2xcyUrXOMBL1gHXiA96Ew
t6C90nN4e8eKcZfWfK4sofBrg+xpah8sMJG2407xb9Wl0CQCZ7xVrS42MnSlq+8041heQ+SGzIMT
OAtwK89enarJaIBIab4AewEzOxKukRhzdcDUWHWtMl3jFpAxUUvryYqNC+h3KLfWWmlIqbvMUBiO
3k7oLWqCUqYyFkQ4eHIy6pJI4YF6lRZAcwr8HNg48v2aSnNwuJg0DncXSrZlEaOIH+TYBPkMsHS+
5IUnlGtdJpl8ZNoxrZip4R3gETB51KdDpNC2YJ2TleJeIbpkWiCmhBJdq5sAJujFG3wu29sVaSAT
FaTR6IHy3OMQ85+JuDYbTpKbjGPUzDy9rsq6PcRrapqFflB7aZHWHTToLLq4q5o1Q99kXVdfAHjr
Em1bly72Vo8iDBVCrFHL7dszVpApVO0zn7Qvi4zWmJYom1uwTrJiWBhylK/cnDQGW642MTwH90kv
efuh8ZSlbrQHN0HidwR7GFfj4tcb29vx83SOmnCFXRtKDjID5+TNYuXcir1E2J2f2nXYZjkb8B+U
wFltUkiflglL+QVe1GsRSNRkQ2fQdPJqXwGZlRgw3cv6ChcnwkmlBXbUVInViXn/6ph4DLPAaDDw
fdL2L+ywlwLdGAFGaDb9AzGoprUecschtqLG2XXoC2fqCzleYjY8+99W+nEgy6PZ9LLQqlKXz96f
7XT2rEV4wLa74VoHJYr1GZ54xWHE89tOokQPV7thhamcuK7S1SvesdC2JrcnlLLq2PlkZ0qECy3W
DGc1YyZ7OodJXSmR9ocSzReAdQLSklshYa1gDoHWN4eMUsL7MTIw2+X2ujwUvCDOJYT0O7WAzfTZ
tnD5NFtvjWbPrJGObIrptRNxlUVdT1XGmsHetVVLj7nHtlwPcNg+rykkBejRACnO2nZ83l6OB53E
G08ZVPjoteSLrB/ZtfJHgkC5GOxjnrwsrnIKISiEhey7WotTLKA8QzvdxTgk9slIfuvG+PLT5IsI
3wHLlxUouaDZsmXEnaW08mzpp9RcYXQiXV8Y7dYu+mSvCcaEQ4aiVhzK7nv5JfI5tOgIKUPFlisn
I9ciOeAQtbY+vLqOBgLeD+iHd7S4LUuxon/Qd7n6k5evsIkHrvmH8TW5ij5o4mUO3NWOo+43aufa
2pMd4b+4PHgtq3Q5qdy3/8S+QQZUKJP3xX/DsVOZPjox2R3cdo7O6RSRbyAxrteeyXvXOE7mNAwY
n4UJIIOtqCPb5BPSuizOGwKxg9JIFwbT8dfCLhIxKVCGUIqekzu16978+SFrYwiNL6Lm2vOiLJ+R
NqZvMEirysB5B7MOcgqvfrxlRyFp+0eXIOcNutP9FDCkB8HO54+7Jg9Na9/Zg1rIVj54CiKJWhZE
ONQYXG7AjGoBd899sA22FzYDx9WzmBcxTbFcGeQO2FCtNlJk+7oxLgmqSeDRAniEwwL57oW0VoAR
h9zoanZY8K5wNPfT+IrjU0KAKtgAWqvurVyIX54VRrr49tqKjVhD0PtWaVM6u5A3wRm/B3a74Eku
aWSDzkxs5AeYG+GMGINuNpxvTDfO8rKxtViHoaBelCEIriCXiFHRml88+FpRR1fW+tebfcTN7yOe
osYkKgJPyI4HCoSZRuFkDC8U286pvfojcdPpHgDQrCTleanroQJInlR2vV64c3q5kHjt6IHy7B3p
VFpeiX+ms2gzBJMHp/Jf32+M7p/JDbTh06oalsdhb/d4p6p5m6BVWpPcMnm87pVuXY5+pzd8+OU2
2N3zxMdJdPJNcCCID8bLPHguwMWFFA3vx0kxWjrFd1tchh1ZCpeDT+IoXV+sJg+0WqaA809+Tiof
TQ1DH2Y0zcD7cCOVN12eEyfVoTuE4WjELtPQ3TncTOP3cUu3NKugfGucVKkeXlbNzVCUSXQgegq1
8EFdXxdOc1GVj7MkfVsEmLx5ndNXYcqCV/ormvGijQeTxoX0i55PvrHuSUCy6HGsK3SVWRwmzH0e
HSEjQY8bqjayvRXR19F3vlH4if132yd0qOvJdhon835qeIe7soWfWHmzPtwXFl+86PAZXVDhvHeY
o5G9uTke8iaHgp7rZpWBqlZxGf+xsIYbs0gdNTQHCwg9xzX+XrOoiG9+Gz8hpYf3sNW3RvqWXNLJ
FZjUC927gy58BHyC/8YwZ4ywKEVY1ZNg1WGSBl4EOSySWfn9ZK1aG86IuaTPlqiNdq0DzADpQBhh
PNzJt+OUHB53dzumc6ecK7xmGmXktoPz8ZIqhvffw4Vq8OFC4R8YdybRcOF0k0Uk3nLiGKv8p0eI
IH9pGUjpcApTuVjXh084Igs9jW4okfWHE+ETtw970KowA1P3cVUmZAOQFacWzctwcClvBTYN/jao
9uMwvLlG1De3jh6O/M0fB884ik1IFsTb1SntUCRXNrO/E4DDWhVHvRDjCp4AMjwgn0SJi7ByoKtf
Dymg3F3INPwUwwhrI2Q8DIejjfOo76+JqPw8kfvv58Eb+HUCIVQeomaXlK0SayM00I1yaEJvfqTf
duHT5HgqfHRF4DTUfWtxDrnj2b9TOY8MDIe7fxP5PkkN1o7ugXoX+7bQH3K04p9fr+QymWh+GIOv
sRK7cGNjICitlXfVF9+a5AGI/xKdO6uNeENcIBINGr5vcP6lOcEinhA7qbZ0zB3WRwpkcjLE9WEI
7eoq9duxTds0DFJPosd+psY7y5s+PTpLWGgNHCAGz4Yivk9Bbqh2/LtY0XYH4r6eptVM8McXX5F5
er3GQu0dcWumhYa869nM24tsxxnLbufKF0OPAYPK8wCQtJAPtleZGthXYPVk8W9ckxyMAR+H7lSg
8f/GcA3PKeLLpMLkfrr5axplHwVHfGem6/Uddbv5kBj2CaGkqiUfjiCdSVY6uP93sr7qN9/BueFx
Ql9iCjZ9Q8qwTbboPOPJVaMNS5vLmIMMnRCw8xeUTkFLdFwXWIamBxLhXYfBDCjNV/p+6sSb2DbJ
MRb1oRXFP4aJZGRKPrigUFTAO+X2kKXaotPuj/Eba68Roz19vQCoSjz9RhRyw28BboQ1akHvd622
K9QKu03F0/pfg+E4csfiVgyvcRIZv7XR9jPeioSYfZyfS4XxlDxl5WwXq9j/bOZbkCeruaWkW7NT
Xvxud4wsCDLj7f8ywdLHwTH1fPtW/hZfPnt4REep3wOco7NfCEDjRwGRACHbxN4gIp6VmX8s9Yjz
wf3Mcq8hSEZfzg6gNkUarqfuC2dLXHsjkFTetvBZJOgpD4azTeQFnaDirVIK6ki1d+deMpF2nfVR
r/tZFE40Zf8n8udkBTdSfKVLJP8toHKULperf1361LqY5sXmfHCvdtXiwwzFNe/njAWr46Ch3Qt7
hpAjZNRXKhJae+VvONZe8C/KI6DU+hzZy8McXEbR+qR/2PzZaeeUWCMmM443RiKu8Ku5UkWbLQwb
E7qqw77IOdQ3NsQBRdcIwB3n11lWUBvNreNQvxGzsnfT1w6J/ppvQV7jNcGMLeEop8fZ/Yqg32Wg
8QDiuSBrTGrUmfIn8aC5PmoyDJtfE8kUPJOBu0Ds9VzdWg2jYu+l4hk8vsh9nnIX3CvtDq0Cyz3H
rEh9MqfuV2g/c+9bSEHJ3W0H41keYkZf6gYQpMn/MGdzieeJ5B7ysJcTXNF7sML4qWp2BCQJY4p2
fqlU07FIGOmo8lbmxR4pqmy+7nN+DE9A0cxTG2d5QU/L0+ExqY2TFuk2yr/wRTkv90h08yS5jsrR
vBXpuv3gCBehuuZLZzGAjcilSaD6+zVH9AoC4VAWgKHQ3M3YccO/T/an/ZpNwC38C0ZUkRA/dLNj
pkMuqcUwoM1xS269cIz5gS07kH4kEGWSNAiwSECH90IvK8bBW8vhkapdLC1fNyI06LffKkwAYbq9
V3YNWREOtGZr/dsuy7iq1ceTPECHlxRLDHRPVRCaxt9IbVZMyUHMgayZh0/AgiiEI/tL6Ld4uEuj
1+cQIHu3HhAaMaeV8xEsIx7/OCwHVBu34RvOEPoojZneV1GgvwDMsGXKSw4AJEEmI8/AYYsT0Ytd
U+wgdh9YUo1ZMH8ikxhfZudyqe2x5hghoxMv7xH0UyUdCHlDesac/Dw/AOcQT3Mr8H7UUP7Q3w7w
HVpvc9vDOzY9deayyI/pOE30tCUGJZsDH+GJCPN6Q+yJPlTf50xTmFD5V+at562CJTsb0wDNFPp+
R6tjseH2CikX0N7Jy8bIhHSBqWUpTcIejw9COPxJI+pJlXsXKLmMo6n2J61AiuBk4dt56IA1DiwI
gz9Dalt6HEhbhUePhQl6EvOkE1cLUS2gZPeUu1KPoCHrQJ/bDyaoebz5lYS8GzFNnhObHA6f0szA
fd+BMiDo/+gkhbiBlEquABhdOXpvEtzSQ+92A2d37TyWgDJTAn2kE382cJRsOKiflFyKOY26EOvJ
ztW6oamMTM0dvN39KhCcC0FbHrClvKW/21YY6Y39KEISZyMJOWs3JtUvPzuVA5YNx8O2LdVKN9Sm
3NXj5i5lncHPH6+8trluOOxzUSA2PnW4XxRCAyyVW8VuvGgJeELMHDub0n+tCL+STTD8U+aCLl3J
vbU33bk429sQ5uXHbXDI5psXiJlf2q6oDYpcjGl7ZOpy4aDXZhFhx1ez+YMqTqqA3oN8MnqGaAF8
tMWQTL5vgbNmIbnwYE7uQsEvrkzSedoMORbep/2RvP3eB0HakXeTL8Mw7eAb/kT+UGIAz4yDba3Q
XSS4gNvqYaOvMwEbk0XcSgRIkp8Jcegxqx7NyN3e/QI8LvzioRXy1GG44ZyPZ2cfIZq5EK9wCXSb
S9Bg9aHZ0vUgaHOPIg59qdwuhkLLFt7Xha20cb9B0IeCvlDv4Sm6+HG98plEvY90vpwSDaZr5XvK
HWFegd1lf+V8SwRMgHjQ/79n8cRBg9BW/Mke3mLYdpAJ4qU+OxoiVGS+uQHzzl70HwTu89bsxXGJ
LDxQu6yXXqVnorf6uToiMTzlfdWxJaXYiF51ysXmqY+zwWv6S7aQQZ/Vl3HMgtJSxDYTuVbf8UrJ
byoLBunogWV1dUIIUSUqzPudzkvj0f/qLaeoBYbGPzYC+5MLDnd9R47jIQeY+Wsg2zi0nTuGe9zN
vu7tAmu/gf4LZtA623x3rt2HvB0iqLzPyQ7JMekKQf+EjVSjFr9cgiRvIrJVctcM9Ecd7FG9dgfN
2DQ2VsOsBnnXlwInzqI9sGQcvK//UPtF/czKaMweLv1lr4xJ+GU78wbak2J57SSpPUDKKteARLmx
MpOdr/pK0Wm5XaE3Mnezlqm7Eo2KzMfxNMFX4ga4LcMmMTeAV19lxQmYzU1w1K+qoMy0b9GvG7uH
TSPK5vJUPuH697HjiEOqCyQKXxo6gt3g1oX/eyYyQFpWdn9Pmlp8POvehzwoYohtge5+aNEhGnLN
zttyh+Mmc5iuS4vind1fju9OBHXsGjsMhHmdGjKD/J7uIIwJ5TJ6BAtXMjDA1mFTMZSV0ikkvqhU
eDy6ksfhm5rdr8KtShPEihHDRKu+UljfkniCeCEXyoDPKW6coAaIbvmp7OcAt5xT08tZqGiz3EoS
RFZbNpOlEO2rkxe+TmoG9hPkNzZEq6KBMVD1xz0iSzVt0fTCIvPttJyemvxObiVa0D6WTY9LHZ4q
4lWALFvvd14IlSPZGZKSsyL1qUjN8jM6vqoDdA768OpXBjLTRMpntJ44ve2rL+tmLvOL2Oadirt6
TlZ6BTtvgqU3Kj12hg56Rve3NSt4VV6pgkNykkK+HLyxTyAhyKo4nGT+MJsiGkxP7/r+5N4RIVi5
+gWt0+j43jCmosuLEtZXvK4Rx0ViGyyTGH692XKHOUuze0uJSgylY1OokSyj9R4porksrexQmr+8
3pdgCOEgfTY+Azx5zmhQdfeL1GVigcYFQR9FH+MTmlseCoeIeeTkBMuKxv16+8xKMjkBvTB+ssil
w3uTIrc2M6dK6pOrPy9C+vo8gP88G4GqvX24sfbKL3MpKE+ABpu7JY8ltcjvqbZa3i6bpF6vslOl
RcMfyKV4H6jnp1SMUosGaNePtZaU1ZSVlcJEwZBki4OWUFKPpaG/WmEZYOAmQUN2KX1TyiL35U28
g/+e+i2btfMsdIJ5C7JzbSLXxq5K8NR58h2IkFGoCBYmoQTWnXxkEHzwTGfrYv5WSoq8A9fLms9B
UzNy5ovWqI/vz3ENBdEMSR0UoWriVsJmboyRp8f1xo5Jubvge4mFdfG/hXncz/Vpp3mq9mDSA9bB
ZQZ8NjSpjOTbsK3cLxFIzWYdTaQa+Yz3ClZL9INQ8/UB2LZxPVfzzBWYyhz/uS8+cFkHjjb8sRgI
VBvDGAKHmF1Djj15NLGMr5DMIRLOvSj8dJkqvVZaNXNFmqC8mVITwTrXEt0gpmMlJLm8EYt2D30I
Uq0CECw2Ywtu4nQdIyoc0gcZZ/xEQYprAJxU1HbNJORqtZhTxciCv8BnD3Lbaica4hPAZK63Ah1R
3tihAKkbW9WbDcs4NZIPNh/4MwVeqLRvXokIbie+Qct7t1kwGJBwzx7WfpDA0CpCqUOaRIemTCZk
tkDZyeKZa+Zthd2ws/VXG82x13opYadlYF0ipu4O1IIPec7n1pbaeD82yRon486QWWJOdNlfdFvH
9k3Xt53abHb4TtxYDkJOqX3sg18/qeWu5o0WLazTnv6XIeco62Rz+zBUkcKNWOpiSD3ACqoHfWvG
obNcl6zDtka0ShSIzgNCgSivnM8PG7rIt9Gx3poCcvSEx93Rlg2CDtD1kz7zRmtYR/edNs1KZAwS
IUXn6L8+am5y8WtqYkw0uZ+Qz5INQqzRDYDojCi24v7BQ7Q2HiiZ/OA92I/kEOb8QQVp2MzbUj8G
m8chpkjq6Y2fdWqg4Zyn1h7njnCIg1xIJ3XZPrGfGj2iLiHsYpHCkUsh8eL6Q4NBYqYB/WjYQOF6
SSKqD/s6y9gApQeQRRrhdYuSC05+hNLrbpIjuJDnviwBMxYLaH1M8DU5dGsdKvK+L/10Q4XJUahO
dUanQZoy4LfrVDMZIBj+COUv39axTGKRWq5v2dVcBdqmtozL+NRARw4PUXukeej0NA+ythjGd9bS
c/Gq6RdHVZOcJ+mRjhe7H8xqrrUpBaSPIF/R3Mhbw9RuGuJ4i3Lad7y6oSoeDtgyJvmPPO/SnpiI
raX2SiAA8oMK/Z7JqlH4Xfsi1/XISc1k2hkt9lfLSJjB7hP/FQ0xxJSg4OqndfNSPAMNdmRAHcZO
omR5SfQx3RqVQGosq/bB3RaO69JWIN+HgHoVgIqMBVikhXl79FPIwfF/88YBhA0YG2PkDbi5jP0s
J4QAjk8u+TTVFT60hjRlURkIvRi61orTjb91DmMqMVZUKGWrv4zMYH6Bq8YyIdoFlIXrN56An/dg
fYljqzB9UJQHCC5G/pO4I+hK0f0Zm2eRCq3ZKgwoNIhktOwHRAhKxNzW3TfKprJdUAv1jcFdJKj8
6O8oOsA+bMAmfZuKvN/jksVsPkffVy51oYZhF6kVOP0o8nZ3YjS6nWKMHHZhojow/JRSUWoMp2QV
VzoqQU0+0as1QsO1jzuqYva8WHPayIg8XF6a5EqwAkPZ8bwsLsgSuBKoYX5oQXCmavjze93SljTJ
ZD0b05LW3xauCi/qsBAlMD9foQ8QIZyD+EcrpkV31HUzeNjk8c1rVGlGAld1ploykmpwMnb4kxq+
4iywNlEgyilqqVAoTuvssjHhYlsroQLBSfAgGIJ6xYyTXUolyYnJP8ZAmNsomJ+maoX1fJRKLOHX
0+eKHM9+hHM1S+GNXFsSq5MuInWhXXtVXNS9wEP6xxQy2HRB5NFTfH5aXnsfMVONho+U7zY6UEz/
m+HlnvNCgTD1rkeBhmEPMYZXc39Q7Cf3zETh1UvQ9GjOzo3uOZD35DDnFa6Iyogl+pKhTO6CALfW
SnwCHQhGkQqKmKl4ifXba3XraJfKf1N8a4Sq+PpM2+XeWrKlrqO1Tx9gUECOfXklEAnPQ7pg/c+2
1sP8gyf2YWapr50qxmgB09kcFei2B2RfND196czWc94i2MD/5Y5Uw9wcrXe5vOXQm72Vtc4kBqvA
SBCVRwzfsXtam3yipVgMxdlcyMibxtyFuJ+/u+PVQLoFbeFDu2aIVTA7wIkYV6dwphrFWBvYqNYh
heHtiS92rCGYhuh0pAtaOWoGYPycVlpisKPaBovvwlkoYKyxTfr3FnO73pI8TNbeBYouM5MMwAFj
zN6ae/a0cphFdFRwUTY+CGc8ssu4VSw3dwUwLf+LmQ5NGgB9wE5gTcZaIqKrQu8PT6AZkZDF3SX/
/jPKaXbAqY6KUMIiRGu2NvfNFZl99bzF3HMqBevSnW/UEdrxelWBRdOodwx7Y9Z23XTtxMzRdvqT
lpDENqVzZX0e4aOOb+dG65e4S7LnmdiiIEMIPN3Hfl7O6UL/47oCxRM0l3vZWUILgl9kq/qKds5J
LsmQKV3RBA+eu7cZSQY3AGDt/R6sqBVbt3hEs3qRAYPCWJPscvnKo34rbFDxHEE47gpw0b75odMO
kIVuDMMp04DL+4CzbtBBTl0Y28poSEWvBUm0M8A9hG33b4bnDxY8JUr93X7p5JHwLuyw0cKjkcgN
kcrwAHVo67nmS/jkMy+jNilUXeAYa5DOJiCk3khPwu0e/BEP+caovK6RxCYJDbB27BX5y4jc/7BX
YZYR/0kFzwf3obeAWKIV9NqXZAG1qABOW4XYKoIYrYQnAjKprlcKP9UdnsX+8B4RyzH7qhSfPiOh
WHEbF9x2bmOG78xFVFUBHJOKkD7HVrZrkIgWuAffJzhYAM7Qe+ZWqRqOnkqVbDXgZ41jmK5gU0NI
bJ23s8tXYz/YnieW8rvveh0iIshWnWyJobJXU3wKCQVgWxTXEyrLQ5GP+Q1S9vdLe11DACvbkstP
E5szl6rWURwXgCnRtscDBjkSIOfxMhjfZUcX2Fzz0vTvwRWZ9LppGpshgQkr8DIT/g6aUrirfNZr
JvtJc8LT4CIBjEDuAACHhR60pFsDepSktBSCf7Ssho5NdQiKrenXo+RScA5QnVoeWgHXkQb3zKLT
ORss0pBY9e9g+PChdOgmpnJQtFCHeOT6BqY89lY/zBC1NU+/D0LIrUV9zll5mPOBD2HzJkWwfomC
OiIzHO/HnnLkzybgglVS1scEDr0t31YASMe1B/j72Uf7PnI63Rkuf6WYlEzzV64/hGuoduV3pv7S
Eg4tL5UvGfumzEtuzK3NWY2MXi51QMZwR756zW7PY/RdMrOIX/oFMml0ybaAU6uNdIq1YvOHmgFE
fxgrmAWrXf6v10DDnEbQ9mmqzDSByED5n2aTNHYP9P5XSXK+2fcB0BY+/ZhcL0wonYOcI1+Lx0dW
0o712WHUwTLPyzxRc9IyxfkvgOLgXU9BlA4ycVXsXlG+VVgBkYuAZ9E4p/F1caZf4MoDKk2spHxV
YoVxC2zUZXEAPC/SIYak+aA/XA3spbb75dnZdCJdx2ci5Xp2UPAoR9V6nByd94EjeEWT1BhDT3vz
FOjiJwGbQW6OOtol4jQMf8tlU3PX7W9WloekC23pPrdLEuVKY7FtH7aQTUfuxaf3+z3VL8epInn9
B6KcuBz9qRQ3jLF6/Rf/SRo8PrfklTGgCG46W42m4JEBbwbRDstYeSHBQQ4bl2I3iCQ2qXMw+ZNB
V0HeAGxfAOyEECY0edSljpacHHSrXygO13a+oYl9Lkma+By7Fprbnytnim+1ua2WqH9XePcMzvK6
A4aYqI13fH2pX7l7nrO6vVqN4iIlE8LOPquhO9ZjD9DuYLVxCjBu56wvR3No6VyFHSyrOEjrKVtl
/37Ct0k4loKZ7g2pl6P4fQbRaSaZT1nwS40cpiGIFoZupjc2C0t38TfHLerdxc9wwoOtqDHskNYg
3cHWxpwMU9G2s4IU8nUuOZQWwb4k9TyQZ4sPht8hjnzMGmgdwNozA2N+PkkLC62UDky/U4o8dpzb
UToVlwmky/PcPmYhGz6CoUh/OeM3dT4R2yy/sh5K3a5hhmDiRcgn87aYilX7NGwoh6OgLsuQ5Op0
LrssvvPUY6iJoeRf2HvujzxNRUAwAp1TTzqgtaMeoa6mZEhl9P5XhcB4cajSF6HJMSgpN4TNVqMl
3sYmejQKFO7368GIetsMbgpKcp8oQYtl1qdmfXCUNDcP2A5KSoWTUZPWpTysvm0JylUgCCeafmOa
D47PQrj9fdDShDKviPhol7X1YRjfaM68Dw1EdrXyAtR54ACpawy98TzEwsdd1bk/PvXJ8JivurVd
PUV/UkxXTZ8gq6JwZG3mYZGpuShZPsuOSRC6xiD8UCVjmaIBy/rAmLThTAazXxmP45KP2gIpvvk/
LkSCaFUNVZX7X9GIzHgfa/IZzebqu2PLNAIHGYEQod1Yf2MYbPJ8H0pH2/SpbhGvzUPiP6fyCo6F
G/uFeNnQaHZXKKkesgmKcniafQvE7CvJmnU481W9mA+JzBwm7Fwl0FW/Byhwzzy1YeeqZc0tfniX
F4WIBdZA5/5XkGTXl54D1fheubOC7JHhMD9Kzqo7L3XNL8PdjCsPLnnmZOd12IAplbZLimgDPeMA
2J0MCmnp/20JQybetCyEZztF8dMJc1v+zwo+i30cDwbCiiJfU0Nuvt3Syx/R2F5y3StH8CAS1Q7/
D5l7IR6Pw5QVLc+mwLuTjJthg5dUSCtwzKej3LNRTJyn4CNDj1p2z5dygCW6arC9Y6je2DCZjMMb
Jvy51TT01ld0LmId7DQVIU3hVzg2NExtoUu8FCJFCm6JKPYAI6+3alZKC1RorNk/MIPWmKVllgX2
n3EKbF7N8CpOy+9etOJujNxVBnKiQQIt7eSEBM2OM1h3v5sJvdoI3DkBlb5KebuHlXnYVS545oFL
FtWkQuub5lrhYFTYPpGYSonrwmxFHOo5i+LoJ/2sSg9/rsRvrUMGpYXTbAXOLHgPATsx/iUHTF+c
u8SggxYU39HyuSFIyOML1/Vt/SIhb1Vh3C1SDQ+CaFaoOYxxqyDUz4ngY4f8OSqkRrY+U4riUdJr
Qtkmmhhjg8AM0yAiuAuWFsYUMexwFFxU1wKpcptfpav8E93X/tbFECoqZ7eUFKnzAGGzGT+ZV32G
y6+M6VwcYEJQuXwEpyuvualnOvus61kIz2kmyXYh54hxgB6yEf73pkcrxJUtU9GuzcEqoWfiyLda
G3ZnF/Q0v0DpvNwMmKFbBoC9VUnQM5N+fTLyohVKoke1JC1gMHoiwOQ5PR7+os8VW5SxPqft1Iyx
ZX2d+UwcC8RAs5j7B6+IeEV0uKAE23w1i+F3bRv+4Boaa+GCfGSlkERml7h5CzYARpz50OVfDIb5
1Ns86+SjSd/2sUFjaqmPSx2RR5N1diimW9P+qvasjbLVdKopuiES7nP6qa7sIDw9UT+UAxW1uXg/
C2RXIlDf8VBiR/mgUfBUOATE3Afhn0cnJk/EnH1V67BdHNWaYRTlFPTp9RjLKn9KviWHaUuiCcic
ALG60iEDQ0KledNKex9knWqqfqqZLQs4N6le4oQkVPxlGTnKhb3gc0Actqv3I5XoRF0pnUHRRDHD
ky7OvIultm6w0ttxdwHKLxpnejQveNHVydzqJ7sugHOOWYMQ/VvW8tFx8uSO84wN04OtvweBGy5O
W8DJg9T5R/VZIxchhwRerqILjtaAa7liYgzhszG8zL4YYRKUQpB6nLgOcHllpMcJGte7ClVLu+6U
C0XBqjzFK0h7OxbXj7ibnVUGoVAyLTtEnyfE/bzAAb7Clgjm8B5VgjvVK4iKWz+aUlXIa1B0FbJy
uhvCW4mb4jYtzTCZSUiKgv/TulMPwAMI5K4QlktFr3NG6yN8UNoKia25UDSX/VcGUZcK3c4TkGWE
Poi0T62SQWTjp1km2pIfsq22M2uWOr6uYGvNIL/HQJqMfJ6ZjHndjZONg0DmUAQhCbBn1imDlkCo
dA9ZtaOp+lCUTPwVTlNuTHDu3kCCc+alePOC5F3YRbSim6mm15JCWyH520u7G1l1IK0OxI8tXs2Y
O/4FgB0XbmlMD9DENbY91RO5zp83gb70RO8jrdGj6gLhQyOWOiPdIQCDCW/0riIRJ8iuLCavrFCo
LGvp5QSuH8RNDh0TXxwDRlim0CWb/Inc+yydkY03BBFJd21hekwQrZRxL+OkjRyFTtRIw6MClULm
8bHXs8FwBBhyLkquO+aTh+vVcBYgTZ6W3TwGpmQLpQJ1FNZrNQNALOeKfWOD2iSzXaFU7qLiJ8oL
Nl2eQLlISncbwEFfoo9pf4M9hHXOSV9xzZRaJ3JG9UrgqMWqSI0P97bNZvmXZ7b0OwUvZfHoudUC
BvreFvphbitkMGZQTqeiaWWPKV/WJFuv9y8gJAj2H77qt2aoKx/l88VDQVeOqxgJgi3GSPjWdl3X
audxuP99W4AH+KCq7sqM1zH/tRAedU7/6Z9h5iUu54Gei4xdnMeyxfH39K/ayEFt8IF8J26jig0I
e3NjkUZlbhef+G2eAX+xgOubBeYM7bsXAVunn3MJKvPbiDelyEH5xK6d5E1M4xPDT3s4y6GfVtME
90a+Wjitx2zhPnomGckfRCLvrn9qy18iqygupSptvq6aqaJqnSOHaglDajfOuUtSitTWG4KbuaNX
nebCCXeBe83cq1FiY0RNhGWVV93gau+K2pClw/P9ouIkBJEm66xtOdmEo+vQW/KtVAqq2F/4wRq9
fBg0KcuweqArx+naN7aF/83WN534RCkRCxKyhBeW99niunZvtbjOT+NXIK+XNgSt2dwRWhG3Ubwm
3Q5HjtjPZV+Ry4m0/vhH/wtyuqceohvHAKeaekh809VmOgZnYLg+2ctQOc/esx+sfdqWhdPorgdS
fABdPkVUgWqPs6uBJHkNqJp+19bpYo3lTz3Iw8TrdM/Ba09G73Ev7TQgVGt3PLMr30vMsfqN6XqJ
X4nWa73bXY3r1uJIGG6a1t7RA0xvQInxyPPceLRWKg5Avo7Vqsql6LYcJYtJCnURt47SQ1ncN3JC
V9ZObRUKT6nvqWu35sSBRUV9UGXFs2OJB0xAgyf8SWZx/JDBb+Xa7heerFBOzkDiUS0wdI4P5jY1
zg5CwP/FqAs4JvN4zcYcdds3kfxw+ZRtk33xFeW9S7uoo7FPIwmXNGpO8TPY7e+wfT0OtHxZKTxq
EE4/8abqGa1neqgSqNLpj6PruJOTkiDuShk8lfs5d6nn2EkEFnsGs44Lnu4sBty1rsiNOHPyiMjQ
kUjy+QEsPqj00jhJCZAjmFYx9UCsgmGkUVPrt3uY5A48iCvgqsF4SXgHEdK8Ol9xB+TTZ5eKNSMU
zRtVid1i7Qaxz+v2NLR4Yp0D9oUrfXQqE+gBpG8PK7dUipOQPI1dGhxRnwNHYFdqH3P+B3IirFdX
9ViT7zxAGY9AfM8knlrK4jCsb3ee4k2YHdViYPS0kXDIK9QN9gIrEVACotG4SwOAyYANo/BtcLP4
n4AKCmIlm6X57c0Qk7rPNLN8NOck4Kc6/cqnQH8KVjUODS18Xbn+IkOB7LOIAIFtpD3jwOFWg4lz
SNecnO0sUEgTJyvW+dKxxl6UD9jilRsWuSOzFJpu4uftdJcfDdeLcvkqo9goPPHfqz5R6XlgaIfs
DDq4IBRXy2RfN9FV5YOyFNVyJnQkYqhWmKaOMEOPxdW/olkjE85rv6VkZ6eK7KVrSq+v3q1nG88k
e7stsC3X1w9DVLYWgmMKvadn+LxeMJMcPdqEzuad0nJls+feNE3qUQYg0rkL0qkv3gsS8vDg45ZC
eqbiJZSRqXoMHCCJ+vFk6Celx/QNoqXuGVKykWhcMhx5DqNHCO1x12BI0aRNLsENuRBo7MZ7DzC/
PGyo1yHlgL+WJnJBOimoZZ4h6OhOxPDZLu7FB2xRNdEmhooy4NXLszm4rf1wTb0l4yLm+lxNA7Wm
7N5iFNqlSYX0EEGNFCvLldAq1yoQ51VCKZ/fXUVMdPdPevlhMWUjWU4jOLXUvhgxLQLQIr3zanlG
v5gInaG7AnrDaY4SrQbNaTBYw/LhrqR5Ke81MMShTFXMXsIqHaMbBaaxRlPRGD09Msdn3yDa37XP
MMSlr9xR44IWWUtxLYWrUkFnZhw9xhL+RVIcCxPe9tZ8crjkhXER57VRfkqlTuEhGAgkY/SDNucP
F1mTuzz7ciJpj9FDS5sqn15i1gwDA7e2Vj7GOPHEuwL90pWDB6DXcLrANwRj9oWn5N1Gb6wHaU3w
NSYcjaxE17YjPXZ09/RcvXi/Hznkgs4v2rLYj1pDf/VCzkwbsvNDziNzFcOpF2bcGv4fjW3WiDfC
VHN/PZywMKm+NhizUTmdkSUiork1Pp2X50JxK6l4snFw5ans3OnfAZAYzzVErx9uZctsUsqP8888
J2Xrop7XEVJE3vtYoctRUjKpI1J4DNT/LwswHPjEvN8ChxhoBe5Oxk/nVSwx7IyNimqIEyp9jqOv
dfN2cZQHpDMDcS59ymxikVEWmJ8s/CHnEKu80r3EI48COI9oa/LMkvp/pZPE3m8JpuUFWY3wqs5X
BylWjjvVQ6F37Qk/eMnD3v8JLxoZjD0cc6RDPsFlqDlKXYtAlrnEOGRI1mMLdoSqbqrw4qX9fYKF
RGC8RCLrA3GBbGB95kB8kcWqJcXQ0k1eNkTu2F/67i2vgGHtdprOaj3CimUa3B/YdKkAYlWDUpRk
S4W3LvHanvQEteo9X5Lmir8ThCMTe/p2KhARsQeDoIOqFa6kY0E5YLz57Rq+OnB60TtRbF0qT5Sw
czZwi/bLJvma8W+xADiCkUObtdkzy5lIJaMzhQbxpS6KS5hfvc6m8LieUHB8KNj1mUTgT2kRvfaR
2RrSLTOL0rZol+4axBPlQPHA1cLA3znY1ZjHmQeUH90IVmdo26IfvCJh0DHrZVRS65vBGC5wM5Ok
oLy8nXQDgMnhzUSGvjzghwRIHl/PH49SzO8NdY59NPQEvUdgIa1Qi4mnX9Bq89epYelYn1e2LLWn
bGvvThH9ngoOo5vqj7BKEZXrBedBAD554fOltWzJyz16tBme1EfPj023IT0lzmO3mO+NbZWDcQz8
iP+HX35XoZQG0w27CT5axNPflNgfpy144IUof2AZPsdEwXsZQuNvi405gn/3nb3Mg65CzfS+2u2K
oVdwwj7kAe4sZDK7hikNVPOjb1Q2G14EgCgndyy5l+0A+38kk8bisgh2us7M4KpvPmScou7OPJFa
fAFEKjwj3LuqxMVOa1YL9HffGn2PH2De5ohQS6ZoavCmv/avgk0M6hGDCUhIPU1tXa3ReiO4ofqV
z7wjB6KNLbYtaDIszsnE036xNF3JHVCNuV3VNcIw4Fw62zuZz1NJihd/ZLtQeVKTnOV2weR7VzXg
kqJdF74+OJd4F4B7MAxxzsoH7cfG1irET+EcDV2XjYcZG7Rc497sjplgClQppJd8vYAvolf6beBE
CZ5j4gw5Cgfi7rPN1spN2KKgi/cbHcR9eeI5nm3eUCZ5AyRxojtvq2+hoz6vWtNMV7vw0d0RroT7
H0ZtbCqu+68UGJDtQHNOsv8QzkEKCgwyJFjwdF3H4SkAKvSpZbVhKIKBGSMOcItQLWUjhV6MDA67
CAvhYokigEV/dume1s6F2pLDeG0G+OvuHrHgDL+eeIUx9gDXCEUTAGrT7qZ/SAqlz4iQm1+gBe05
/ap9TotaGYobmvnnExq0ZEvVfYWNiN6bwNe6zpsfsHBCFzxdJA7j6jK2B8+j+d6XmOsaL7wubl0L
3YbVKWLlNGDWlAO/rPRqu+Y7UcrWLwth7uV7m6rQNo0/k4K1rVzyEjRmdVrRugmjswsjqCX+e4yD
OcE97/wBxWAVRtqX4pVnWXN7Y8zCMjtVPrP5Vgtg1DrL6O8RChDk7PMlD5l9sGL01Sh1lZNUwFQ7
kDN1sqmHWS42dLDkqeQB/kzRHR4e6xVs2Z38Q5XR6f/YkMTcAmDFmPtiqhrqTr0CtprKEhNoW97G
XyyVv2lqlSTeN4t4zz6Z30/BfatKYRQV5RSYAzBx9oDl3iAtYYHp/xi1PgIzrpebexRdSdtpoelr
hHzS3CDElrE0EqMk3+d2hCm3W8E8RNcsRWJyd0D4HvKuUgTnv2EET/hnhWFE/cfNbEUJLCjKE8eA
uN7wTS+OthFFiC3HUmSBxiHRkDkuBmLucaBexxbVXFoxIiYiLorrpALHeiFzH919qEaxJyACnNds
NZr8ccQ0cYGgswSlZ2j3brBPnt+HoTXBT2lI/nsiDCRmyOQMu5e1enRSN86hjeY5bFbDkcJTSXFk
YhHYxKiBfRZq31LCSxjwp3IoPvGO9T04LTq4cdgeNOFcCERjdKsk+kcZgRwU7pBfeFzIRBpS22S9
CtEeGGsoUMig2X65ftfjVP3rg2MG6pf0SJB6kt45f//1YiFQqs/qXv8dz6yin5INzy2FRtmhhWxx
uI+37vKLHeg2yz/sL7Y7gAVmcxGHhe9D6fKTROmhVNkaCmT/lbzKO236SPWPrLVsNnED/JGYTEAV
MyKYggkm+20MFxmJkiLw/1Nhqvy314DasWGfijKTAYsM8xgT77CSKDs8j98FOFwzriAOL6DxAyV6
CzUE7m5w0X9Cg2+UP4+hiCYjeRTdf8HeqhJ3ULH1X20PySX/09ltWcUhaO67Shyo1wyeAOdiJvox
5FWSN0RWeEgOATJSju/+SVNpaYar6ML+gCTyigrLYD+AVkgvdgDiMFdty9PaVmrZcowReciZbCne
hXTUA/3eAVRHSXbDgLXmWdW75RkpAQ/JVeEEumI5r6OwtGE4/iBw2Tp/T05iOpk3PDDylRfHv+FK
B4Ja+VwWeOLEq6S2Dcn8MMWK7BNmAVEODyxEkap5UUMrrnuYelEES1/q0h4avmOTOMV7FbsUAS41
w2t6nnaQsUlXxGvvcN3tfuossr7N/5kFjeKYrwyDCRhqQMDtfEhcHDXCmYC6ib/qajIDiiCMdcKH
Q3XB3Zlrz+L9tTN4d1NVAEUQsQRbND3Of+RFqqGfVcBRGTEOUdZmZ5eVlQhub49fsd3cVRIluqwp
E5kQNXJACWRumWa2Gx+MuPJsV8iOpevwNyihlhpNt7XGkGmVUWUjViai9f3rHISCVAdDx6oty3dz
EyoAIl+JlKUQkroxU6bZtb+Cjoik2EQo+gY+2e9qM7RofEzOHs6BA9gSijPSFY8Pf2D+/bx0LR/+
duaXeQmefbwKkM+GnqIUocB6+IW9fJZpfifpITk+KDlsKnCV3Re6EfhaOXSYLjEQV3fj1sJVSP4q
ksuic5fkVHBmHFz3zhFFJvm1EviO1T4OIL2tEjZ8FdOe0/McBCe17ZJXyN3RCHG3pYDNwSKLJgGd
cbx9pxH+1GcrHAnoql9DPFn2rG3UAxFvVg1u+/Uq8iB0ZpBZIrMyzPmsDZD+P30T3EHNNtwZn2lV
dvS0yTIWoRvYiNg4SCQF1bVKjpzEJI0vD1U0QEcJzKL67NQm6JFY8Xrr7/DZUOoP5PO1oTtyNECn
lJr0ZkosjSl69pxqzyj7E9bbDNA7wkEQh1jeoQiBCE+k1j67djF6yeCGI7KMZ5+aihSUtyXGlcE4
ya5y5mdDQqOtYL6D1Pm4vUuQmT1Y393p920uJR2OFM2zGfZWj2wgGb7VzttxgNhMJP8JimqJpzx4
ES+uocXNH2PFDm6RCzEnJ40Nq5iFhCDphHlheI1GboSIPz3ZKkLQqKT1XzqSWpcMYdT5YYSIvx0n
z/ySh4eEXfm2PJGtJrNG7B8IGefekC2uVJgo8nSRHQVSjZ6/WgSoui/R7UGIr+8bGJECefy5X3zO
5mQjZi9E/h+NElzr1plj9ti1jDJUj1KU3WW/82z7xAEvdaWgXh9tNXFgpbs0uyIxf1zBYLTqtf/d
yvnxxVr0Za/7kdAqy1+rNkgmKmo75jFt/qPKebJFRNIYZi2qJIDFSVmJuD9IeHFPZ0JQhDTeIyX+
1wT42RsbTqcC1B4UXt1PZ0Ubi0Xon5BdsbODN11CWvfI3vgiGp90Mb4OmQeRgr09mJo6iCMZf3Zu
zorkY/2hJx9LO34MwWIKr9fYknXHx/hAyR2tNxvtuZdMu5ehJgp94LfKBw+9CxFgeS7FE5RIvp3X
jHmYQQs96mKgjb0wdz8mb06IXgVKSAAHoo+HQuryvkjF3SP3hfqAyicaspDuc475UUwoSsEbEZvE
90egi60VHC0uEandlxIrYcLW0kC8N+CtEhbsFHDbEXe3SBkVdpSwTl1Kp7O7L2Ml2e1BKpFKmxkE
ZMqVe1OfDVXLiKx6cbqeW1n2JI/DU+jH7Vi8VRkanvxAUOqbVzEY0UYKDqKcrLm1W/A31GxBJvBS
uEfKm+22Du8t9WbZSSaIXo+e1jJN6IOAL7h0nUkejmP8XRO/ZFsAS8A58j+KrVbJCR2P7p3qHTfn
TRg2z8CYzxmCxEIZsWuak0uFy6LZfDHjiwAxRYnBqYqGe/S1XjGBBVVHYR+NRGEubYP3yiq6QLmM
4AbdWn6r8pvybVsuwkmrABODTUtZHVnru7+UAUWj5Gk/TMkOFDfTXMbvb/QeQqwhf6ovE3APlmuC
punvBZrLUw1LcWFlPetEv/1LA3pg8qKaBetiSzsp6silaUAyI7Er7+wvGfLbGAqotA9UDFerO2YI
qY4eVjHtzfVT9hr0/45ucZGHGQg9GoTLj5OiCS6B+iaAfGl9wpg60ycI1EdPLNycS2I6YiDFqubU
DYV6di8E47RMZJPfs+JkP43NF+a/rV4dDPTXV4L39w9kS9UiNdKEtaxRKPFcCWN0Q8HCMQlngEaw
5dUxyeFnb4YFffz4zHD1m/BqlyKYYr28LzajFb5Iw5DqzfRKkxPvO6jKLoxu72w3JNEhiCiTH7bD
UWEJBbAhw451Z7HcqSz/0OuB5yC8tj+/07No7qaiGHRIe76xTkSEjnszWzvNgxTA7YRP99HHm7gV
041rB95I2ReAvwPTgshJ7x0F6g+qc/6dRbMEzmxtPhPBlL8xpjc2FlTwNsmROQ85PHzioREAHKyD
0POboy4G0JLC+wPD+myr+g/o5+wy0kgEOi23B0mSc8uwHk1yawkoaYX+aUgeVuDOMKO9kYF108Zn
h+7v5leTOMyhVTAkqT7kiAdNYPe0h6cH2Tvu11Ah0T9AhbxctVd8n2WyVI56QXGurlSE9t9WzlHb
txaLyXSGtDKCiq8pYFvEtEnl6Db72s7JcnAfEJDR9OivndQdMAGR5XqgUZK/d40Anlr+Uqx5nW0c
HoFh1eFK1OgwaKiEaC3vW3lOjAq9KvdTULiBApfJRQstbdsvn63wVSOhqAfCGVZLFRPpA8hJknXb
SWNmZwvNP7sWze9sFuZ+tyJTNOKgu/1rHovno8YSkexuTH71RFG3oycuDsrGW4IVi9D/0Co9OUUI
xDDTkE9g5FAY5BKbBcbqyXLEao76KTuKNuRW0NWlL7sCTeIaPM3VcoNGqOVvbPKEbOVlyx3RSpnY
fimn82+m/kupRrOqC67uUA6IJ/5CKYRExSJDKNk6txL9qVJtpbmaWq63ZeIdlf6kWvm2HfkmQKk/
GEToX/RSBOcVKX6fjk5GvB+wZFIArQRUzlmyg2Ro8NOqmsw53CeTfkuuhHoA94O1JvA8B1V0ihh3
gXrkMgsDcMPSMyRKCYdoS/HM7pPH1YBT0+EcOhpCKP2RbaCTGYitpxcKTCCBoI0fxisVcY6Iyzjh
wqPn8KOv9OhpTV3cJw0HxqAGrNnStQMvn8zjXvheayN03EQozfGFNhWu1+XQZomtTdxgrZcww79Z
Yg7PUmouMMkxiUJqCXG4FYM3iWP8EV5xvO2Qv2i/nMfJENY2EwS+h0bcqfYZCqaPKXzFfbz/Hcsi
pHLYvfbi1uZ4az03/B32Anb6DYX4NXeogt6QlkgimpPA0Jw0Mq7TNeCR4Hu8t8VnLgXSD2oGBOlw
biENeyltrZbejKCDWhPkX6GZbiQtQjs+T3Rh9JCPXv9jfvUUGuW4vkqY5ARlpwg22DRrdx9kVFkx
8vzPEezLUJFo58Su7PXdOYoVHwKxueC7rB0MhTCPaMH/d118WIxd3CMi70N5r+stRufAg8T+dRCe
uKWOdJWPSD0YEgKbvAgLbylgVPXe7GxMFqx7clZIBwqtvmk0DgjLkweMKFTz2w+uD/vYfB1qsNQk
XAdGx2hgdHMIMNmMpaCwmrNXpGxTUO1jhbGgEsSn9jrr74V4cW69x6eRM9L3dVAKR5noGY+GMwbg
P6tIFlT4DdFdjQAk4d/7qiprZ5nxHkaHLNbg57/RV2V/HO3xbpN3l92oN1miYWv+AHTKMB5TGFtq
EYxTpf5XYtyFOakLX+GlWpRZZbDvuUri+DXytsC4DQQh8R7JnIRfZhsvc0ktFRd+NVKEtorB61PK
jV4kypO/JXtUV5TEkaGH/hE8T4xmHVCEYWfNlNxirGWB7bEVUHev2xJNAwo+d79/l1NLnPuqdxvG
X8GBD6GpUrIWPueT9Le21UhTbSETHDTiIE0o+wzaZrdZD3Nk8zfyaI88g1JalbBZP7qRYPcFCMxE
wV/ey+0WGU2UOg8js85OgaOJj3mFpWjks8z32MyoiMp6UrM1AB6BgAmjr6i0xJx7piNBT2Bz0GXv
Ku/GKzC46sJPNYGVth6SKb2h9BPrPVMSvnkdwDEvX+vzHYECy+5OlyNmPFQ6KKKj7pmxVkrnDBO1
w46IOiy5kpjxVLXurnUGlUKpwIGxdiSaPvlwk0yP8EugvHnuiM43WumazuBy1NebP1rzV4E17udI
PaOMFws9OSzWP2TrNjQvzetXkuLBwVV/i8zd7rRxc0wZzrHHhvVtHuYZzDAWnK06quXROiTD1CB9
3jHSpW0068DprHe5KrWrzV+ktAf8487fgHOAxzwOlfpr+c8MV6vDvEeJmc0p4HqjzKYChy9aaa/E
ojHdHenvc09qLSyaCo3BtI4hXe/cUNoX3tPOY4UwnQVTHn+nQSdl579deoqVr2+5OZgQNn1+u1BY
8KzY19G5lnbA+btniwzb+YgRwfgTFKTzPREIq65tBwFf0OBaDpBv8rPDpU1FII+1LqT+iGx4GcfJ
lnghQpuIcznQJ45KuBZFJER2dFRDAykgTu+afieHX3ZIsG3gpWVR40LKoLxH2Ne7cvF0lXWotYm0
+e0dnE4GiwVaRLocjwmf1MvzKrOR+zhZoRBiasMMajseAFwmQEVtLlY/5Jk8NrVB+0QTY6NE4neA
/bj23sws4TlzT6H0lKuoqPzzn/WjATSrH2/m8M/UozC7YHbYt52zbuyMaXjxNUnj8EpcY2bMa43j
VoDI4zjKzBYvv8qt8A3xDUZoFR1dp5GJvVKxw+dkpxdx9zxQKDOwMkbIxSvYPzwrNXAA0m5WwPU/
8+P7gEM1tfdO9vkBOJQTUKT161XgnwhjI+/DNKnhWqpS3TXIFfIUdIJ2bONPlK5E81jmsdqJ3b/D
+jmGgy1d/xsGt8LHvBJlRsJwv6UQg/rr69QZMOW7OXywRQ7Sg+l2qPQ5PzXLC8K2Y7l9i3DvBfz6
KU56xGS+wgrm2BLH3Zre2lpBxLZPXvKth6+8ap+WS/KZvzbiROiQJcvjgE1jEndjxSkMv53w03th
GsmGZeQv5msNKGBD63UvRMSVTtroycwJspMTp+m+PiS4viiZ3rh4CVC+pE+4x2rHHGHj0EWORlZO
uI7nGI27qbykqphpTdct7DVzd8Qhw4p7FLRTO/J1stfupDKuhpJ9WqFccED62NmcbqOsCNukpRtO
CpTSJmP23ZtlM6Xzqoio4s0udmvL96pkiBxvlMRR0x+4rzTPr9VAIU2We/YDV0C/LTwAHfX2ouiL
f9mIGHjS4xmtlMxGx1wkJ0kUulajmH87RhfPvQSl8qZXZHKRLYj1jxDGGWpvB97UPWSXgvPpdG5X
h4L14DYAa29RWHuXPdYLCNeD7x1Ht3ZqwRje3RLsbtXhfT9dniGhlDRetPyQXsgLAjtjkxWw4l4Y
oQssoj6/JIFwFHiQQASFASJ3EHyOukrBoRGejkB+ssQLywZCXBd4mwvQ5JMAO/MpxjVfOnyE0g7i
1+1lEDb+9UcIF1nTQZtSALoQAfRDUeUC7YjQePQNthBZzuCbvNziQcyoQLM7wNB3E7aSCgqRXl8Q
2DRVJ1/u28jthOxmN3F8HrjmYn5++DfvK0Ji+CfYhu6DQg5OM+uMZRZncveVgQLgz4jCb9093dp9
hoWMBhVo6nhIiunrmmilmn7Ee+i9Ap1N9PiTBAGKy5MquGFx6+xpzO5cIj1+da+wryYd+eOnEqwX
Yj3hxAbBdVVvfh4fNd93B6wzL+eLYB1AmtlcptJ5RDLQqgDUMraait4ivRlgYv4+aHtQ+mAzXvVO
v98WGPW5yI6XgL7YJF11gkhXCqZx77yJ8sQLKZRIhTf5rm2bmzoP1WacfHVXYe3vzRJ2W71Vftke
pbhwWvfkTlYm5D2TLMRNMs6zvTUuux93dSD0chN5TlEBHD+baN2lj1zyy6uG7dQqtRJM3uyPeUck
joRZ2l3kEm483189EKd/OGmE9yDYJr38W8I45+ELn8W0Z6iKOuZGB2Z9l5dEcudLF6AvZWOQ4Oog
k5M1YsEkQDxHeQTp2biaXATlbrzQRydbG0MFGzy4L9cPGIgbPzMp5geNnI1rzXn/yQsnBQDlb1xp
ucZGC2LqMMWtwiI2qinz5vCJ5FJYETXw1B+tmhgwnvJDPJD3n0GAQSR2x0ZjKphRPODCDm5tKrc/
XSCKvi1FlZcLnUMp0KdGWtJtVlErFzcO9Flwh1dt+1SLLFtm1Sln/m3kQLAqznHumaH0DpkznZSP
I5DZPTWIfqTwE7ZPd00UGaggH9AqHQpX2Au/ynuArE8HDkasAaRmIz8KaHKl+pHnE502UxUiVO8+
MUQV0/UrsgvUlFHuV3UinFKtiDiy58FX2zgG3DdXaflDPb4X6FlYiivCu2Ruh53adiK5zhL/7ue5
SPEmUqdSeYaFQtpK5HGlIbervWvkbECxuTA52q1WLr1QzSg6O8XGHtLRCccmuMXmDWLLT8Sncjq5
H43zr75a31FuUcjJ9PAgN/jOvzGAmd2I22Ewn6lITIj3IwlGu8vTL52oVz/PK+N6GVD/qaJW2akd
RchAMgCbaEzhwtYQLnD1df3x9xNwXDRT83dIybXitkdVig5l0iD+QN876hg7qI4oPe3IrnZBDNE3
mZo/9EX8fk1vos+DlbBAdmhAl6C4cVqUkdHKDWmXMHozUGYjaeqH8OsgtMEwMTAjiRNRl6n8tITs
CreCCFV53smbBlinPxOuS32dEx3gE08nJGChdc07qjj4eoaLF2KPnDY7Qgb+u3qlnokAJLznldQk
7APSADsz2pqUgpjiHyqEHURW5+9tbO0nm7HRaTowQBc/RfKQDZqhWls5YlkSuhTfBVD7dTTfp/vh
gtvUNat2MEiQsGR9+Xby4mZ97BJ8HGbM0MFKfnZDSjRLlQtfRd8K73Z+IHS6s4GQdsxwyEvSvlqw
dGvDwlcUn8TxotE7rU41Q38AohBZY3vWBwor5KmGrI4D5OnWNSqBuIb+VfHXYCcovtOgwlghOuUz
4JOKRNAdvwdLtcbuugqtuVhXvzVpnLeGMObhJBeF/CSMUzOyKmyLF4j6OFd+WBTNr0/k24bf09DF
dL+0Rj4sTqKn2eGjY/ZeXuexUG+XpNckHDDYndxcqRU6GRfupGBHXq2H7aQbmxlb/5ufbwhwGa58
6mPVeVbUHc4pGJWXAY0KoC61kb2pUPglN0e/ckWc8/10QGzxPHZ+VJoZ80k34bFI1t77jn6PQnpS
OM4BneCKKv7EKBz10gwfp2ps+Lx3R0NVmymclcpVI+4wn3yqpP1UNIeNsi6AHZG61z9hI7vqU43a
BGuR6skgrraEy4/BDz/zpec0XkImNLgCjCROOeiDuc9zw9jIeyLYMQth5rnrRYwtp5i2Vz0tKYPo
oU97fNQOglN90X1Blm//W+u1eGW7cKX38n/KiS9YQkOx+Bx/8IoaGUYNgaCGAsaspceg6yhjOQ9d
ysDhQigalEZ04Id57nfi09uUhBdTZr9pKkMJCJvHbEldFN6oRfmz9n+sMUSYnImTUc/+uTOx/3Yh
k2p/DmBYpKXWu8ILwpwuogMBzKHWh0BfnRKsDjPXPFJ9nc/BwdSwpfQMb+WG3CuNq0d0iENMq3v/
EVGn61MIxm9iS/YnaQrzoUTMSkddBRedTxAws03Ho8XqBwK2CuS7w+OasUQxXUChkAa3vz0Q6lqA
F+OCUI9yINpoRvjZZYHuWj4ydrzhWN0Hkndsd87LeaMTY+DFjX1Vkx6FBeEY2/sjgmpwecLZ4lIj
ZY2lKcX6r/6Bs3mlkUwGSNde7xB2kHCaGYJ/88S6FropTPkEuLjQlegrohgGViuwMUJn3CpLYrJQ
muGKH9mV/gWmQTV8EuMBnFpdDurnpzJrptRqd+29Cd8VEO6N8JPZuCEbaBEMmdMotOv6vUqIdy4U
TH6KLXzHbSaQXSlxyqzsvwy1/J0jKhV5T+j/KqgY5UoXz0yrWT/IP5MQp+QHQFsTkpSxfBXgDVhR
7+jJBhvQa2ZX4lYBYgPavEEeZ02ygx2Yk9ca4YJDmYJ7VJn/ucJMH+rzHbKhFx73fxL9p+JIK+EA
LPxugogdMQUH+E2q1FdoH6FuaYNbI4tOalZWCovhI3Yw1w66xMVt6H+itIw5d7LQqCTMuZm+OujO
q8wkY54P64zpnmZuBmbjKRtf86uKcnSxu/26DOMbNoDPjxYF5sofpgiIHzNeXvoRcrcnmp+gXVNp
28os2ernX2FhNLPypK4BeEsUyeqP86goWFt5hfpf/H2sRDVcuWBanC4qeCAPJgQyGVjIiq+77t51
P/YaqwRe2ExF9SgyuSM7f1Mft24cbNcolLfTODq8ZhUeGciSJF7sU98AUDTK+rKsUSWrTVJcmlm9
eKoC1OwohSi1CysFORz0zTfWWI0FeMaxvxLK/F4apazVgSZ5AoUfws4HjydYZFmK+bqlWRSVXoS7
XKHHJ5rH0WtSeedkgqx8ZRj96os1yduShRXfOmJIk3MvFcMzA5H0sca5hzQVrRmPgeHZmhlH5gt2
UbWLmriCqXH36w/UgAYXhyWOALVlgVTuPOwwFXTlDCKd6fLqtpmusbJ2fgRaUZiRpQZ8D8Foigcl
xLBTFaYbq8aQpBe/T1yPnyyzhuqyaGN8wi6tNQSvzGF5rA7zkFzkkmefy5+8KkWd51sLHIcTaAN8
ryNEhq1E1THWV6Ywosd4G3yU2PPnCQr0zWqI1x5/u5vPh1GcJyg3XtGVeDY5FFGNxsoSnVKKaF6+
dRnxD63ebKE6ri0nsP3X3W59zCW3qpGs/FmJUzmD4gYqngqfhtp5I7U4O3Kj1BWyNB/iA+q6F3qy
vo0h/DYAcmSWU3Hwy0qpCyFa0pHIKxk/PI0v4sZOtA3iXSo8xQBPcmPpnGVoJjSIu0pKi6spCzuI
fIqToWzNkdCjCAv/K3lo1geprLYYOTBOd9pUCrrN6+x+sFtRYgqAVfoKdONmz0o7iMkZnynJEz4p
y5fTxA00Wtmy/AnfwZSyqR6Nr6+f66sqXCCaO49ubCNCmNBW58cAjXH+aTc7eENmnknZy42V5JFv
j0hvTvcjUoRfFL3zAuO4SAJNgNbNCWiYTvzLMOXDsXb94i23k8Pk9sXHTahvk28FN9o1zl41YclZ
yrrytlj5IBuK3aqON7OcQHYitp5+anB38fC5j8XuPb1DoRdspVwA6YkIIm7HJkgVceEN/wlQjhcf
XH9UDgbNK9X+0ss08qobiBznrf4jAPcED4z8I0ScBmeGwbG9f7t0gMPTbmAwbZZ7MX3JJl7zh3gp
JJMMyscCyh6oNMvqyn1+WFvVtqLh8g0+clOJsjaNYiPuyh+5gv408ayScIG5C0bRnO3EJcPBwqZF
L65rTlOMdiBLn5GPMR9L02cRELJjKoEYBw3krUqMCW2THxlilEwHPSM6/LhJJanS9Nj+igw03GmE
lQXIQWKlEVeSO/I9aRJ54bDPjz0/u5SwOtfJdmxM9zodg0+ZRf6j4V1io901Fk6aubhZ5SFAsDD6
lny7iwCxQcnWGhW+iJJyVKi90skQUWFl14gSqpzpAeRnJYepWMXUfdQNFVJ8VcXdeizLKk/MlxJ0
+7ZJ4mBHJWo1TNMAzrX4+jR3hYBs1CXO5BcDYsN6b16OI8yds6+8+sl1XdhGGLYCPbJq408xzr4T
x8pvCC5z33hsAUHW+i/nlPVC8kh+hmgGEB0dRRWGS9RA64VO0RNbV90N63XNPGmQvUqt1iJGTZyu
5JvD7y/GBLssxpLOQ8tVE3I2NnCz1iKRUMMBkL9Dmcz0N9fpLnMgBr6UoY3ZK9Sl0VlQKrM1oTjg
38LPhlr776rEmp3+ngifkYbHXw7jKip7iuYVvXdQBoWdJ0fGRrvFj6ghsJi9LBLP0qof/xMe/u5I
SYR1Vp9d4wRQB95BpxI6nrdtcEZuxayhEjK4Hz/ybscv8IoLLZW38FnqFZugohEl5ojXdSfAqhi+
wPTYtcjWJoY3si/6irZaSObOj7HQ30gaiubyKtj3fihT34GSMwRuuVANRcvEH99/uYcvXc8aUJLS
vExRfzWMpBMqISEgPwFg6XwbMc13/dK6oyz32M62EokcxxPyRjlkw5FL63jxviJkrlZ2rc32fl/n
7T3bwqgN+PfTNJ+jY3YP3KCFsHMd1y2amXKrMyPB48289Lk9AB9f3dljaJZgx10mGBGpZtdGr5I5
Przt+xd3RtdsTPvmCTKckdIRROOFfZunZV6x0nN2XNaSjFmIwV0CyI3dsaStF76mQVjkyo9vpO25
d9TXqd0LTvFIGinoD+rsNDB1rZtIpDOO8pfU1MP1JMsIA0O35fEKyeIU8UB4G841Ldd9Wg8HDmO4
UZYud50saAhBSvINmLJPXBcf/wqTNFrpJahPFuxSv7WKVjuXpbi5pSJxcJtXEBG4QZcxTZRrlfbc
KMIycDR7zEW5foK6bIwfDcx4fc09cmqQXb63F2tiXtK7Q2lgtCuQ6ilCk384+7L/4iOAYIZdj4RZ
GmA+utliZg5fy9AGleHXhndLsz+zH45aPBuMzLGp2MNcK9ACJxNvUPRi9N1DGKAPf2Xg4fovgj+0
1HyBEvF+7so8gP1kNHTqTXXs2A6eec8p0p8LUsWs2l8nHa6CfUI84W5oiv2b4hUZwOdenB8ku9LP
lE0MxQpL8iL5Eu/WC+m4L7ewz8WhYEv+0jeFLR/BWX8I5G0rYq6M+3e0L9kZ6UT1ZojWrZH8t4dU
QfsiVVjdsCmI6doxgbOnaDqC851dWf3wkVaHYAheRixnHMENowsCFvLxoItjCs/3C7BvX/trFLtv
cD+nCZgD32sEuRwFOPXtYVhTYvqqsDHaYLx5ij9awt/zDg+EiGUIQoegB+m0LuRIbo/txZL8LGKq
jrj16Jw/VH6E4Yq0ZeWXXaIZsGxmKqaJp/UXHkYK2DlQkdUBLv32Ab7BioCf3iwzqjsQO5FZC1Y2
OnyiuNFz6Old9ENYBzKJi/ULQwGMv4OEgiwR7GvubT1Z+9RGgtv/F7I1RuzbPXWSvTq+ecxfaXoK
mpfWzAgyloyhVfiEfs3TOQHlin81ZDOR1XazFREAMNKa2bl6jFjsCRbzK86dGnS3kQLuDURRPIJ2
m6iVbq9lfbaxkIaER7zyeGf7fzREYxNnDzjpKNoexnlh/mT/jkqPrr1v1x4l3ANSwqJFvjKCL4YK
9rR571RPFlLHKB+jbJmWvm9LsN8dTvR2KMVSQL5OS8z7qLcXD9/5Ul253662D4/tbDOnmyuJNoyw
Y8yBLAYFaJYK1EYrTTT7axFliId+YgRvklurVUam0bR9hit3XHiOi4eJHhLgRLS8YgN53mxy+8Wr
E8wTIOYBYoqhkDXHGZAFeDdIN2shCVU9WZlTqSu+WOoGFfrMqUXty/UlbEUXbJxSbmAS1pOtf/TL
H1Rb+yruWhDjE2fnJ2be9CygaQqBV++TgwdlJP2xoEJ+tVYTzVJ/8ogdhtkRvXZq+u9Vy4oejGWl
0MYpaG1vG4lbcQnsqZMOqqW///tZGEXdKtbcnhnuZbG1vjHHJAGnXLhzJstihwL2PIKM+ta5Luck
Jrbyk+3Usuz9cA7oA5S5zKeCyazHsQWJN8rF2c4JuD0weFsexA8NpK7znXuHSKykVjchOflayBH3
uTSK0TDZND92Yqhze701Ok0kxySHcu8KDaPKPLq2HYDEdj5SyADeil0lV8lsoNHAC1PFVoGbeiGy
HT+ow4DL98tmfOF/bRNhn4ILR7V6Bm3+jKTfwxMqv2dYBAn0a5X+p+ErqMAirq+MQJe+wnwF+tYp
AIZa44dD2sX5SpCj8iRvd+dSKyHWGenJsHfE3Azo5Pi28LNF6jQ/kW81+QEbOSbW/l2BAI36Flml
MvKj9Qvn1QaGpOh1HuV9r4I2E66/RgxkMCm0wqURwmFxyMPhl2B+6kFlmm40rUYAt3FPo0rny1ON
z1gXt4YAC6PWoVoXdKDxqgkMAYltuHE4sTWf3ZPy536eIgGhJPtD/FV/DuXiP96TJ+5FZJiOxUSY
rox5Z7nrduil3anLJ7CJ/9H4MCfXOu7qcLk+UXCXI28j355KKsstgM43fOimH1GsdRkqRzM4qYU4
6c2JZ7FPhTKTWXGLcL7XB/nmqCU8bH76VaJWZjE6IIfpXwAtql5jhXzhWKa1LFOKBHbNze2RW5Qz
eYQiu6OnvvPIGXw3vihUWlJqTdW/b09NMvb8VPT7pSMnuswN/GThVgdFavLWU0y0rWjeUrAYw1Jd
QrzDk4ZZlBHo/xhZF2zv2iiHcHEExyBvq1FIZ9XXn6LdlnBB4H14KbxYb84czxPlla1Ej11vC5yp
FflJHtf5SegGf2TAavCmgAuVl3MeFn6YWso7KS7/yGlj/EOq4OtjOTV26xNKz8qe8xT2FRk2Qx6+
jW42m/mg9B0Zp3k2o3TD0fB3OeNKlXApnGOxWdGqV7oFl2UYte5TLuvIDyIR6BoZpW5xBelWqwmE
mOMBV/QU4Wn83Q/qCvDO00wx1dm+M/abtNhIhu3Korh7bASgjANz+B+H/SoqSJOpusBbyXI93yAe
YQoZkNugPOL6LmLcOlt9gWIssr15qJuYrmWyRNj9XCSfVBbM+FsAaIohlgnYuKOtF4MSQSrikkgA
WmpIKww1RV7eDUsDLY/s7ZwNjyX1ONxGkzZFNEpUKxlVrfxH3Po8ZdMaSO947TDnfFJ44I3uF4uN
sKO5dC/iCUgeb+nWaP03R4wOqdtbLmfffqqKPaAyx7escuhdt56FOOhswCMGdvdfNRC4iMXcKFQ7
U3ib9mR0Wmk+nl2nZcOWN8MKJLjBgq14oKALmJ8E6Y5F2Isex1pGmOFrZp5jEccC8aYDbEfF8lil
bEeqhINqs38ncUpzk8sueyLWzO0V/HZyO/9q/xSabhtxVc6IRgElbrId6EIqDQkM7CZ+egE5fX9v
wBk93Vnf9STNpmDBnvklZJrsM10IWOTJV31SsvKaoOph56gNYm9d+mJhpMMcGenTnm6rv/Mj+G2U
AoImELNXbmbUrh37Rq0xmEyTXR1WFLWittfTKOQkfBSptOKIZLeamS6Ubhq4MXRGf34+6E3iXtY8
0u8R4l4CZbHzSltnOQl8oImvUIBb1oHCoza+rMeEjuJuGEkhf+YSWNHqTzbirM0t8/bkFGBDq0z4
PzAoYmKKFNPuBaaUmfhhY7XJMwOJ+homD+0txHR+JClB5aCHoDYo/gqd1vuhmw0L51Ybul+EriNb
R0LPoYxklwzNhB+LR9jyFTd3u/3HdoSVhWzLBTO7PbhmkSaJfKsT1UO5Krofpp2QHwscZ7Znt8UN
8mBuYkJV62WQycLDnUh4FtrOHuHHtRcBgWGlHsinkDdMHWx7o/jAYXO66u2a7gOrfl9zODcYyK6G
FmwsWW/3duCdI/OBNOQ+UKuoOVAQjLDLWzDxB+5R+0OfV8ieckidD1f1dT8sjOhblpO/h9An9izc
pYKJITj88efH+/BzSvcj3EAq2L13D37mpF+GWnNGt8CQ7AonE7DAl3j9yIG/aylzdQiuaezLm+dk
9t6JtdeEjAwjPQ9bamhlOxxLecRDGtOJmXujSyNlfx9m6QxsIlFgAcL3pc4145epAUgbdiXAUkXD
mhtCyDHz2ClXDXkb5M9Td4ZZjZcYt2wRqWG4gat9W4gO7STZ5EB629TQfvgJyYGgA1BU5zF5YGgT
wt2FENe4dz0COMoOYfnATh5cCdlMnC+P4ic0pxz6xFPoDdrEL9JpXMoYFqIIfyhpHbmA0pYvj2NW
Ff067T3ygZcZUli4r2pNay6jl9kcPb+XD2bxwaqzBTAiyJDr7gheiYhYOkbpR83aYw8uGD3AB2sd
/4hUrfnIHOf0SVoxPi+mMjC9twezJTasVWu/Fp4l+o6VVQHKrPGX100eUsBGAnD80JCvT1AUvO9y
wk0YAwQPXow8z+DeMfzcFeb8CzzNleiJCw4luyQ3p7i2VCfJi7k7TLu//e3JPeLKOqYG/1uEMhKl
XVPbE1axvXRvjOoa+tP7wL5s3QRS+I0QvjlubTf7hMMSVNL7EIEC+Wgbz6KCVKke9SLrjHEj0V2S
c1Tw8a2G6luRAYSd8suFyxT7z0uzCe/74x18+GFmKlP2CZ5Q6LZ3L+K2GW5r3R070m/umC/9dQdH
sDnzzJXl84dXjNZQOs8+k7PjTgM61Zaxg8lyl7M1n6wadjbVfeThqR06twai6PeP06i7ZHqPOfty
Tz7TWKkbAagt9WM3uG0c6UPAC68FSK3kiKDy8z3j0Um2Kk2aPJD2MfSs0UUhy/WHbMmK8KiRMhQP
qcUDO0ag9nJs1PTKZ8xPSiH00y5yxlbWanjShYbjW/NkbwYfn0JuT1oSBZE5FkxMMrKo8PahzqAA
TqDGPkZyXb6ugjmSWnpMmjRy2plUkVZ0QaIgZga9zvqkwoaeJaRHw8RAdPLKzwP+KQOxzxGN9dGr
WhpNsUYozh8NXFi16fyewdaCOVJszmsUXm0Q4eHqx51mktoF/v24T2c2SySiHaY9RSO25mgOjUY1
5rOZDmIaWgI2tm6Pl6Zzt2hWoHorRwqaejYvMgl3YDtfyU8ewvpPJ/96oUy6Pc/pmc+1ACPhguRd
z7hV0pLVWPkq6xJgTJIqNbjZ95YqExBxx0kNleGp0u1ijnZhx5zeLZg9EEqlaHCEt+yMudldZlkl
Jh6WpcL0oxjimrsyim4QF110rwrdWg3fm481U2UDeZ7YZOEvR8HHafjRyhPmAD3rmJ1Lqwo7BJ3v
iJbYQZPgGTu9J6b/7n2+wHWKelrevw7/JKjfknLyIfFq8tI5rfIkqnf7nE6Xc1gGBPbTmQEf/RHX
N5MwUNhXfludLr1k8VXqaUh0f+5cZE+4prYgOg22wuu3vM6zF+EaSLkcwu3VEO5cSKLFkvO18BL6
zK4YLlcW85ch8h8bq5LBtEjBvskL4sxxgze2VBHeKIvOq/eUJJ/nLwn8KQ6rikaUX0q7auz7Qi2t
hT9UPMvP0tKMhZQu3mSMOle6axZh0KwQu8nF1+uWEFozlKHjNPBGTIxTl2ppB3Xlg6S7ve7X3ZGg
fGvH8UEhdqfJ1pY959SjSxSNuTZ49NtmC1gzBRW4ruHIHrDeEg2MPc8DVHyC6GAG/RPsKJCuWDGC
qzqxtRgnydSkpfDhvqbWLTe97/my7T9FtglJDCDa8lubbLRZ8ojpOUhqs8/OzIJF03Fb8meMqLb6
AtIoGTp7lvSniwiK85PENPzCJu/0wzZtFdt7EMyjQsAOVkDBjJmhhtVSyWj7rJEi3hUEuMEZURi3
2hXBmmrN0TXieh5v1sH0NU17S4d9H64hjI4hv3MHwL2AJ8ZbBw0WOpEVYJqO5zgqzF6UgnvMSk0K
iVzW7k8MbQ3UAl3qL9SqfipKemJAROdpyFfDHg+cSPwxcVdmdoe/vSfMgbnfEWD2NEfrvKNBKLpu
lt98rZyMdgNBnKhP/GqGdv2ZgegDKf1FtPUdnPXSMeCdov0LCnudPJccP/9XZulmdvtUlzva4L3W
WW0rRoLS5pFdHr4CCW+ecMdFFWZUR0h3GQJXIYbdVu6LyaKleby8cwk/VDRvR/L8RY32lHJGClBX
EcMC8DPtL5iRgZ+weMf8W2ypHILafMbMB9FhOZyItszoMnwSs7uATU0VyB5XMsjpO8IFvFEcCdxA
wsHoVS/JUEmEtm5XcjaCngMiNF+3+wc1sYDVpNNV/k7wEKrhwvIRUPr8laNaI42ihNmAzMmemYnr
45Vh6uuwRjA/TDqZRnASdo262a2ObMtmnSfNT6ek8kRG5BZrPgmD+57L+hF9aQ1FJ5fVJbiEexDr
L6U4Q/IiLKCtzrgh/3H6QQ16KbC+L0huaP/a5JTJFnl3rLm8kHPKHrNv/Lx9NYwe4jTivRxcODU/
4G0AZ+KdZD0021J8liZgKuy9Cduda6bYAyygfkSItP89vAlMY/eJZi3HntcLSocO6r1ASyHsY6D6
Ec8l9s9kEvzM87Lx3N+iU7yV7wdpvRdMl9vbGueTKYcUIJKxxtA8LZ5ooDRAcik2cP5UB24RIdHG
FyRitgfG/JWE4n3bqrlYRYARnMzLqvfXvWl45sMSpgBK2uSyOPUgKB+6ndX3cfqgQyzYGt3+tXI/
D2XpuZJm2+KSZRvRKfKnPQriTyj/cDnS7Eippzjdwi76aqHgcJJv6HZDaXV3Gq13wyRW8rNelVri
hKQQsVRmssdhiZF4Ym0PFXO3mR0ZpVqQkfMJO9D/rGU+twI81oTojj6bD75zPVQM09FzFgpKt5Vy
yWEw2BKYqkqfO+MYWP2OSxvb7E1T9XI5ymOheDioRXAtexR7u6zE4NBOFNwbFUAUII6c9/F2w5ZY
8jNT6urR/VflluWyk8YYyHfd5xoxMMwvM+WkAg5qXstFbHBoyikG0qcf/n4UBwLvI4hH9gAkrrdf
KSzjPnwSihQJGotbKq0iXNYLoRqEhv9zVz9bum9rRBNxkrXnBE3VMp+UtN1PQbETncZiId8XVacU
iq7jTJUpvk8XFeNYU2bidwNmWY9t7KgNpxp8u7wOrFm5IYqvzrIcSeXvd70VdIvCrIbJkQByxzuV
yyZzlL0pAlksKe4+LK3mytuCDpU15EGVs3siNSJ+K6RJ0jsvqbBqbnH1oFyB04JskrTQW2VYjfh4
qR+xQpJyVlAyBTFR/FuxRCyf1mxMQCIBx/nuB0o6EuGXknijQ/f3oNre8oPLLaw/miOvkv43GtT8
7jJ34XxsPscfbZKn6vs6/rs2xG7HUBpIJXFI28kpXGnChL4EG2qSxGIy3srKTIK1rCKyn5bxm5gl
lyX69zOA6jf8276UituSXwgNE8nnXLrV1sZYBBOggbvcfAGrwPk298PwDmP9YSbIp7BEdwfRK7xG
OlpsGzVuemK/lPzWUc4OfVUuUZgckvvo8ETj9vFiYlTe0YzCmWn86Wm2tVHgLNH/BADdW0M5fyka
9OdzhtamXrGNBPaXggy6zUriD8vMFuspid6XzYJn6TK/S5+aM9DLFir6Jx35SWC/1POGvaJlgogT
sTlYALOKnns0Plqx9cYcyvf+3BpZtERuQJo52k0g4GD4vRvk5CFMPz45fH093KKoiMBP3S3h7Dql
enYV+slC3i2nv1SG4Do7D318yAPdpGoLFW6eNuH4WkzqP7V74FDWayBlBokZ51Pb/n7FPBbnNwjK
yi8foCeXyId9L72pbcP+g9ezFK3sQ3gOWAKYsL1/LPiSJUXL9w0WJK+7MjxiPdbLZa/LfToCwwyT
jHIXLcM9npFZrDcySww4u13qlHWHtbrkJMOD+yOt4CG5d81yx5q5gqo1dFRq3uHJUUUjrno1ZVbZ
2uG9tCAoA8wZWhcVrVltyMVNR42w6ycjLdEBUsSbuu1NL4uPquEeZd5rzXMGg2hpy/OWQ/c1Qykm
PK5d6Y1sKWs70/+ZjQBYSJjC9glRnd+YLCRK1DEw9riieMdccu3cn+UcADpcbvlorLP/5ZBU4vOc
3m5UMba8ZfZfMl5gpTVp1IJ6YtvahV9eQr/9yetXbPf/mhtatCI63Nb327b3/uvKp8Zm7Os+ZUfF
9yqroEDKvkkw5Xv/d3wuCwATkSNfsGoK6wtuyoWU0fV3fls10UZqxMQT55v/F6450Me57vi6CiSB
SpT8PXC36KcPqjPMAWljbVjC7fGP+hycmV/eCA8zZG/2eOiB6DUOvm1buVugECedVWMuSyyuJ7p8
mmU6WgrkgaMm0g+IfXC+oWMA8c63Jz6Jy248BYmASCQFQsJvDUuU71eoDhE57tQWF2kQp2bOjj5h
hwGwvrTuslYrsaOLKmbWUyXyKmh5R5Fo2fk8nTSi3Y8mBCb4N9VVWI/XlruFIlVQwJm/ozEyqKNi
mGTXugICnMrncTHvxTtb/1qReaGcsiZ21F0dr4VG8U3YSFQG5MyyyAb7EMoXHn+zcVjBtOLVe5oO
BttrYV6TTpl7Osit9ZVOMuM3AZwvjUq/oYLIME7o1ZZlep7uaM964zpdIloFAS6E+Sf/zYI1mCoi
GdqET3XLSI/PftAzeTztRGTQKVmgVEHoICM+6k96QFmrLiYAPBxySBO7sSMqzR80bejhUZiT2TL7
sSvATXZEid3YrnFMaas1hvIUWrdpMRbtSs3+8weqZVRlC25MPKyv/X/rdFMt5jwwPQAMZkCujLln
gAB0olDAx4Gc6dvfr/D67bbmCxHT+Ak3/cXRwbmYu52xcf9i5K07xZNtHo1RVlyLF6wEfpsp5/4D
FH4m5eNU0/UckaDwws+vkvtjdI30jsFGKq0QAVE2sQVmOzbRf4VbYuRqkLOk8OPpZsOCFYF2n7I+
aN9W0rEL0LEvvkIb0EJw9OUb1bfvsiYqYrg+o+OVhoczXNCiOGz0MpZoPOC2/zWavvqltr+pGOQq
92AiACqMt5uBDaqGLEo2voDkUjViaWEtHeAlkO2eKlccBrPyOlolS3Gwj/Q1PqbYOJ3fS1cqizqk
rZv65K9zA1XgIhcvU9idR15e+FYUWuHRGZzy0/q4db3128sel6WZiN1gCETgaN84Y3HgtEjT8c91
DuyRU9sCegNmyKXvdmaJ59vaALnNn/a0MpC2F0lM6J4WjZBBokhgCKkXr7wdeb3LgQTtgU5Cdd2U
dJygf4WIxX2bP36HwtXJA6vBaquFyB8ZzvPZ4Qw9e2kojjgbojpKeejX1gPL8lHtfPM+mSQIL0WP
MQWJcDBzUqWzKIEddmDBiQlwB50rt06g510Q4KgKQtxixTrvgUl7WlQtX1ygphScKFn2MZzuwr3q
OFKuajzpZMRIU4BOVlnReMDGWL5qog8QzXP6Yc4ibaV4i6EJfzE+XBidt2j0zUEBG5b8x96S3kC9
3eACONmPUOYrvy5GRq4apdVLxWrF4Bty8a2sahzLESC2VJS6PL0JrVwgYCoY9NUJggUSwJ3X+afp
PkCyp2LhGxxW/4RcI71MoOB3OUOsGAuhMlttbxw/td7e6eVBoeSybFTYLVAd74wSw0rlkWMWpeOg
WRoSZozra0bnEnjuqe9lezw4O9K4oJK6L/rPqdwcZnsSDsgG4FSEoZXCvKtGcntGePPdsXPuKIxP
ofv6rX5adVu/EoGadMGBqESbl1Chcmktn3EI24smDS0w4rxiKKmuS4eGJdlRf/7xzLojVU6oR1LK
cT5d80WMralxcvah6m/pPnp6lOVQbehTqymMcof437qAi9saFA7uqvBCdpNXJlX0zklfqu8v8gQD
lL4uHKoW3s7mrlzAoOWj6po32Sj7355sQFcKhJmjlAugIwOaXQhWybSLLKjUPtpoWft1Ivkqgnhf
T1ueTaH9vzlbU8ffFmEUTIZVql/cPqhwtfcauf8G8MgquGlCQkc+Hou4z40fqvl5Ij/1Ksr/9Zlr
+XJp503b0iMzKkZQrnQa61vKURifQ3FFnv7i4miqILwhyQbwJEATtzXQnYEZbL+yaeNtW8D3teFC
IoxqXEWY02z/f7iRkjZTlkGlwmpbLK/f8qBnbXiWWNWPOB3WQhEiRjWYSkIjg1csT4VY1BPRRq4p
mHLx8MKmSGveWgHg7AkwzRp9lkeSz/uPuiGAByJLLgJWLz7Uu/brcrHOS8MUNIiNLFD5ib2vEsln
RlLRKnQFiuTCK398zWiRwn8E1uVnJOLhWO5a/Pz+LYgvLmqXFxnJz3u1wN28rjjQtT+o+OBQFLpP
EoC1pxpk9Ohi4yJmjG8XDLZQkZ2dYwHqtqsdCpb2I/ScXKK9qOg7eyT2KGsMyAYno6Ge8l1kZpCY
zLNwQiQXuVZr1H2cDc0reM5W93alzmT54VOyTys8Haz+4rKhXh9vWhPnNN7DZWNQiyIurwViJQUp
P3/sgijvcsySx9U8fBwNnFZof8IhTZwGm9nelZgYF+e04O23ByiCGyzRaVSgKOSZ/4i3Ca4cgg2T
bjxJYk6MtYxc/MWA9nodPvm8cxlQoVJMhF9AKWGFAcKExMIN9SJ2hHY8Q0aU0NvCv1DlbT1gpOfi
60ms51odH74dIGl90fbEgSMcBOsNNafK2hsVnmeYO6EvdnmE+d63yEebxhtjijNWFYPaL4UuH1ip
b2xwfCCbvZrjQoPg4uKUFhJW/M2GN0Op5JVBZeBn91O9J+SgPV0jCgdDBVk0uuXiC0hqjoWhlQX6
TaylqmsKCtEGsH5eilRJ4f70BYkEt9rdMHApr/E5sXo3n+91QuwMOSoQCBEjaVRIXMvKJEvsesOw
+68bGzxv1XYd6XETTrXTTadIzSmuhwQJGXY/82TDYXgjiC6hJJtQwUo+YpLKqNpLxZLconEOduJ/
KNTNv85mnjpIG921IjAoOF1DtSNphrq5zrk6lyLC1Xqg1lbeIg8rwP46zP4GSk4/Wd28QXG/+jR0
tI8LfcGoXl5f0YO2arKmidhODFodXEwNroB/X4Z7KE4E7FUstgPVdeXj3sWlOvcnZ/2x4XaUwjlO
4e20ksyj0Bcqu6iB4Ld+IVf1ZG50LyoCRpQiXqv9ex9g9HYkuIGaqkFvlyhwyWtUIaLP3X/bKsHB
1GLDzpxkqWiFhn13TFKjYUErgPcMzoD4xJ3tzJcpcdj1GtpLcHZOo2lIdZaviJc9mqw3KiCgmMCP
ZXcXeSwAV1c5E83A6waxSj/Nk8s+HNsWRkBs8OiM1gM8qKHrAaEDFkNoSo0EB69YEEQ+45os3wYB
ySmD4SrhsC0yUYfggGQcoeDcXEyP94GPMCWBqJKfjEscGQZCi4Nztg2jwLQZ4Ts7UaCgKn4xSscK
VRaFCVeik6/hrTgRogg9AP43H0825NQ7OW9c4kLi+g5C4yPOcOel6GaWFApijx4Zyekt3Q7u8dMD
3lKnI5+FBecni68vugLmgG4dod150060ggRRCLH/oRVnmOX/yew89x0hSnAjuEkKhdHoq0j6beyw
HU+o1KIlkurF67I1JZb8IaHIlGY+YmcQsVeTTMqtJPS52BWnm9DlNXZHjqg54uFNrmfqfA/b0KB3
o0GNqr/Ta1yzewTpO4NZ7iSx1Jg/zLQQVCb20lfFQqAeGRnDBbWor+zrr4rL+Q8oDx/NCZozTTty
l8PXzh8ltmBclAJbuA9aVCEXjI3yHDt6xuq7cXrI2k/BLv/b4St0lc2xxmlGcT5khBG3oetja6zA
tZ5q1ium0EhOuybO60ebjZO4mjbCYSiJywaNpqAhxiQVkwZ4aHarOoSDbbRJKK7MAdEMobCSneSq
5Rk4Fh2GlK7FvOR9JP/9cAuYiEs3wVYoQveXVD7uL5L6V1fnAQAJ1hfBL7SIFUr8I6cS193XV/zb
Zr4KU8hhJrjE5aT26l3cpd0vLhD9Ciaa+Txiq2oGnLnbCoLRXqzS7SUh+Kudhab3W5RutUf4QsJV
viFbUH7ljGSs6P+dSe55w7f0yLH5rMs/109OXxnkmESfsYspU/3A+tTXNohx5L20Qrbm1q2UfMd7
AhGXQxfHnX9/7p60yop7b2I+2Cquw9ZFyG4F1DuyIbYQA3/FuZyQQ3S+i/gxxJHa7nGm593AXYQI
yZYK6p1yZQih6TwTINZnw/6YQovu2So7yh1sWps2vr24D7N0DiHPHonbROL31JlQ9Bnf737UPESf
UZpqQzAyZ3Y8aX55YBwlc3wLYMTBmf5cRlPuInnALqYrmxG97uWfuI4Z+3vHTUdRLMiu/zjmobXM
1kbYnLX4mwVu+SyYOQMYcj8YjYX0axmRVXAnIdtWEC2YUs/9gvi2D/rE1KVDIJ/8ZhyvmmpbCK9u
V+lCXTZfOt+/OwJ7VRER7/89av+gDC4r0saGSWWcJobJ0I2yi3/yb6Ce7eM3CKaMQvUj+KeKn2aN
b0RH/Uj/y8gdorAuEHWOhHWPZ6rYP88/7RTBCKHnhw1QF/3fiSefGdyoBkZr36laiziutvW13WK+
4r7d0WAEXNbsTYCIbH0f2c0ZCW0ZXLCpBNxLJjMcyJlQWKlh9li8CPl6YDt+qsvXAf7+Pbc6rTzx
coXRs7O7a/GbP5oP9OhtZ0WWXW+7EvSfZ3lbF1UJbpNOjA2B5KLWezvM02bi0U7qJBrk8Xa+ibSM
udsc2MANyo+30SXXfEeh+SM53X3Ht9eiYRzBZ2dXad8ExqBZA83evd07ijMsieIaQrPLh/ajNB/6
t0MbCPr67W5BFx8wMV8RUNdJI0TbXV4dwv/PrSDmnw3TEBaofF7LU2Id37QN7FeNDc4g73YC/Zgd
zEFG1vkY4n1KFtEiN70vGhHW3tugyE4S8t0SoxVfRFlZD6XAoXmU6VtLmta3YRGdqAOBnXbfTZJ1
jl0pC6XIogizmk9hKenJNxD57INZ6xt7pAg7pKnn/BY+30b/YQcUAkWenvWBIOEI6h9BjWQ8E+HQ
gQR1jthc/dt6zM/6uAnmJbicTV2OlCXYJ48REZxxI9UUw1yUKtutH2wWt6ZV6coozrBxZwX/utXR
nHyZDaTAJ1qY/mxeL0SJLWJXHiRQIEijkSK1XwyKE2xcyfhG5LgpfZ84fWV1njre/A2UD5txMWoG
QLGXCO4seucNxB+zELxjApjSqXmiKpqqg4dchRu2x35In6SXg/r03k49UQubk+AlbsG2MJgxGKFJ
YdWdzFtcN3wRMcJQjLJ3r8M+svE89bmFchvK/y5Qc4nTmuGalyd6Xi4JvXj7rHwF6cDWItdrYEfQ
EgybBsU+HHpuwZxXt16SDRZXTER9mMa1EiewNKxXZnIeDjUsLyhiPXBYOIb+vNx+11OQhXaNoaQZ
PFEvAmDJVo5i1wwKHcWnsukWW2E0dQ370K0CF5IZgm8iQeLVHUtpAdBMQMT4owq+eglReB8OTiux
u7lIdrrHee4aDfKvoBdou+z0xk0jd3xKIypmLH9cS0tUjGO2VeTCse8bZO5ya/ZsFcdBmEv4zrz1
tNykBq2UxkHTZ4PYueVWVrn3TVIgBtekYJyD03VxKqBi/HO9R/taifG06WcMu7j6ZpAJakaYSfwk
/9rzxH8dW4EV972EMIeEFYqUhlueq8PwVE+HgyE4pgy5bfZD6tTPy1VXPgM6NDYskVg0epq/ARXi
iZrdvqfeX8JhR05SHi0vVOJSXVEjuLcAGiwUPM2K5MhnFQKbAQfl4LApukBiATpxLxmrOeqFpLie
KcNUkdAZxNlPk4DgVc2uDmhIwejfaMzo9n7AtNXczgNwumPiMVSQdLZ93sKUz4RGzCry/h6GOIzY
vWbCKnV/XJRoawxZ5xLVBDTyfmsQRQ184gQtV8lEhz4/MiDWM3Dh5zpHVjO0Id2TOlIqe9ItyJKy
lZFq5df+43dZw9Px1g9/nJmm+ZEDLCYKpVC3oVEVWX+C/NR0tNHrnjQc6u2E5YNRhE1h1SlvYGNG
UA5NPSTQRwLK3yfrrbVF2P+5aWggSobgwJdrBv2zIYLo/5wVFjGZ3Ykc9Am1xK4YmANumaSyA0vY
Iu/mO6yP+ORbxbEuZj2mTB/rt+W6Jpi+KKijs1ZMU6GUUcNURADWFzk0QKErOctUMVaO0AYKGVrP
2wnRJhS+7fSrIPiV+QDTUnSIMvGQh7SjAfBHNcifzp5TvQ8Wnvwa9k8MHn2hpEzF/uV2ZB+YW7Z/
o9GohHXOOWMdnnOLyDC4aq/R03Z4xZtwBKf3CBlG81HEShxO5h3lvTfliEas4tDZ27/UUuveDe/o
6TPbUn3hJwucUlrQkTlfvmavJMvklEiqqsOUaYM51KFzsMSuTmk8nxkrgib/Urh09aTh73oLnIJF
PCSEUfbQensApwhx+pzafaM07+xkpaXGPK5SyeEMu6SZLw5xyBMaN2ARZkv/SWs9NpOhMz85H/xf
GHbm/U3N7adeG02K04b204YjMOW3SWb+Mo7tE1jASnAJ0XMTD1uSzN8imsNMT26clE3hjKtblGca
n0Ph8ywODkDO/6SAzKOZ/AWkbviKueA6vMJOyb6NG1MIUj8LEueIdNLV06swm2C32XbBqx7GnAWf
Fb5evr9h0WtqS1nCcBR05/9EsQrqzkgZjYbLiDCovNVr6CS91VtgKy6XfByV2WH6bk04T4yNNfRJ
ao6o4CX91uD6AAYhoOt4/g5EDNwfEWcr2PIZ2hw+VhOFr2THYcx6yfykiDxVxissTi3LdCKxNc2q
d+DUcnc7BniBt9/5a2WopQ7GLeHvzTxJXHUufebqqBDpHlKOpeOWfavYAhwI5nv37r2WuoL7D3vQ
QP2Yz1b2vNYyj0hpQBf/KH4tjpVPRnRdJ/Mcobj+GlQ159JfLonzihUDd3D0ubyVhPXQXh+bGByX
i+D6Hu4T1brjagWKQtCR6zGK8pRhYUax3vf62CyI9TLRQe4YVSjosfTlDZF5okaoYN80PtGXtlS+
WP6DgJZ9p4piWox52ZMIfX5a52QL4/2cL4bHqyDj+YWmTd4e6qSmAJ/LYvwvdTJvEqIUEIfTdAoJ
VcGrPNVTm8LWPkEnFTYhPrEFYBtwMxD/GhVMAdgYcKvaS2hF77GInLH24x7sfnE5vg60ZSQmVPKM
ZKfJ1H0k8zGneOTCTbmLLUSrE5+w/aKrSsMOLDaPO/V0mD6rI15OlOnhc2r1xJ8U4kCzqBHkktJL
TxjU5AdhuXOpg4Mvtcflbo/JcZQJaqBMa30e8qGzXQrY0zJjLLvpeU0c01PhYyKw23zkkLnTFSZz
LhJW7sJKlJJAy3lw7xuTvpaHWCuVgQIxstAnQr1WHwf1sOFP/kMZH4yekSuccotFqpaKNRBFXEKX
fGjiTAfuv68nrJGPS9LJm0wUK7MvM5wDTOGa/123WqzMLouoKouiA1NxYwtj7bOsCivahMonTCNb
nSddQHmEEuhm6er+I5E7pKhx87qGWU7tpeAbmPbCsgSVwKtDOPADWfEwqsAxQgF8Dft9d+8+L0D6
8u1c3XwIkcX10pUJjV0+erzCNHWmMU/pP0xQTFaeqpKok+bx6B/okyeYo5Nb4jieBX117rttzRRc
5OJIdyybNNjxGeGA1xvPvPEapaJBeiroII1cIikob7LE6LYMQZLvjHeb3IhlVBkUHKmeANjn2/0H
gCMRilTinac5PTm04sw2sWlBEMgGbc1cVDOqNNLdl7nKZrNiNMuD2fQQLfJ5oqV7Vb+jGOrZsPlt
GCJL1Z1qf82eDBFlJ+KCfzhIjv5Xq+1yz/97JhXl3HvREZ7hQht3q6P2zAo48YOmek9xKZyBS/vj
2kAOgKnfaqqr42EunOZgLrto+CLaQJnIN6TrYlfo0lIyIfGbM8umpXkApsD1JTF/Hsmxe5gvAJW4
yrZq/n3CZ9fLSZV+tKde3Wskowe2oWMQM5qbXXvXsXEE6i85CQdcXp/sN0NSxHRb2sbsOoVXL2ch
M7V9qee9sGLn8AySoEJdKsEzelf2AiwNW9AHQSACHKIr5wCKs1NOxe5ZWal1z+6hqDJ2/iYYWpgY
JDFNRyR+yj8f+we0t4JEwl4dcpDvbly1J83tchUw7BGiXUERTw81KoPz9Yh5oUwiz0iydAuRF+kI
jq7/5rDFgIij/BmtpPBtz3r7WCzbu2fxJ202cteiXGDbSIsLqaKIQ1Wcdyjq6ppBkrKauSQJtPl6
FJ+v4sR5Oxhn8SjoTahZAI/NQGf+qQ4nR1i52eUFqZrspeAWSPCgoLAukPxBZbXMXnfM8BT+rI6z
FDTkQ0vSAiHmzs6Moo8h0D3pggtBvalxrtMZlCQeQwqkwDkGjyZxSyI17W7lkQXtTa8I7tG3DOBL
wCMHWpou8yc8004zDLAJUBtPjk2mukw6yIcE0HAoaBWDn1bmrYdwTiMbvXSPyKesgrJz1wvufJCx
jvDA7XR4+r+7oizKIGLu/rmeP0kb6xo3VkJ057/4BtUrsrcYhjCcl3qxaklvhzLBUIAUq0nQblpG
SUr7SvnkCZtLbwxdbX9w/hF0sdahRqoJBt21GVTEEznZ2z7onTNbKc/wcZW5J1ZvcGULdrvnheQp
buSpnMOvySIyo7fq948YhtdC+OC+WbdgJ/Lz8tEZ+linMNFxX8lxSHWoOQ+JegPCXqIv1EZNyXTj
98HqmUkNUyLHneWYZFCYkyVivbMLYNNqDWaogqzfgHsqbzBmxOtc//+jDJ8NkULrV4KfxaeaJPE0
v8yYl7bsp9fWj72ruJirAgAT0Yv262Dz55hzMuIQDKTB59IIApw5RuJCdjeDAc1QMllzyELwSmSR
lr6IQd9ENPeopmeegPIDiRKPafo5dtyGji6iiIE+OSSvh0Bb4BTO4Nm1rNDCAh021jyJwLOPSUfl
Hdjl72KYH22Q4/jyK03XNqX8YoEbFIJyAsWsZQp2yiHTEVGOW0a5qR21+zMe6hpbZpaBNH71Zb2t
xc2p1Kk1zzabEDnQprgAHMEIa3RLbWTBQaMZ54tam4Gr0mOKp2N83T06FmArAsnYVqWj8LbiTMm5
u1a2r/2VHivd/3h1GHRBmFUaJ20FT2h4gDlu+vZS+aL/UP20Vb7eKRVJLEQNjSO2+R00wMuNik3a
whgix5HVlR/dDmMNDm8GJPyDrdPcWtYDd5qHI4Pqcj2kRabl7HHh8GT9qqseggOZ32wV8OQpliHT
b01FiAeWfjxtwEB+sVDsDXskZt1kR3Bv6Ux+K1XaLEWFtjDZsOEvqrLs+Q4/zuLvTMTFVmFkcG4g
YxHRP1OxkjQRQR0QFSYK7kJ78YrntWNp/A0/wOCfHNzQG9ggy3Wxp6iS9dAXcxgBOS9vyvUblmdu
OAP2pYm+Jp70nyha/0SlA0+JrLMRoTbDQfDuNTW6BBN8ZHi77/hR7/oEom3TlTiLez9MQD+XvaOy
ZU1gknW0EPDwDbeENTP94oHqja/cSgG3yhuBF0D2815Jzgd1vBb4XiahAcK3Zu/vsiU99XRfIJxH
b3oLe930uvLTrEdAoPwGZEjCceCOAk2J0xcuRaoJQlEVFQwjFSMS8/zof1FmEk5tzIpwBTLGd7kx
zQv5H5VpXGd7qX95B5jiRlSWdUH0d0no4mDCY+3YuicEusmndqxso25VFNUvPjst6Hy8HI142zRx
IgsG451srFaakRf6RJ2kupjCbne4jKUz8bMfW3dmvbmDzWOMhMP3BOfizHeVmd0Osu1OKsGaXDHA
axskEn9Kg4dgMRNhCabXbaSgVaray3va9ABS4slm160wSvPsVJIrFvJqxkzKkTVjHmuQOwjyIZbv
4nGgFOlk3diDXQb128l7S2wQyxDCYe3i3wNMqo/3qFin6Ar++WTPOGqFUbdZZoxXFUu+a6xLY3E2
5+FOZPCZxN7C+v83cnvkOWCVaJEQQyAgZiFLpN77lje+gIFFh4hduRTM3p98+nbN/Unm+dHxSoyt
CnA5it5r7nOPA0mv/bPD9n5JRfr3soZk3YmTXqymfAFYoO6OCh0RZXZkSvttQdsYg1KHUsB8+vKk
/zacmCk0AMpfp+CuV5zF4zbnkKqzO1GLcrB3gRfIhcodHSdwpWlKnoZEjbnDBxa12Zj1RgJ6bT5q
Jg0FZXNfFTJ29ZWyfRsKrvGZ8KBD6kRhR/+JcjwJzDTJAVeqjIkMRnymWDY1xX6ECCSu5kBXhfyK
jRVgpdagUX58CM/R8lETXkqdT7iZStMXm9jQrdXWvLX2Cu1T3/Iv+oIJNwItuIffEJU+HsyJ4sgv
/jBHwHzlO6TGRsayrT/TZkKkN26MzIQmzndWKb9Kg4NaFeyuOPh8Dqcr+WYWf+v2PQDPUXieP4K7
tm8OZeU6qeoDY92Ig0nIUbog6JCTtyUrkz34M67r+PzfYtNhc1anvzfc6YFBwT+nLEnTOMooH8FO
Mq1DkHg44E111S9V7ClwCXle/AnREI8POGddMtQxuG8LPqSmLZcLVVLGt5w7jzpKe97JCTQ7Hlh4
hJjsIQ+abRuahaczZkPtI2bbQsFyL/Ms2FJFBJhu7fSK/5zGi0ZqFwX+xTH/3UgLkght/W8PqNox
FuisB0zHo/CVRl8euzgSqbhdjOGfLpNciaqJTQhpQcCcItslTdU3f9v1VYUGhcSe2TSyyWC7Fn8l
EXXDItaQxsfM4hIeimMEkugszyNmtlkayeenM9BsS84OxJ1REmDvDaTRluXZ1uUmLJfk5Gfn2qIQ
t4JOenMSHNnfvV/9vumfe5yJOp08uVBQxYC4eIJ+SxYgKk71J0jIRM7U1FRUhCN5n6BYEix+FSGE
wQn0uy8ifgBDYvHUdWUw3GkuOaOliNf5GW00LdiKMu3akibIhN1GdcNlBUnS4bKM7+/t1tFo/8Ae
POJbg5RXUvElAJ1/r9yJaa1fLRNylnGMTowrLjYkyJiWRe8H36EagdTbJ+UINDkeC14JOmwY6j4b
6v/nUx/Wc5XxB3IXZKH5hg0WKkCWUR1e54s0LAnpe45y5thcDNxYCFuOfigDRafUnDW52eqXF0+u
swX7d3VdomilrkZofOg+jz8JAkEv+aBTd0WvBRxn7hTvIWp2eEnNELbEq1QkYd4dYFRwE1X5a6hW
3BNJEurMsR8J3RZwQlKjN7JsbQ+uWUxEWuHACNz5BRIudnos7pquMo1EgLpvhSLoMFgVJlz2kwz9
b+NC9bKSzvqg6qZ4h5skS+2PSQ8ibOWGffo6Gf6wfH3cZNnJ5wnm+lXuSJ29OVjv5yUp8HaREy+B
01ZyYM7Nb+RC3/PiXzUjomg9b5+Nk5xf+Mu9fbSTO81AtDOw1YgQknv5a8n1ezTnQ7xKp8d10ou1
WU0Bc6HqyqwchqtY7mdpg/nFAStgOM3c84Rb+SryQsLDwB4RA0H0K/fUTLdgBaSCxnTv41AauT40
Ky6zyjsBBTMIavUrDs7U7q4G2UNWzi8k4U9bspFTRZjp/Av9Cpx0IvL7f43v73gcwZXudF/Vl1gX
GQ/tTmM0QYFXK5GFulSfGQx4+fk2GA/iJR3QgT9XP0OiwEH/QtAbdcUcm6I75OFnOcu71aWwgyL1
M1ufgZ50ys9gzUWbaWpDWT+gdP1ZYyLSXh+1JIhVJTxMt1yT04SGPlV4FELClJmac5u1xAKSKEnR
LLhIB2n2TMVIwULFhiYpKMhThnyg+g/6YSymbJOcn24iVcdyHTi+GkuCBMbmhU41NPTmMW4RWGxY
N4z98AonQNl/uaai6wTcjLA1nPIa7D41gWCqsJNfeoGBRVo73nVTm9IeEgAhCPfdym0UtFxxyUfK
82gfyzFLbq1wK8MhaqeCz2GmU454/z/TzUOxOqwCsLPKCrdZN0Uvm3oex+YgpHVJQEQSXCXct6Vp
FqdfKFRGLUrORFUHUzfQEkNe0yH/5bjQeFzvAW9mOD2FO0qO5kwfrbEl7IMHhn0TF1y67mN5zwd+
JpAT3lSVLwoD2+p2u/dzbUVC3DawmUEqtjirSvTtEKcqaaFWK9Hise7eDrnI/lxVOr9cWj8n4n+r
lLEsTCAaNUB7egRiWZKWycVZt1pKODdZJaIep7tjE/KheCCMJ+q9eoFH3H41PRGdjXHFxY/RwbIM
Etw1R7TQZNaRd6C5Gs4dSRxn/+n/f1podNMrmoAtRB7WvqYP9dNRnPDinuaVCa9RKj0SChiecfaY
G6HWprX77XEHubfnHd93D9CDJ9+c40v0rSMt42cDlfMzAsr/iGXGaAurkJSEho5zZ1l75SwahMZZ
iLdlG0z3n2+EXCtbJFojWPIldBVo/jue8fgQ790umNOepiCIGvnZkHMKarFqK7k6eo+BFzEWGbVc
nG8DJS+unzHCFFZDyiydaxSMsvv7Y0Ui6sSsBMLeKv8iHt3cEStsFlmr5ECN3vqJjrFEee1sCO0b
FE9XztOcizNjKBgA2zUI3xrrq+hcZ9wBupCFDnvoF5XI/U9gqo1CtG+MvtG2WEZfBGzdfZjK36g0
T7/BHg2ednq1+aefMe4GvxgWpQ/5leSgjrvGUqgI+yTXBNoaypyOYJvFshUfNjpB7z9OppiHedw3
PKD6f8uVSEOtF+oE/bNIPdZabx1pau2OKKmNltTmw0Ybw8dBG5J0MI7LfG3gByPACeVeXFJNzfxf
OlBLccdX/uC3x53NYeofh2MDKsHCOVtTwD9XqIu1EM7X2YmyaqXVqKu03J0qpdSLOv3+Oh5KNXPy
wCAw7JxbfsSKBc9rWCEFb5IBwyFXNRXGuhoc87S7U30myZ0t33qvsi1rNWfUtvlr1SGS183Qtcy7
v1cnB27zmIkuJFf9Co3X61BTmrCW/4hhOajEAp1fsyEZarN29SUIAVvmExr93cfulMLa6eFDPz8R
EmkGFgee/ugqr71bVVKLp4KpMgwOd3JyATFQ5hzJmU6fYlJT/93+ypvvSVV9Icm6bGpTiSPMeeQ+
z/7BAGKrI1h644/NWS0q8JOYkFbl8QDtnUE4LMMsKdB5ovlxQ0PpcYrW6b1ULd2qgIdVXrZLQxaf
3kQAoIy4oLY9H8s4IDrdBIS9+N7yCA0ufB917tDHm/mL6MZSe+4lBl90nh8hGvogNnJQqJ1f9Btn
amry57ow1wJ53k3BGkpUQKzvf9oW+Rg9WBAwpgq9HZULgnCnfr7vJtNzGO1vwox4QQiXWNX4GmmO
hfto7hwVttPGeyqJ3N/uu3YWljz6ujiZAbdRtKkdu5tkAu6FEranJntcNBgAXpHNu+BPo0Z5JOEz
1FobWzjdH2I4Hd4xvAjpaiO3W1k5jY8QHWIILcVQ2fJ7VjD4pQb3NuFWAmDeXi7Fv6laGzbPjA9g
zJUa+uRn4N/n8LLjKXb+ChQITV7NCfsbpSayk0EQRzvF+MetzSinGGM0NsMy1ubxEBaBsnjbeCgJ
hyLC6BmbF/VO/rFInGJjtHIMXro50/Pli1fxlR2jEayrKj0ptEt2o0ioWALFto3UP3iCujgajOwb
OaqY+Obp2+JiXGqlgMFEUB8k3qLq6NBRmVCBu7Zd7sVQ3JEHlUGfNKrvXtmjSv/k6D+nNa3w7gK5
rVtlzouO459p1JI+trRKLRzvT3oadWaNMtuMPSC5GNlq7nzVsw3dnJidqC02/Z7XbOsZY3viwGzG
DxC+T8ktanta34md3Y4SZhvva78RrD3u7gpg2NixtgJjHDmlcdlCJqCU2gA+muU7Wuoee7PuLLBK
fBeY2PE7cAducijFtbU5W7qKw6IiO3y4Xt5M0KTgpiuqal9gY1LsG3sgGnFvwXaX3mzYEpK5VefH
8OeKaCcasHvh/vfAvMsPcME7oin8dQp6/v3vHuxzxKe3nXZ77kcKzk0JO8oKNRjArKPeFpRGFGkt
PaI+GPsmDhH6tpCyZmUeKni4VgZ84blFVmL4maNcWHKRv7Qan83GCwj6HaOMNWkayug8hJtIdgBW
RVO2LG/9SgXSyGHnSD/OvMcTb2qJg6d6ZBoZcoeAwnhQUJjc3vjelJ8Po4g/56A7go/3ZyJ9Px37
Qpvp74c6lVdVzNChL0we4Jl4SuhqRR8jFMa6aA5Hl6j11m/ZvQDpu3jmaNSsqic+Tz1jB1kIw40j
uy8PedCugQ5e/fCIqh7ONXs3fMsJytLSWQRls9L3Bnso7C5JdL1QlDK2b1YXy8OCYwXntff37Chq
EgO8Nf/cmsKpxLY5l8cMdgEDV+wiv7b3kVL5S2pfHmGu2GDPc1HEvvAicOmH36a9G8zzJy3SEBGU
3AJ4huQD/MPTg9We1MtplJ4eMP1LXyneRm7wYJxdVeybUriO+o0FP3hloN2iTdGV5Voxxuaduryd
dMCGZ7WMlLX9NA6Lgee7/wnbwfKCbGDK4IJReArRBJUKhaI4VM0cQh0hgYG76YkTsxmVVuHRioVf
rSJGv4ISJi8O7HGFnqHnfSxd/DKoJWfT61C2miEmTfAwF6OzoR/NUeScn5OLGHCZyS/S0p3/FZp5
6mHtdSY2wwMFYgH5oTfvuCv08iml/YBiNbNBDN52VlCkR4EMK0QbbxqV11UjHI11msxCqBekoP2w
aQCCYOIc9euZJIXSfmQ7mbxI4AxErZSY6upFw5AkmICetYya4sdTmeg4OLibml7ClZzw5C6sr826
I5F1tYRZ7MYPupN+1HfqEXm+K5geGr1cee7ek0XQ7aFKR5ypAaFSHGTRbfkzvOJBM3AZYyf2ocaK
KNJhxxGKB6ljTlnSwfHgjqPaMVBsJ5CIo3AenJHnZIl4DxTSDgbCLEn6sqe125v4tzs5dODROYrC
pc3rNlyT7P+f47CgjMpTZf1i+Y/kZvDPJy/IGnxZv8KcLuIJur++sF4IcRY/jFk34h5MyhNsQW72
DaUZkZsLvaOLVfdfCgzbE23BkQVhvazArgEt7oxZb6ZBHQz5IemwBkLdspmw/xNpsyh14J4d6Ndw
CVPm+csD5GTX9VAZQCJdV11RSTkyXOCVSyrhbdSJXWpj+/H5RpueIAEHE/fNxgVmG3+d0CN6TDaS
9FH51q3o0WkxpBoRwyVVngwcCzEdLh9no1VfRQ8b15TrYfhB4PJxVajEMP09FrTkFikVc0seK9F2
HOFN73kWkB+50H9d+JBk6U2FGqknWyy2Xbn7heDMsPq1T/ZVxtLHNx+yUd1vyk5SnSYAtBn3/e9Q
4VpAW0oPPEjtYbYThOuknZrHyqk7YSGWEsXjqd2blnqMnqXpJXBsVzL9XMoG89qExxLx6i58oAJ0
HDk24s2SPEDnOMZxpYrhWBUtvIi9PCJhgOSApTomaghlm+mgEyqdKmG+BU9n6FcntjOCPH/vghpe
4+nME3LUxvDqjwr3aYbxkUnBH3kevOOSuFCwedews4Wbxze6uJyvZoEf1VCF0EzLLrgNHgaNWiNT
bu7z4GZqz14gHwHlHEvCymWi++wN+AjQRY/B4fYNhVrAsqlwKi2NbQ/VTj1GuMwmMtJgc8Y2UlcB
XS6yq+HpDG3VXarjfzEakiObzD16sjSoHYu6JCDToiGEtMGKJ0CzvIxUPogpu5lyZoo4rnC7iIjq
4Ppgt8rBtUIXiihsoFMp9gNmHgazE6t5oYSRdOrnmKX87bc9g9X5Wia5IO1h4lq80LHTsFEBwLOt
YHHn7DddDOVpsA4CfLqbH24HMiLa+QqSu0YlJK+L1F5INXCQg1fKFSlAbaZHHvhq23BbuXTxNJwR
gxAeY9NIqmQ1QWkBksv/9fLjWpomUbcxiyJW8rK5MpeT3KNl2MMEW3eWvVAZh59q+qBXFrXDhyCJ
5Oq4UWn2vuZzdJlIKXK0NKioV5o77/LCLYayud3vwX0opegUfL84faYYi4gQn047/ssU625yi1p0
n7egRy0iYUEx5OCVLK4sJNZmd0dM4qLRYNG2zopCuJ/jvjbGCrtS6LQgRROxIF3rCT2Fprq65W9r
rrC6so9AXlT8QLmKVnrh+odtH2NEn1vREe5gxEvBxMKXCO5pMCciBDJU7dD3zwykqpY7921i+Znv
K/MjElEIneCEPSkmQqrFDIf4j1o1bvAp8+TxONdPSnbd7nVwi7Q1keji1JOaEOlEmbLBhz1eTpeW
p+xaf8y7fBpxEtouCNqhh6MdsZDEC+F5vP8yxBejDVyYTLSm3W5Vl9zxS1zsI4UE5M/33iTuOZvK
NvgDZrSnCQ1Yhw+ih0YdFe4iTZljKCRb2xXYgD1m2oguW813hvjhfZTOSc7Z051KkKyp8REHJ3k4
vngJG1SFoRWYU8K+iT5ql1f//4vvhdSeLohdPOw5soy9dvX1xWGTHb1Mij1W1nr7ifM0XGnYhPy7
sNrC+hfsFvtAMSgHL1h2Qm73pJO3ThAtbZl3cB/9MlDJbKqasQcr3nYTJyVDq7LmWY+Do1RCsU48
Wm7O+DXObXBTFVZz1b3jKz98CCIoyFQBpxjYePlYi+SvPGMXAt3Zz6gYNOLNg6MHOGnQX+xA+UyV
Mnx5vDbXdI6VD5rl/6mgwEuIQij1izMiRW8ZnQpYARZETPn0JWLgdBNKYesgrHeDVMz/48arz0Fp
QHk+14sH9o+s7nDg/E+usQ/P50XWDH4QSUkCTbQJEdLTfvbCEvkvUpF2hw1cWarvIsFnVsl9Xx4L
6GFmXbZEOitx5WevT5bsizgOmGSATwf3yT8xLVYlv6Hlwzny6Uj/lswSZ+JvGR9pRbIcCbHhVG87
GhUdZ1UPwSf6hj4ku4MzmyZYsAAP18an73ALqGO5Gc7YgLOv5GZrMN/vQBmISmrvnjohhjdcqux4
Ju7hT/LP9/y859BRtCOEKRAszjJWAHe4ZDb9g7mSUbbt0KhqGdbHABhI2nzv0FxIGqYFV+0UHAqD
PV/abjVQVDHzt6e+9a7eOqXmfkvfdioh3PO5S1Xs62KwrELUH+8xLzPyzqImuXGqvP/aEathk3hh
eE6DEG4YlLOneYtE6EqtqJpZDneDw5CmPQZqpgV+2Y7oi0Ie+2KLldxXFhKRiSKRKpQ5EOMQbrLE
wPSGotmVwC8RNIhq5mILJHD/ohV9o8d9Yhc+3yl/Ex7+Yu0XJwuLpCusN9UEcptlyTL0KdrzB4Yc
JWo/9YVgP0AG3Z+qkvP1zNJQ9FZIWXTKn9JtoLacqiEln0/wWhJ0B6q9259hKH4ByJnqQIRGddQ0
eoPUVGnnavGwIJTdjtjDZ2xy1NctZzcqd7Rt20S7p9VEWhuRNLbX2bh7C8m6PnYCl3ucFuAGM1u3
JBkAQWD/dcVz7ev7kE/APfkMHAj2f1qhNaoD24MeoDYfMSUNOkzT7rIViQxOlQl1kgbVaQ2nPjvo
3+E04EBqQz5C9k1zguRiVqgCsfhxZLgU7IVMyo9l4ohQVISpctXLoT0bYAhiU8s3aCCI9BrKSrqb
TUvFlregskh25yDJyBcu/MAWjTTOg4RbEoNoUHKOy7yo8bX5oYMv1or85+NqCz6U/yXN5QnGCtM6
wI0AD+DxKtAVeW5uApPLyCAIPsCldRJnXqF2F02RTlksC8zdef3mP6ZLSBeX5ZPTsqvzzm6O0Z2g
FRrP2GXHc1OyLHqPjjUe+4kDryZNpRdzgGHqjPhno8vxE84DZ/OpbUojhE5FOszhQ7t5mFElh06e
A26q3BrBcxEkc27d8kXPP6LwFCHBnST6RaauxsBLwXBBUsoZZtfs2UhyV6xyhmjaVeK63H4FiuFm
lNqtA/L4eoj8Mj7s5sN5UYl3xCUdYuZ1FxiEJ6EnjCnbYBawXY1dRA9BkqWKNqFNHL4snglTtGk5
dNCv9RLWUZwMZmlY2UI+H/0TD3U9vOyGCcArXmKy6g8GM9kDxixwL2ODmhHT/9tY6Hws3DobZPtl
wBV5lyvF5zv736XiYTZ9izeHCl62qtxVv1/Jhd0Lt3IL91+4hEQAF+ZHSXWbpAWB4g6cie1z0RCK
Qh+dK3tIOr2dK+1+YYwwoyR18QsMhQkWHOxDkQzS24agn6KoZtcluSzHgXYe99rPddlpnhkifR9j
+oJ8wcFCbnwHsQ/Mxhz+bsWgmFFyPZkzPsLd20yhXO3zUpYjaYolCErArXKT7nT7TTuMNPuGJeo+
KzoY95/DZAmPmm+KA2j+Ey2IZSzEjeUsW55qSbQ0ImxJbyO38rD/ERxO0xLbmyr0ssDKDto3Daa5
5XMNLJvEyOfPBKFgfuBZRYgssLXPB3lJO8c/ok7BqAzHe7MyXgZuOzhA6HunGwAMmMgfxU306bve
X7s7DZ5zcAxQAma2x/20kXmqgjtdHCCpNp8OQUgUDdC61ae1zP0RZr0ri5U1XlpciO4/bfA/se4M
CiPnDUtCdqB5y3mswBc784etkBsrJO5CAV5xvQQJk++AnfFdeCg59gHJxwNlSr6Zc4SHMH+tv+3S
p5nDupHN1RxlJGKJNf/AFdU0nzjWzMffOfKfYi/7ndFMJdEkE6/AiFHdzLDPvTEw3251WYLBqN5d
5lgxvqaljf/CV5XVTCNLoJYm1VLFVBVtA3k5zSIJE9RG9MhKigNodR3OjwnRwaxbZ3f9BT+mfTTj
Ja5eX+Rmv5yKppdAWqdT5yaNItuGBcJDtlh+PzDro+L9wjY3Q1Pn1Com4I+ZUsgL1n9QODoEKOLU
8RdpbOoc6L37/nugLP1zhJisWqvqiKaEcsS8wlhlNaMzNL4gonxH/qohobnFe5oI/9mWuWaHoa1C
boDf6xqwRXtOP7G7ZjXSL+4513UvzNX6crfzQ7YJ7kdQZV4dUZ+bZnK4tkjtV527gLI3KsmZ4VuK
JUx3bQvKry9XQCubxIJJuFePSf2jvA5S0R0/rpTC6WNYkEJmJRuDt6kqjQT+YitYd5nhFLRXQARp
8745+TNM5X7XflfczIlhv8rxfxmWOEIO2onieDcTO63eNuX/hR6Du8tPFQqN47hftpkK1cYyt+AW
bqhEnXYCY+8Xnjy1MH1buxsPhPcAhLMJVOp2MNVLpEfjtUEFjYePOpUm4QvEQiVpfRd4LcM2okSc
bvFSobU3M8aG9FzG7A6PiHsjbMRnnonhMb61Tm3mlQkI1IgYoevFT+H2XMyPg2B4qojariqEdecc
lFbWNdLOyEZs9IVksqJh69qpkVYcRlB+xtdskQel+eh8uluwJ9F7PYFk8l0aNJC7GTSY2fBW1WDu
RQQUF9v+8JSA4G9QhSSkQEtQzdwxRf94tF2sEKhlwyMVJnR141CEsme9TzsiZmM+O6SgvTE6GlD5
yBnbAw+3uKnCmJUD7r4ux/ZlBynKJuSr/dyUKL88/4k6iNigtNnNi69r2F567Php7h87ByPV2qff
i5ljSao6VuEeKaKECLIoOA13nonnGk00SwyG08sYyJ+tzXVvzSbPf+NgbBPCOtlf+aYLkMvh2ESm
ZH6+lECzlvHT2awURP2BZtnQ5vfMwlOUqYGm3RQdyD7Z80FrDZhBIwLzz1GaZriBrnm4JxlZk9iu
Sx5Ret8pAfrSNi427w/zTxlMxZvfDOpo97AacqF+zqgekoYGTdqbDw88tztG6o7o1VFk2RdI0GvN
ObKenzMVm87CsJni8HHnT+pH8KnoGSUdup6WCc4jir/SBLqjwa6kKwSOpyeL+O8E9vrik1gSncHB
E5L6CCoqhYUUKh4Oc0IV9bB6YK4g0O/p7N4fKEacJ+3px2KDemHcxAmH/Kc4ESMQX2d6VmemKrqS
IKx3+YfcnqHHQVyzitHYUu0u9jNJw6ovvPYICE/hvAYIb6MpZDhAHhXwYEeYgp03ywIBtbVz3FcY
obTqaNVsB0hkPL9a5AnC23KYYIo9ZQ776AxFquY0j75zA63wD0aOUQmaceY7VkhZBmzY+G2dx/YE
Nw9Oo4Ug0VoBXx8YgY7rRb7+E+P8pbuu6FOTPQjxJ86Av42tympfO0mHeOs9ubY74ao4k9ZxQyNe
zt3f5hUeYD//i9UVVIq6K8xO+oLLDBj0GslMyD1ekm64ydCO2USRvQJTPf0J4FNSSjILLKNiF2dl
X5wP1KvW0VdQH7c9jVvmIz9hgo5yKibwAiuz9klc5kjx6L+SORsblvnAoHtHKtOc3xIw8+LHxxhd
Dxp820XnNGan7uPhwcBmenMfsRF3G3yM59VihZsMJyM2bqUkt+zUgMWauY3gHY7yZafvqRvI75SP
klmmyIzUw1Hc0a9QGzBL0bOfRSu8iLo5J31Vd4tVi7lYIU3SRUQn+TpHfFG2/Wi9O7bRj6M3oXAO
vEHqJt3Yl6C9XMATzBpLK2Hi1zJR/Qim8jd5rcKfbo0qKE7ozCqxDsRITBV1EEmdSyqFSO+V8KtI
W6N3ikKyq4RriBzoYFUPp4ofIEntN8GZjqv0C6m3OldTO8oju1j0GDUJVYYB5Re9ShyyEfvwrz6B
YHWPIEjLQeksHoMmgsWFes/5h8AekptdLKFtHi7HV+v1GNmYKqgjZZTBNCvo7+DqEveU2oiFL0JC
VZvODyh0ICjOz3TXI00ND8226elHZwLqP0TEGiKOC3OCHXyF6LbynSyVXlgzu3VLn1hR5LqI1HES
kYJphLkEL0qxdQjnIjZWEzz/EFgT0OvWaf6OBkXEYg6B0PPvWoFncPbOvsNaKbjVX7r92umZxjpW
2mw1/BgGEbEGkRg4t5JX+ez8BKwbdTFv0vW32pUVa0IQCVu9ym1P3Vq4lY+OZAA0t9DrCWRYYm8t
f2LGShgXamXIG5i+rRHopgKE60kiycqbgRZg/nhe15HZ3scwQrHw3HuhmKEO80mC8dsyAoXF6Zqz
iF3YrdgTqk9tuLec9fGu7L3JNqCj+2rGrmJ5eApWNUvLj9wo3e9gVExeN5yxYwuFa027YoV7a8ge
oEGogEKwxHECzfo7F8zwSaA4IANRZpHiqrB6agKk+z38SdapnlmARveXJKEKzhs/O9y8BZC84erV
k65vZtpQIA5OF+D9Tr0pZ6wIvtHmj+EXXot3IxS9iCVXnMy8LWm1C+PDkgj/ex64pCIPE7ZIhN1B
BucHUJOa1lNcb67c2Ogdq1b+qW/UFDoFFDJ+55OsEOQ+cRHpV9/J4lwM8fitmXSxvmz6JT8ZgkKq
gFxsi1uoGLLVt2zK8y9hbYfVcxE3V6VVt/lfO7c/ZnYCdKYphOGXPlLY5EyVffFsMH25C3RChqPf
vLnw5FohPi11qO8flQfNd/KlfXeZR19iA5/qGora8xBKaO2vH9VL1/BzuWQceTdKpkzicqYzGfrk
bDSBJ6WSD8QSkbHmCZp84UwvfXFCGBSWpf2DP3b1341gXgxTAR7vvoLP2Jfw0tgYYQMagDnCPFk6
Fwlx1DtzngCrod4Y4TC2d5VC4aqiy0RO0SBAvrfz2MAL7aTYSACWFFFTjMhvXo+m51ryWqAKG9wW
PQ+673+0voz01t+t6A0jrcSl6W2R/q2C+9CEe72GKsTLz2QH30YXsgIW95DWocZWjenviY7+vbgv
8n1whnvO7B6Ner8GXWfY/XZidHXX0vqXj3EI1JCfhIEkUM+fZxQApao+3NiIa7szeTL/4M5wPfNO
su8Jyrmt6npTSNCfnR0ZGU0zL2rN/+LaprRsmusME+yCeYo3Sf+0KDRyHUpAYq1p9+e8+miXeyhx
LfQiMj+z/VtHVRbhTDlbdfpkhyfZGYxHyZtCAId5jDHTLG41wAEUK0JL5skrnyWQjY8clILfP4ga
+PcNxZ9zUhiw/ENIBqBr+3HGMD5P9+JIniHljaM4mtcd7uxRLSEzoyHRGaEau6qcTINm9WQ40rdK
YTMk/1lRZaw+3rZsrG98t8zWLQUWCfqri4K9r8EkIjHFtUColBfJt8z5v6s/Vy1psxMwEdrhp3kW
yTTuqAhUTHiRumOHkAjjzYB0glq2LkSbG3Q9/vPIbURID7SLKEwMaAjoL0BAuun7Sl/UVKH52NC/
CwpJoQ9jgSwZDxeceIE+9o/aju0ilh40cpNm9PqZnFxUBSriRmJSeP8fB1KRCQRoDd8RWJ3qNp1k
MGqqmykwyGCW/TzHH5vydHPk43abOlZQTpLohr6Ab6NsSlZme3Y8GNtxI/frebYCtJlTXgUKGbNE
pjzDB5fy8Htv4QQaQ85XtTPJU62Vv7PBRL7YdPNL+mdpaA/aBEG+tTTLuNJ9/73yYd39mMjakOaw
FINtawcI90cqzjZksZDfP6TOWkF7Uk+5JWGXI9sfqo5iv7pOP0qzDNcdEgxVXveEWLQQ3Pva6Q9u
cvNOlpiRJDkKeOwtu0xt97Uh9gBuQzc3p9t6lsxVycEywGZuutlXFPyU/J0XNt36RHs3fXKqprBc
sWyJmigXkQRgWtsfmjX/qqSMqX5d/FltQKdGSWDP3jiZsv60VLJmNERn7ghiY6QSlDVtzvzgbnpk
W+8VaPqiwNwzHLpAAhjHZkI/+FjBupbEVbthd7aFio/yZTFAj1mqjuUXUB9r+hnLlDz1bORphKsm
e87455GT1gevBYHKGhuh3edn5gkCkdvzp4KGFi3RDfLaUHE5wmYn1Tq3VgNLTwXnCneA5oZbcMsr
+9dMTOjkvDWKG0YFZJpfUsakMyybUj6R6BQo4+u4jCW/zu8QN8DSjbZN/pmHJDExxlPC64L33XlC
F0pkgrwhYoRE063pNpRyMRaqkMZ+wYarPbLzpp28hwwFXvHxO+syQ2/k5KZD8/bmB4pdBBNmbLAY
9VYi9d9q28bsISlnTbfRBt9sxHmfcUPRVl45ram72g4Q2/3FaGsXNUN/Y78Fc9VtIxQQfC4nbECa
g69tuLEotralTK4qtPt2GT5PRIF67wxRG7YGDkrZaIKDVSOYOkeK6y2H3Pqj0hRmvtFKwxNwxZqu
7aBan0XpDfRQLDQQUIS2CYZ16Sxg2pDFjkzAuMR2hUYSvKRbihPf/b23QQ0A9op6ebuOqzSS824F
NT7XA6Pn13wDchX3zbhlffeA8HbavjY5kCorXXuRSqlYDrWDw29xuemuy0o8cqzHo2LTzH/UQG89
HmkcwjqasKz+w+lyLG6mOZyJL2tCRc3Cr9X4SHSTxffU2TAIK7KFHUAbIlQU2YGTERR+vAGL4/ZR
gn9EFsd6+THdgsLnYvmP1wZbwJ0ZUshxY7K2iNll3PFHGIg6tctUCNWW5WJcrca/bx2N7lYAFHzk
lmqNXQiCYrUay6suqnd5vWGg6MQL+qSAETdk1BYL1cqb68n672pXM+tQfewOJGTaSUci/D9weQRs
xsJv7m7PxFyTI4K+8U72pohOnDcFo2AyQRrVFbvfiY1GYuNBaXr18HM09kUQUd289sCdd236n7Bc
RU+/KrCbWWC+cZSpi/YmFf1QQolvcKZqcGfki3mPJZhRWqe0eYx7wMg0FTLZ5MOQFpzic69nGJGt
8KdM90MpUs/2/85rHUf8LYnMgZtrsyYAvuBAIIdndaepkaSzQsev6tzF8d7mnFt+dZAOZtrDCm8D
Z6UuuZuzFhk1Xnx8xUx8Szpmk+R0TODVfekRvcR6dpCH5/bmMXSmlw1VDGQh5VTVsdOh4Df0fFl/
2MVG+7L5gMkUd4rKbnA8ACyP0E6k1ddSARrC2YdQc9gM2dy0Ly8neHxedyeEKtlB6mDoCt1k6vfe
5za0Hrtf1uPAe4AMhdZYyIxfrjVIdnSFJcUzI4frya49i6hPtWirvIxNNAw/Yj/4qwc4AOHfdLEO
gcbmo5Ybz0tN6fcL3DFIyOwjf51IxEVxVG5L6tkZ1smcI+vRutRH8QSUAMvoBGsWlELioHDv6Pin
eDYzg/9RbqhfQ7+Z4KFYxNpLfolgGZujHj85kEOX7D5AGAT2ov+Ct5Nsx9AkqxNgTx3KNo3eRWDp
1SFvi1Up5RYV9M40zg2UMLigSJHyC1UYhnSWwXtlKEKhsm0k0u0xwcoPkE+foH49vbREgpvmgeE8
8lUIsa6QXXDdhkN0zQcIqhNQOGBrx/jLNNGPnscyALcTC4W3FoHL7BriL2JcB2T87BiSQt3cJXHo
jzsfYoqUnGt8WyMCCW2R0weMlAJ4QXDSuhIXvy3yws1eXNortrm4cHK7C9sarrAezycTllazzFsg
ZqKbWhUxi7bLEJk2dhYvCmJ4NUI+qm3zhGMGY49GMUP4NWM9XBNG4vUMeSXslgsm7P2ONLGo/Ep6
EXoGxi0cGLeiObh0O3D8xN3PcR6a4qPzmaoC3+nPlE7P8gphkQ7xnICQNcmh6pT79lb1+4UOUXdi
VUrrS8UY9Yvtizdkn5BdEeeI5EZ3WfQLGkFUxmHFRrCAFG885Hxo6ltuus80MqwI+XDoWgmU3rnZ
Br2ZuGRZBiEtD2kOdOIz+YhcfzW7EX8MN9ZG7WQOLcsQHeXi2ljP5LV1RuWg/iIE9K7UWaRueDoo
2xrMc0NZEYsls4fTeW20u8CepTRZlkbt/RGzRT+kqIWB4Muz3GD0/3LHDCMDKVX8QDu9XFw9vIvI
3ISsmlKhpYwW57LQ5As9EeUqFzjh05Gd0B8P3f7iH4j15XUWo53gXiU/APNYYooHC6m/IQI2zDHV
mc+PyTux9fdZkhf3olOdrF2ekrnhDFPB58qrJg9eirXmiZkKVBfpTDMtoeNwmtVNISaImFkRfHuf
h8F4fzACTwwm+amcqHMJGCGeE+G0IP06rRWZUAcrbEL5Cbx2y9xu9NmQW0xd2s4pUrHOCjPmve8t
PuetiIYptF0cz0mrwV2LTYCLsDF4xCriXJZsZPSgv7IoXMGHbnRFMto1D6fzTCsv4NLdSKWPkVzm
Aks6puhxM4xvMizmnQmwypl252lLRTy9Ut+qd1Xx8w5tQ1EGPRCzhqf9KpcDYhE9gAhlhDe89HPV
4yDVoe34TvX++pQxyQs09FEdnmgV1j3MNfuG/2lCxFfDj2c5USDMvgtfl6ybc4mx9oC1XOdyM6Du
ocO/KFeOR6RnppnobQdTk8jUKJUfsGlhwhgyZONYQ7tRd3Q1yNSmEZ+D3m4ewz2HGhdCBwU84H1m
Kfu13bLoofAWKqyTmlrkkmDy7uMd9sgp9S2XaQuS33the+Bkxq9jQaWxofz0Z+wq40UemzLIl/l1
JLZgTpnDxfoOj2KgMS45VXXNdqmfWUje3ut7sSc3NjFa13Bl296zHX3z69VumOCfvaj0CIX5oNBX
1lD7t3Etwb2QLQ2LoR77iCjaXJh6OFimzdGTOEH7Hqgr/kcrN8yZkCzjZUhtEZLNjDRifKSz4sK9
xX9GJGf5lNIPmY1qyuy1JBFVUckRrR0Wq3m5ZDTOcCG6rcUC5m8W/ppzu/tFuirotTx/62g9Vvxm
GsurkVJpSYW1AeNhETDeYWtuZyvNkckzFriYy+9JrOpZRM9zV0rSvwoDoxDgj3FzBpvBHfmv9OLI
YDTeuc8U11452/+UBDZ22/aTk8H5GUCXhkN5bd2MqPopBCA8J8WzvuJkjTepxDiCL2G6esmy/7wc
KcuPr+ZBm51I1ObmZvIB9RVnqOA+ldh3RPBL8kNJNRCEHb0lb5j+XVij6nxA1GJCTdTnOL9/sfSb
O/lo0kNkDAWtyFSSUGB7bzb0t3kTZ/gQAdH12tXU4EWL5mC9am1b6iGK3ygf0fT3LCqwNNaQSYYF
Y/rzjeuY8GfypgHgbsyCij5y4zs5geIPxsgn6voxpHEdk+Z+bS/nVXFGFuV4YqoobUWiFn21FYZ4
ex6HlZ4WWOoKXgUQKSgCgn8bAaKqHympt8V2BTBut315+46fln1U8ttfu/7HiAE62EhtK2KoPY/D
BtHjNiId6L2MkM4QtwZ21IbPub4THEIczANjyHQg6hAPdYFCVaODB2KbRyV16RQ304bsk1MaZJyO
dXaG7eJDjNPfmKdH2Plm43i1+gDXWjNVVCPJTnPGHvcUhuk+mcRWvYPe/BOpdKMrbOVEv+y5nzTg
8GsA7l7PQH7bo49aiIc7Xu5Dkej9lT0jXghlidL/nxAVeLYP1hOA2bnSd4ry3tOzl6JugnwjMqGn
v223XzMStdH+Jdod01Lx9jPQ7BU1l7nT2oxUD7/v/SEFRE3kxg9tAowqqkLlNiiBLIQCGwnR41bJ
3enS+S/ijw4zv7Baxv0w47rr1aouSylX/g/o2A91dImn2ctitaH6anjxQ7ZdcDvKPsdHUkWCMe89
6G+cvaXcmmmtTFcJ9yIi9qHLrEJQDmtK+zi7Zq5gWxROA//83t0j3IfJmoXciIQWusBDi7jS/3hC
TeBb8RtQxDAHKpoOzX0LaWZcsT81S4jWQNqizYCmxDkgCl8lUKs7b9dYnXn4GanbuSaEbSdZZ1UF
ogsyVQPbR8M8T5JF/0j34PrNkkC1/guccoU54IJO9GJz13Ze6L10oiABCRvPw9kPRfnmkiBNUrr7
yr1YwuKZRv8aVgb9ucGiz+uAlk30qjkoHEH0BgXRJb3sWtEJjTybeLRVJbBBw9jFwsSV4jop4IVi
/5cr/EVLw9P18uiBpG8skJ+HaPcRpBg2d2I9wB81YlkO6Wv1veYthITwZk0a/eNbExFMezwVM7zY
DCCxiSlAEbfsOAofFmUdDniDHuxlB9Ehvxxc2/TyufoEhi1Hjg75+57k2ruxWVpkcvytBx+XY+4X
dOibraNp+tQpUBFB1akrfBXHmDVw9Cs53gImiIu0RrriXGvWm7r7ddeByXCnKu0wTmd7CJxQ6ZpM
Qp+c+Ryh/J8dm5NGe4KGGNCGW2WfiGSkZ54j5tTn52vyomBDA3LiJGs3Ilz5hEDlZkT+Qa6i0vcA
zlgdsHiM82IwJ4jW1c67NYGHP0eT5MdoaB2GyzkDBN1qVnCFdpHbrWxrW8wtvhJhBd+31I2J0dzn
TxdWxSCLDWFBa/Z4rdlE55JU0C2QUSjh9hQmGP9VbCwReu3nZHQaYlcjNl3882TbooTb07esfhtB
vRx/ZNcgrgjLQ6DDE20VID2HuK76+uSfLciB7oZwU9ttp4ZaCEHiP+HKpFikHEWwE9/dZI8cTtuU
ar0YHRdqLRuxceIjX9UKt056V3hNGPebBsQIqSy4rYorRAJWgphrXXcUjIZtHN2hxn4ytj1SJaht
nNyldd5u/brPsS+Pf5CciMZnbDjnqsmyGbwHCoEU+IqU/+zyFFZcXf52RN1LNQoZAwcADIU/DwT1
NDis19ophtzWpwg/gN/JXhEIXWzNpWkTCbSjPZun/0snOvDHhsBouF8aiCBlH7QGa+ZYJ4iCXMa0
wrEcZquNDLHDvTCPn7ds5XM4UtnM4USt2tVs2L0pQJ+3lFYF6/tdbFmMyaVYz+Ungx0CBFEsxo/7
qlghcfEv2VaCDMWbaJjX9f4w5qQcliiQuvNiuOgLcm9V7demUFNeWNqFUnAmL9T+Q4UxwfyRCe9o
XZYE9qp3HGpMkK4mKVfOGHJ3158vmUfZ8gqhPblrA5MLzC8okAwlmIvt2Q8Dmtbxoab1p/doEbcc
ESVRFxRcGy8YnrXXdOYAleIMcZ2bizRvx9Dy6ueWkyf9o0uziYjUBVDEWVoTbpLHPeusUBDgBFBm
JMuuQzBaJdvR01r7EZhM1Ddz4ReV4TCM552825iNXwQF1QV8J4QtRlIQLiZ8XxYY6r/DFTpHwcG4
T45psyv0k7ZBDEZ+jb9gBbzdV1ju2xxSFrKVUiw5tvJOJCAmZDiYPTp7j6MlUsrur5a9fsYuIy5I
VM7zEtwtOTuDg0yQrsl9AF3qLgDUao8YXd0s/Mhm42CkWykBirKblw1BpTJqnYy76xu3G90s1SYT
HQedqUZHxO/tPGkydolPp0M5ZUIQswoWyRwtApgxZH4X1mia9DS9wMydoeydjEyVakGmBmOjxxww
txZkaVYs15j+GOXNc21M80FMK7ISpmkjLVBaBofA+RNs1+IjGzhILqd+pW5gG3hovorH4XFytO+L
5UN9C6N9zNK6iG0mUsnV6bsPwBnzYOjTj0T0W9qaIfqRQPtC1TwpgOGuA/zv/xWhK8RZyeHAalyz
QC0vkQiAef7HAiNoiiBCWVtc7hny0wgRp+7iVdbIhAnap1wphw07KQd9NCJMOL4ELSpuf/JANuNO
QAGKB5q3o64mqUkxuDH0eTYXKxFDZ++DzLCYgt9WN+XQxWQF+jrUAKjZwbFvu5n4yUxpbADoSt0k
JsPZy92ynzQLPb6m84zyFmtZy+ORPTAf1hewJ2AMuS6brdGCabrJZRpllFxA2bx4QYcyPfoKlrGu
kcf3t9OJVZIFDGtUSEBlNoqCR78vx6zH9QebvxU6/7aytGh2iwwmco8RyM9Sr1DAkZNPiUJ6bE6G
AAFf5Ql9bGug4MZ5Yf2yNmVSrwDQP0PZrKgbDUUDitKKn+sdD9m21hcgUMasfc55FO9r0SafmqPb
cuWBeQFydIOvzUQSpKc3RW/mY5JH76TfcEvLIQDZ5jE7PJnn53JwjiX53Z96RILSkfSf3+T/9HCf
eBExDbo6on/bHwYc/YY7SVSbD71mSEBgSHSNMexrYth51EmAyDHoMU+yQa6beRgJnWsgx9Wy6YSA
C3l8Meh+SFls6cvTbprdxnC+DOpcb7L5Qo8m2ZZSuUmriFGU0/DbuD6o2akm4MmI5RvaciT2+1tl
cRsyh3l6kfXqIU86ho6I+pyYbutDWrGwjEJinnN2nNnEcLov13I1k90+YU53SuGmr9A1LVOv8875
P5oBPRYtJSb7q1bJ2i3iPa78melpusSTyTsLZKct9gljcGy4oh1X6CLYxhy5h24Hsn5HD3TCj08X
Lrra8wnBILes1yhWmhNfQb9ZkShUM7RCmM0XF/oLENL6swPjS8U3DdlgAE1/cqRFEF5rslP/nSjS
JDpTAi/Ozm9w0fvfFJAN+vFWKx1tttmP0unOemZMCRFAfD1z2b3weQboEwr+Jwf035t6+0T4wUqs
A6Pvdu4JTKeJ1UbersCMweuXpL0RDgcx0RejA3Gpw17GGVQuV5iFVfSGqjT1UAbxxAlF+es4uCt2
cndD/ziuBJNjAbYZ0I+t6hYYqUOjA70uCt9c5dCdiykGlRlB300mec9twxQgCFU7zuwN5v9zc68K
GMRu7VN7+HA3Tbnqmq+tio1eUCi/g4krsT+VQ/HIllwKJNb/vMmWPgfRnLQP2IG8BLHHgALLVWxG
6Z6O+a20BbbXZjPONpiZe1/kpEBkohMBhEY9WJj/kQfUJO8ciE/lsU5mw0QF2od9a/p5DTbM9eCJ
f2VH3IgaxN5gMyRGbkS3/oI9W5Z7DEQCGky6V2oRYbgvtgkcVnxqD6+xQamfw8LOSKe63y69koJs
OGa8Q0g7MuXwtjissqenHHmeBT6ZzxwLMEftXdq0L4pst669+rpyBKCMeqOkHo7/aH9bQveNYCbX
qyI1+P0qSmeUbfXTVRLWqJZRXrvlNpmw+puESjXJMpjf2D9tUGTiYRZdFlgIJp3hotLFv9230FY6
Zae9srh0s4+rvXuEIJVcsrNOI/8Lys6BmfSDQU24c7z6LZMPVYRYZ3cLHagOCkwwKWDmgYWsXZgU
jgNAcISATUvi/wVm4lWH5/2n3moV03o4XQQJMk+GzKe9EChO7LXtAi2h0fO/2CZBhf7l5ub5XkQx
hNkyk8f1lCT44jGryE5ZJaySAFFMF/TOtp6GMaM4LbP7MEnekcid0SGDQ0CY64886XCYYAEumqn9
GVXFo2hTgClWCAy8CNCjENwgMI/2smVRbAP2IBIlJvy1cTDNCpfjnhkWzZ4UK4Ur2U9gciwPawJr
nlJYPtd3eJf2KbfNSHPJ6kAEe8u2no5rmoNK+4x0AhdpjgHOub2OphPZethaNj09c72pLzpD0rHo
+HNNPDdPaGmLia52jvAGBa58fbFIyv+/XbjHvBccRyN+IDzKUtSHLT/MjhLry8CgImBt6O7gBK7F
dqy2p1/OigycroJ6L4P99r0YC3DxQR6eSBbsLTLwt3d5ka6UN/gaTb/TZ40UK27CdTLLmXCKeRDB
UfnlV4yYy1vJED+vW5KBrvVdl89b5PQTgwcVNOVNMFM50IvRBzDnbrcdEJI/jJ+6lVBvZBVfQt1I
M4n6wmLW1rj4CnB4rQK5BKyq1K3HkVrTh2yChOdUbs26BPI9j9WalvgPRxo1asGmI22X0jOELFfa
D0FGG3vgbShYl4pV2W4kJuH+FXn4Ac+LCQVV+R6ixcZEmMlz6hjVnuv8KKdI9rCoQBdaukMnsPHY
JR826Lw1a9ubpfWfnsouFb3c8Qc9eaA/0wSl9wQZr+fi3dRXxOsGbs/mrB2ROLHgDfZcYtw9hPKn
yu6T8Mh87el1ZkMA0pP0RJQcP77FnqzuVk6+0t9eRkDf44yRBJPwBmkkARB3XT8GXHRPYKWy+CYX
WUvPMyNOySIjJqg4s/NhzsegmtrPHvo/ShSS9QjvuYzppsIZNTGJZAg9zZBsKyQu/YIPr52a2V+A
vZJD1diAhfXYMlqepJKvigzOF66kIGukXrw4+sPVLtK8oQRHp2ltYd3/c2Rjj01r9VbkfW7C7l5B
RkC+IrfMEUjTNIZazwgBBylMRIcflQntC1UYA2G986auMIYnMwJOJ7dvkw124ddLhTQ5PdVXX2dS
wetw0u92aRf2sICAiPviMVOC5t+6RxF2sV0dC8sLOnYdEFNw2YekCPoxn7c5m1LCPB8DXwwXUmb8
NIYd9+IvdSVDGOVE4yAvKXlsPEllGxyfp9+/xTBnwSKldKKrmEJSZjnhWegqHIwN8THh40nWJ8ZF
5YfH43haUXWD/soRb4IqgvUbxcNjgunmeH1u4f51cSRjq/JZHmZIkJipu9PY+peRDCwQrKw/5cKs
ZGr+G9kugbYd60rtaE1pWe7MqkTUcPiIKZY/bQIje7BzyjfG0ikLTLBP9ivj+Rezwqr/d/HauRxw
QU2ZUI9SYVsxvsOEqYckxT94+y+9XdIA0LYVOplMFmx3VO3EHkXzJ1wHQ3/L6hTlGrTtA5AM4VVm
GkpwX/DYS2YL9tSLaeHWFh6txucm/AD/BbP0sAEN9Xu8erwcHEQrb95JJgU8jsdc5sKoHw8KkjsP
NVVwmACiRC9PhjnHVWNjnjWRzBzxwEZxyI03i25a2Ae6AWUZ6td9VcgV+rEcNuDcUXFjSESdmnKN
3pawr0WvqePSEekdBGlE+5o7YWWrMGsY26BO76Kn06DLDKFsH/BGXzv/kXvJGix0MFIz6gk0ibTj
nLNTpeGayJ4IIYGFDl4QYaFtsT5K3ZPOxvopF377lUvk6T3ErmcvAFWqf30HWeebiEh+4kXV3qNI
DGkAzjAq5oBROr9sEITKFeIXYx0IhJLHOUAStkaMefInyC1vpo+AatoEV9TdDFPk8b8YvuqF/4zm
sq3lHDPp9BCBbVRwybE6NbQx/USKOz4lbHVgkM9YIp9Kmio9rMA79iL6ui7mfmD7YqvJzZ6qZKuD
imikg2bIImgXjqNryYS5JZOTzthTTfrlF1773AWJsPC225Egs8f+3V0raHLmliBzcF2A4XZlb4wU
xteUDxjugp0TikMPY7oVXSIh6+JQDKVRYoVLINgZ9mKrK0dfCOk720ArOP/cHc9kqVPGVMH1P/bv
Z9GjBwnNfniinvhWoDfTsSAZQiTNFT35ep9Rjz3JlSrOP//NiM7ehvOXcHYDP22e2TsbASLOM8pl
JZppQx7Z74LKNXTdCNrO1r7Xqv1a1gYQxomREmCdcX+tAS0zTQs+qiOWzC6McoPzcLiK7dmxjYB2
rtM9g/VCnN43g9u9KTYiZJbs0ygqqWWyLB3Jk/4pld1Xp0FR7fq70Anwwewr4rGuROysAL3AEJsh
7zSgfys6uf3IxoXD2vtX2dns2vCKuGj8B+5OArZGKvLun7HK8n4nvdKaYkhBm/KFLyyRpi0snL87
qCnTQThgPS52cMzPrRyHe4uu1z9UvaKB4TFFBKT2LebsPCnkAXH793MwTkFKQ6fv50hDlEVRAvUu
OV6/hx+hf197W/wcSQKpSuYejGpJcuQb/+WYTi01sn9o5cIAfvnDuJvl4ZVAH6k4X4LwBPRz2fWS
ZBBMnxwCw8wfPh1eglQg2+I86jOaAas+9ox5v+TwZX0jVB7p07H37HQN1D+YLffUo79qhxcxuTbj
MXVjNXhSyIwDJp08omryUy0nap6+11urfNy5GAOFQGhseHYTTH8R7qjY9GeFNqTEUsxg62InVYYS
ufb78rPsUYoyv73mIza8RxBXkS2UonXGKkoGvHKFCmQ6M8E4fgKFLHVdPvhcW3RlrFnYZql0T3ws
exO4MwtuZ17eUtI1G0u18KZS0uaCLWCuRGtDQpYyrl29SjAPua+4PzHnpAJjVlvL5ahx82+Ij8hp
zmKYx3eKU8g6I4aL7xDYwUh3pfHem1AWORlgcUq8CAbfY2+slTQ9sSEbXD00JmIpzAYV0KVHJRsP
P14ak3X/11+C9Q/YxUBtI5OFfo2l7ifFC236pDt77hLV/qP8xBy8NiPahX72/nmSZ9zSaThjs+GN
bAM+XJ+Zh043lFNpjVon6Z4YDCo5mtcey6EEn5oXYZGqV8rWkhOWjo17Pt7W2YZ8befAQt3DVbbm
kicGkcirzbEF3vaCsGjxCQCAyenK0fO7uQ/Mbt/1p8z93QLi3lHOQLjzF7AcUqV3mvCJFo8vXg4w
RuI6YwLEypYE8j0x6ElxGNFjfC5Xj1CIjLtQ0+I2ixs2VIyFEYjhWcsT7wNZ9/O0SYwRg0iJSCRd
XJfmEWBKv7Iwe1pE9FeFckMkckrszD1wpLGarXT21zdyq/dtp8nLDUY77pgkYvLDRHc5bgKZ1UsJ
qaMNDou1Lf3I3uFYlSMAjhUBqTwKw1kqTgwlIGlWWE7gYu1Ru0StdBxX9idQ/vl48oS5hQ7Ws4Wu
KPZqEox9RE1ng+AP9nITW8cz4jlUvdihkVw+lWQq0/XSsJeyLXf+zXbqzwD8/zcTYDV6yLx48X4J
uiIkIr/H9H2b2fMwcRM07FhDQxSGhaTl3e3E5MOLndoVvlmIuCAZq2fDUbyCb1J/ExjoavNqVIYh
+II0011ghh4Y4IeWhkVD2/hzrzC5ZbX5oxaY8qLobjsVUDEEi+JzlQZZZTUADm4XbkopB+1Q2Xyf
zkvPRlLuDrSuMoTIoZ5Iyr05HGJw7Qyyfqnx8b8er3CWZkKNouOQqbwib9uUZlOO8hipJBvy3jWW
L6J2S1y+aQLagANzklhyLztiFKk3/q1LNba8WHbzFI77Jn/zUhDDf7PP1qMfnqyFh/ajl8ZLXOna
WHhsHSFEMAIVhnoz+cI+8nOkVsObPAYZfACH7A269lJn7DY+1w+ZGCfsGzwHCyKO0qyudvHtn3RW
ta0e3gQAGELYqq2R9cicC336HwTyyk4PZtYX+ZPptqP6OF6lV4r3uuN9Y5Q2YBThxIX4fIjTeftS
d36e3I7oZOVn5iCRgkLiVpNCn3DWCma1V22HJMcrHOkHoOXivfTeusxSCN0FZqUFFuwzGEFPhMOF
/zoeRufy0Tnzd/9gWtKbmPqqRW2bLDzP7bdJoHJUtnXxHrvFQSz+ZW3zNo+7EM+lJrg2Hf7AMK3S
3qGxFyF9S0C1sRQhzK8pdRGe1dQTc+gYJcnBjYu3bQRvEmMuZKwZZ3sIdSy+47vrcEXzhv0VrdkI
k5880RAwnKNTgYrcg/4PAE1UtfHQu/Ye9t7Ikbi/+sMRGkRt8QFQpa22+pzT1IVPeSmOgf4xxQzq
1XFqB1bdmG/2KBXfvnPWzUI4UkJ7jrfeBUJVhdoAZihhMCMAsWjQ9qKjTvjlZ4AlYUj1pHoodp0S
pd27EO6ATj8FcT1wkZovCUXWCN+ukbHfjAWX4onsDnUAyOiyZoGB1m41oR85ZeqLy72WFOCExep9
4XMMqgfn/EUsA3BDn0Wq+0IMze39FTaPtUmU6obhYzSq2S8lgW/KLIDIbGT3urpnyziwbKLOw0eg
nWOP6ex2rrPFAjqeOXIPjIKbyzhIGPrg0FTPkottR5aQ2zZLsqGVZWcJ/ZakHRyxAz/dHySF2oG+
HUs+LWLGED1dqofBpTTsrMwlQmWVGqOqdgE++x+Ugq+iykcJa0xG4Du2gLzwqoT6UdPj1/Wo3nCz
hGQTg7iiOwpWzHsBPEYxKUr+cSqS4U3xvcNB2Y9kJewGsmGYuete9Sc3+FN6qj5A2zmMEmvyOr4x
TtCU+FyjQ6Bg8kZJQ/MOqn0aVOXuL50el+Wtklxvqv+FO6x+6H2tvBbS2N4Yxejyh7cDt4QUjDMl
4zm3Wv5tMH1CLrIvf0oc7oqN9yoBUJs28pUnsLC63JnLHygMr86Kf3ApdGt9yHZfrjJ39BrbtV9s
TPGirCGCLIuILNle/TyI876aIDricnfH2ZfGwCvbalKDOt1VPsCph1qIkrpIrHicHPugJXUl0ddD
6dZdYxdlTpen82P/i6kSmLsh+GWeLqyHib8onMv9jbdW3i1bHA4NCthDSFowBOKqoapE3ANGxGVp
rTCjbmAAwyN5vxzuWuKl8uDXVm7zSfDAwbI/1mz6RkxsLy0WZfs4TZLqzURgssDbxcLtw5LIhUpY
ToA/GySeNo8RztEwT8PGpbrTFV55iLNX0sivXO2z0PaMipeAFV/Y3IvX1Y2hbi6E2cmVMuaO6b2+
s2ldLRDKyNGwiifBv1/t+sZGoT+Yvk31QWa/gr68qckN4Gp8s6OC2KLlUpeaVvc3+tRUmXr2MleU
uvtWhLggE+oekh8454Cy5o8AuCR5omfohHLgNteNIlq7liD3pwHLI3yt8sZ7jHWKMC8t7BgCg8RA
RltyfYnWuqkpPhwp5ADC+h3iW+tLg36UdaherrKIzuUuY2tEpaD69PZ6tkEOOq0m7xVZY+mRd8Pf
p5Vvjw+FrfSSpgN/z0GUoM+F900dZXBB75Xs9jAqAJPoRY13vhfH7EJQptGH6T159PqmBT56y2bE
2GVF47rRQefflWsSrjBGSNXs8I1QHiGldLJBak4kYEvmWPc/Gjfsy81IpySKeJM2b7hSBrNDotKH
e85TmeJZusnCqnNQgvESa6nNDWP3ypAyHJzvNaMClpk2xb8p/g5MhIzqA8Q+kbbZZEHQ5syYFZA3
veH5e/rGNyjA4Q6r2rYG0IGDNRfmm/3u7bWTQ2Efrlxuz3aiO6XaBe28LIJ8XD7w7+yEQN/JAQEk
4JDg8uKQ/0wMaifl47fZlK9EKF6/3AA6fNhSv54Eaj3+YUH2IJWiBgrH6a4TpOhNaGcgSJfVM5If
sX0bf/i85F6qoTEvEFsyzIXZXCKYrkbkAFxMIOUInTjx95W0RpbTgr5an6PAPGpfQgOtqP2qRI0D
Ipka+jqkLXCvJLjOVOF7nLI31x3rMC7ZUVFsDqsbQbuuSo6VI7qHtax7GSoQ64ltVDwGNzM5ASTQ
nXwGpW2T/U1GOCS9YmuTX/JN55Hh6pH9UxzaLmOg463Gznop6m4+wPPeVIJcAk4OSaSqWOHBjqyW
pNrZbCJjsjQ5QvKzYhA40f52g8BtaSmHHvAa0Q8KU/AX/Po9JxImHC+uCzFHBRTO0xsegf464Cdq
Z2Igy7efKyPLTfEaOreI249pgQqQ/S/UmxxKgqXmjqCRLWPcbZijHlNDeT5mMB9tIPA/XTMNjDq/
ZDbnf7MTwmlEv7gfY7pcfMu3OQ3RZ5mWjsaOFl+y/bBNrg+hU/GqjVttUxPoFChDwxHg5zG/HBhz
/LnL+agp7DNVNx96Eej4mHxHL2H6MRa4w+zVU2keLa20xMWeBP+y9vykcGW2xTiu50g87JEa6Z4F
iEGDQxuESbT+oZfLD4dKjSeHFdAQXA7Qzsmps2ReDvg/iXIdL4B867/GluNuWofZRzQGUQC/UdHk
+Fo63mYfGDZ/+1y8f+qAFW7s+XRGeA+qsrUZEbt+ZfNwcXLJsxCWL1tcGntQ9YmkZFfvvJQppy4T
Zpdc87OJTM3+laZ+Qm5FaZ876N0IAsc7k6viF667WkYCWsIW16QsXK4vLPQDqd6YoALmSAP8BCYs
SdrqEXzE4B3Td1wlKH3hAYAeblY7Q2Z6SxcjsqQuZXPeBrD2TrP/P4VIOhmvhRs76Il+so+QxR6p
LOjCBmeTnCc06ai801p5P9pwMOKM4WW/NCgmC1jK4ylAsIW7izvJU43lV0aIXdjaO+Uot8WvSNYV
cl4fMkkvvb+PmjXJAMPNQ32oGMF+YaWRc0evnuguKFeMvT0DXMADTiphGkj5wuYbny8kPrmSheBX
LloDGNnvfXOsz3CfOKLfIlMn5RQNovdq3y/g2n6aN53t2Ydwv1dBoPpqvqsHeygKEs+WxU8FbknN
d2y56rS4jrU3ZeYX3SAcaMZkuo4KG9/Ahjs/jc1mO0yo54eJ/mPzhNpVP60SX8zVQMjyqODPfu+X
yYqF8jsd1gMm4zqa6WAMFM8KhuiCdBmaYt4VrzjFIDKAESYY9iieZYPC375OhR/xSBl74LaeID5+
Tx0+FhRc6q8k9qZCBUyt73RG8kf4xnqfYLFmjhh/asy8nu/LiQuXixQfYoAGkZYVAkVG9X4vo+kB
tIaIKFfS7GVoWoE0GBTNB53xNHIXZNa8Kw+LKJjUp2qvQCjajWZrlNZ+49J1r790QB7dNQ8Fmx6l
Lx9hlAz24amL38//inwAgMzz9pABqcGTp+wYhNS49khYgkjWzdquPem/VGV4og2AM8nkbH7XK+P0
y1ARWsEbxq/+BhBEtymvBTERmPcSBC/Qh9nu3BJzCNmQZs270dmhHsqXKy4X0iCTSt5n8oYwTlvs
BwqeHMeEMRx329MmNAt9bJzoAQDaWEmVdKHRNwFcGIosq2k7oHeZoxIwp94ChtL56NWef2mKQqJu
gMwog54UOq20QBW4VeDGEJN6nuVhsYXTAblnWTZozmwjb6j31+h9NibeH06e2lC73epo0zQkyXdC
cqC//sPsFsfcDy91KIv88zzThSUKsn5B5UqmhsnlyUju7aPAWmZG4cObR1zH+4w9vBhwKqnqJWYL
3in6FQflwupXOVmjyPqR6Frhw88AaLdVyMLjM24OcC3I3LWfb+CpW6rHXvTNw/hn6DlGz6DhY7gk
ga4vnQZ25musX/+dXoijEdMB93MeDYdYo3CoHka91DLFENV/NtiUG53+uihxlw25FnPvXHy4v4Nb
7FX3s0pB+Gv5rY8jhJMGFaXTDraKs539zcoHmZO0BcRDBglfJ8PstrmehQkAAUWuio/hSR6/UHPh
3Ir+3rv+svrFZIKxMa8jNMY7KRctiDnxWGzbqviTll2Smr1G5ZAeHvJKVfNA8E17y6hRo+cUY9g8
iQA7PSSTw8GyE2DIUceVCFJammoyLxAsW+q7tIxVLDxOX2KWrLr7K4azHD8d5oFSBPj4Ny25Yr5Q
CZjQzxDswW3/CYBsi2YOH8RcRX2rixdPcDL2KNIjOJBCqYnWIlNgEALLbXam4AR/SFQdNzEd4+St
D6+W6mdsbpWct9slROYQssdmEcYhyBHUDk5LflVb2ddsQtEu3rDVwV/T8mXCmSvgmqjMAccuWmrw
0a1/dgvPQHYFd5QIdikn1WYGAH5iymEs9BCw66PMB8kI9XMeA9yRTdOlESZfgdRxcvoptLNnf+PN
XuXWVCRNR8Ug4RdgUy8lHRGhrQXl7CXdZ+vXoORti4Gk8bfUgxWIKwVI2rdSUQFG3fU3MXqBWEU4
aGDF4R4F7HnHbwWtd2HCQ7X0rnSXWwBIL5VFjtl0IckgaRtFMRgnar6F1+F+LguEbyKerSakPDn4
0m0KGRnM1HT6hRubA8Q1AiP4YRc8NQkIu3ZTRhhV9W7K3OMGca4yYjhKVvFRi69S2rhrHlA+LXYb
lebMRUMsB3S/2PgS9IVTokfU7EUrwG69NrACPDtspRHcGcaV0UMb7AOvgnbBLSHd24CCeTc5xwrd
CNV8k0AUAJ/b7H0TQJIDdh5wOkhXxcZQWzGKP8zUVH0zbCw3KU9YIH5JsY/lLKQiOiIm2ClD+2tg
Bi6wVdfDxJjRib9ooC8sqdpm7mTHw1jux80bBDUlfq2ugMornv5GTmSycUgslPGOPL9AAvhcchQP
/xjgeTl46Si3qAeSZTmIN3p7yfqVYllDr3mdsc6fWWJ6Xy/5Nj+jw9PR5B4PiWaJHYRoxWOuBgyx
cLAkDbrt7a1d57Xj+un5Zt27hwJezFyWbV4b5jbBiLQLtQH+3tD32ZyUmXi8BqL0Is91hFH5yMWd
zzmYuI/55vLUkWImwWcZTnHwnFx9dCt53h572P5RlRqzs6qCldMxNqbJ2yifR2aTxxIMzUPYCo/9
GoztFVkU0IBP5rwJgNjin6hqXF6A73GP19CjjPoius9alRFAIrgaUGy8qbqrolr0gT4/tyUAGxLZ
gJHxl+btOLitGA67NCZqVmaIM8y5DnbuV/iBn8YNJm3KYdSATWAS+JGUyfIVtGVq8wO35RbZ2OMB
9wtYd3I9bQylKZjXt8h2SVFcJ/LcCggYy86pt5YFEex8eVU/hXTyQOf96SFdyam0aPQtEi1IrXuM
vUqZjLg1Nv5j0T9dGc9qALfbieEG+4ET5LOIzbyI68Auvsw7jstJGL81Pz7AA0Z6SqnuDDNNFPaG
g8J0p73KmqZgReKAo+HdcUs+deTkMIDN8CxQzCdMHsrT//v2yot/rSbA4GLSspNDG69apATHkjl1
nqM3kHpELJYhFKeYq+2dhhAXwGV5ziuYRScy36Ko6eLBoFUzV2lY4Lft9e8r5s1VajOgiiGlMMdZ
QOxA9NdiT8csXmYasgTTyqzUCbuXqtjghq0O8Dj93QgpnsM/uPj9qmrE31GTDpWwIhrIU8Ex+cH0
QoIGDr1qQj/bDgGjNFal3FunpwjytqmMxNXBRnFxggWtwGY7Tb/Mx44dwin49cwkJjgK/ufbYH9n
9iaDLk5S8yuuS8hvTGzYhp1guP2p+zpZwGG7ORS4+h/qPcvU38zJR6zQtJGkxSMUPVmq9TMLcII5
RdSyOWaHzX9Uxm+CCZIifmnx4PwCNgW4Z5+c14VTGmpURkHKcuoBXjBarp9O3U8UTwoRUsnG8dQQ
h/Fnx4rfn+xzX7/qHuT0wGoKMbJv0dm+mvybiOz0bW/rh86Lw/y9z26qw5UiKgfkQzp/cXLFN7OK
MlJ0WYXr/PDDHw1dfpt8LKgO7BP5C3LhElJ4vmI/XlAprgHxMLO2mRV3IUtkUHhQ1zKIWX9dXu4I
4LafdOLXG68W0YfxcjXS4EM+LN4kCmQRv6Ha/QnocFIM0aWFdbvMmJPIqZwKtaQuINXzR1swrHdp
MkGKgR8TaOE+YNOkAZy3I3NvVYUTUQqgIppUqgWm3eBCKBLU0TaszRMNJEylZqspKH8YHFlPtejz
BUEdZBNLNXwpyjHNaylkgLnaFVRsmw3dd8YvSN1f057axE2F+fDaa0M/W4KIQEzvBrJPDf8EPj8E
zaXqRbmakj4wNXhx/KYt/umm+OU+MehzYTNs+a5a0kcW7dZKNdI8DlE5fVaYvx84+slovQ/d1grK
77PKnNUhiRx9nZ0olh4tVic7w/icvyWH0lZiTXkX27J21Dk/MfemzsjtpgsJ9fa/v+UcKCnEYbF8
XYqbLZsxqHYM66wnnuevZ/KLe+rqJrvjr4mYg/+tMmeqgafNftY/BRBBUVQ9eLoT1oJoETc8OkhN
qRxq1/YDugrOMbmy32Sc45y9cm/QTBh08DFOVB+XguBnXiIanDciQu5jUMtpdSsjJUwL2IH7xyH/
0EBbcC1zkMA7jnKJMbLuevaXjvEiu9+oztc+72MGoGT8z6s9kBJGmobUMUMhQLWLURBlSrQD3OyC
nlMCuud0As6AfPztePuAY8O4qKT5zbC1+Kqhv7hQzA8PmRJjz7CciDAipcdLt5/fs90FHIGD2RKM
c5xsmzSjJmO85dqiDdKjbyB/X/ebaX8rzDO+bnvwxdU+A+T4+W0ZCDR+ZMLPouF5piW2qzs1FwPC
XWe4arpZ4rtvFhiSRVJOA0tyFBm5f77n7JYGXBy0MM8wvHn0Mo3Q0onV7BuxEu66iwR1QX3dsNgf
bXhUbpsbG3TXLXacFifZ6BeacQyTxDu0lf3JKw96Yue3DdY/9gTGh/QulGVk0wzxmwv0pLDthP4R
cPCqIyk1gmPGAW+vz53269q0Q2bMiqhGDlZiJo9wsIe63o+3Gz8dOw6/fSHVM3ZwFnQnNdA4OKND
DpS2C8dzMh/mAf5BwwNBrAX/mJR8yhcotCGPE+7kNoowly+/KLkPU+IXgWe9BkrGF20C2Qsxglil
aGhHNQLry5PvaH+1KRie4JbZ75dgaIrDRkmvOx+/AJ4GF8VYxMiRb4AQ7hOM1u2dZCJ74obn9zRN
neWhR4WqyElELA5p0h0B9e3WpBFhQ44FbO52kBxI523tp0sT5Ef9nM1BtDCjdsRlZC7gTXjxJRWP
KudvElAvusEhviQR3Kdc29Ip90fvbJEMVqUNVkv+JF3K3VU/atV0fBTaZDrdbOvPwE8tpKuGZB0z
h7cbV9WeDypGDO+YjLM6sTXEsZthFsSFku0rIBjU/hvOq6QyMQ9FXL9u8kMXc1iupbGigYWRHHdV
U9KRa2GhSZ/jolu+EUnS2DqQrK7iI0O/59xjnMMoOdjpk+Vv2NGs4/9zkLp56bMBmt0762vituxf
gntLYIpQo/AuKbDxAhSzTScC0Q53vCZtgV2eIVYE9/xJeIO92vBWBueYMsK4R+tVMhNOyBlUKSh3
Xoti35iF4VJ/OMQDwn0tCsr745gNfA0SROFiP4qayWAm4FxVQWUchsD08k/gfRxlpF8z7bndxhjN
nidiG800BiQD/lthZtHcIQnVBe3ME0xbyAdixJpKTTukPvkHqQ75vddOWN9QebAm1GnLClsiKhMs
4eo6QjyM4SkAg4kNBW+8Ue/+SCJzLw8ocvA5se6MMVawla6WNl8/Un6Q9NHpu2UVVxGfG+7nfMc3
mqwPEj3LOiSGyRxK8vPohudGnYPV84dBMVw91wEYJ9WhSTKXUMyVgbve3tTo+ZN1RhpA2FNIMsJk
ChpsZxm6YmGmpoiOCbHj3IBRX34jMLL0DMh9a7hFaWYkS1XhC0uc6UF0th/6vEna7pH9/3PLgwJr
zxpYHDAY0ixwvBmKkr5hU3b6yaA0LpOzsGFcRslBb/j63G2SI5Zu5nHrpdzJ4mkfRKFl5xUGvUps
QHaxow8Pk1yAFah3mZCuJcGnbSsN3nPvxssEkq7YlHq+GImPluqP3as2qwGen08ZJPNsqELGWk3j
vBTS6V/7XIHERc0xgD7shOZ891uC9tb43YVkZwkK88Am1LKmV3oZRGfMUYtksjXgskbFMTVOyzsq
0f/rtbv35d7chtCuAsWGF7YNmhICBe628xAiggZYlzPIqDrd2WhUjc//hZXByuxhLLVsQJmj6hFi
k5HS6aZ6Rxj35rvH+Mtogrr8ZF7SUY2G1gV5cl2efoE1eKITlLNBi1eI9doB+s+EB59rpznus4h0
S4yO94tkWWy0JnXifj4j1bmyE19D1zvYuneinnNrYUQ3sefEVfCWrWUiEtYDQz306UjIJ7VNJ98e
vUpNbFfyQl5sfLtxIRNlMJXZyeO5fwsDs9uj3I7GZf9vd/mjnZ5bHHkTJHhtAMpDAm3LYWetvQip
O2KBSPerejnE9gZ49appXlq17ZSvXu9fb66CYjOb9djbkfxnm1yVam4sEhl8IaUkCU10F3FGeUTU
U0VtXmFXt46d58YwkrdhrLqZMibGs6AqlhFEwijSPPsdwb93vsO4FEIeyI7HdwDzsyrb2N65igPs
Y2S0lGVrl7oeAvCYH8X1FE1UUx7YhUMqDB6akwZ+sQ0Mb0ZsdpnaQ59+ppJ+SPfZhun28SwegPPg
Ppfi8qZifUiEE0OR+s4t0oqWxnJ/6yElKSH1U7y/ot3Bt5sNwhq+Tql5bw1crLvuD3d4Xks5l6tz
ZHBpnn1/Seu1cXwNg0k+ySbnvTtcpt95W91ttSb1aBP47CMUyO/md/52FBegZgHUTl2tA587kPaS
Kz56o9e0dSo7BQFp0gpQ7pATo0AI+RL1PtAddyNrP6PV1gzrDJtKNdPPenFgW4J/NFPVyuribRVT
6kbI6tw8DBPSoTWaS3IMiHJTTNcuNtCGg+pDt6CuOq7Z9M3UbVUZvsN9lyYBLk3EpUHpVhc4gOd0
6OxwjamNSBX/UiVifHj5z2LceQCU0Ci7igFaJXUAu42HBN+rW0OnYI5XnlhdvMkalKpbjqtv88hF
X0cHAVGwuh08iLm32+9TofVRToG+z/c/5QRDRwd+pKuAv3C7YYuNV22EDzzbh0H7uzjb1CkkhVoc
GoB4CoXOs+c8vppy5MbiJDgfJRi1JpL1FgLl/mS91UtIFFxJIwauIjX2Sy08/256oqX07bm+JzHA
C4SPSSsIrxWNG2Mu24Y2HtiJvSplEPbJjtLJ0sEP3oiX26ca1IDAv0gdTjBQ7N0ZQIWiyJxjOlmC
pHVJOcAQPNDJ/Z6rA7JXnU0EV5ZbY826j/HDUTRoy/YItxYYf8g5Da8d9PN128kzUrjC3bFCQVmE
XzsxUKgZG4X45wCNqeJZ+K+1G7GEK8WruRI6wXptPrNRKfc0YKmieZxyxFvhGMpXwgAUwZ3OxZdF
dyGTw693j5X/Dngse4136t4qqrrHykaeYGA5qTbtlPxxOgRcSso6zA3PHsTJ0K3L+nk8ePUCsFaQ
RYrZOym8FOmVUn5fZ+L8pOr8TTCXp85xRl8HMfiu4edfEKTSUOGqXfFFIfT4pd58BS68UXCXIc23
uxdCeZpQL+aRMKCMkUZgibVrftAUdx4SszO8k1bcUgK8FR/OEhDOqXQzjqZf6btP3LxpBluisEXc
GAoCkgpw5mErKb/KPdkIYfi0wM9cIkZwmYVAH07ylyZj1VZLJBj4qskwCBA0KBZ2oF0K6wVaxV1V
KVQFkKdLrvSJxFLYQ8jGY8QPNPBKc188VtyccwVRdQ6HId1qNNd2pO9F8/++RjPfQJVCnnX+Qv7A
F1NsCUwbBTg2LnNFkMB/xQSkEBu5OaEW5twgq1srwpLt617a1C5BX00/C5k2R+3aX8NMMQqWGT+4
bZ3KfYJcZpcdJvEyBYE5fNl4F40vOIi03YxJAnKwT4vKvmHsmst/aNkSwHoAQQa2qcmh65vhX++S
/M9Ev7m8UebMsoVz6Ws6vzqcz7doaOYYhSZVKdEhm/bn8UltR/cFvwMwrh40bgWsDgGNHWMhZIfa
toh604NutI3bNpfOp9x+w7sH4YAhrd8Dkn+/GqOVFvb2eDAaohUBjipURxI2JfeN50ZMwFMVRln0
Len8PH/gw6+uQ8uAZJUkElEkHZF/fNSkycmyIjyrwydAh2suTs89WNcAvpMi/E+SktR1/qiTmNsh
K47Zv9Z3wng6N4sHHAt33E0nkmgTDivhgpvadVYXuHPifOSt/X1+LHiPyazkc6SvotDoEudvq+D7
i7fZ1Scon67M4jMAe+A0MS4J4c5+WkcXf7AExrO4eAiKg8NIro8WY1VZkYrkZw3BuX6/cseMqeLy
M+scVU+GPto2g8b4OZbMq88Zrsb9EUJ6zEbH+LRtnA7U0O3096mLMBLzotmG8KG8XU6vE8009xu4
m4ST4KJEJ0gvHLv9yGgVd7sCIRrGm9Mwffm396tvQqdvpwgqQ76T5oUZzrt9mSS/8lZTRolHW9hK
UFm3+cS+BfBWi6NXmmUhV863PIJLq6nrlov3efnG7o8GGFVtqYInSHfnNEWwZj9WQZfSCCBlfrOR
b3vA4ERb1p3kcWvvFK4L7fRb9ey/O91NIP0SMPWaTJ8soyWim3jhG9OiycK7t/lq9tNOgAAmYWHQ
V2EkA2CFMAEMmDfEeln66rt0Mcbln1mOoUtqkxikAZ1HtBHOtiVlN+RnpP/nUysB15Zsrz54arCN
6FglROsjMgg1/pTJ4O4yXIBZjk449evnPFg3bCX+2raMqNRXL/jWQsBhtAhf63xO4snRvoNL1NZz
KheYBjc57ATY6RUeCeO+obGwcWi4Wn9KY4ODpiym3Umii0cILTOde1JhvBw2pkpoZq8V2sobDNge
RW9pOfEy5tY/b8AozuiRfhvzlUviz+Y6yMo3yFdOQfKWBPvdOGBkj1elswTrQZKzOfjaCEAUvMED
BWJCtSWZUJ02S00EeWHPMqOkyGhFSd5gjuqXtGYsg7ekUL05b8t7JzHKnFHiTWR6Su4ddUwGmRaY
PX6Lnzaf7Aoe65hj4hhoGu5kpt7YrrLJVGIefODxPqizxhjKPG71kaj4zn0MDSehFpCmSj/Jekni
hPOtWwE9yLL2KMaKTQgaKPdvbOuUuvL9TYPzGSx2XKZEuS46xKXvTq7mUrTdapCl/UHj4jgSsMSZ
OUUg0fMeRlZoTcJWCid2kXP9vLXfwevGWskBZReGFbWua1xTsBMD+MfRIPIctpJ9bOLnnfpL3pOg
9v9QS3EDmAQMs9Y16fdTHjZ2HxgSsxFkrbFS4ifPorJjLVCdI9jpbx4wnl75NiwzLZfn5veAXyfF
Z6bpz0izmuJ8ya9Sp3oHgMbKDe45RLxzLrn6Wn9Ue7AXe8d+gqHyuFJY2ZXCjA/Z4tliw2UXFoHB
XBjEptV2a1cLtSR2f0xVD0lAazELvgE9JrEzbufaWcFh37r3cDEnvCoOyhW+lAnT6bF6+Ske7NGw
rpzdbpmFVIquzyaDs28ZKxTyF0tC0h1cQq8Ap9dygWspwrME34VdmmjpFfltB0Royg2N6Lj90izn
VIOqzdaLLOFaGeA+UPFqX1hqkHQCPJgdrOGHPMGCNohSj8esKyzWJIMbIEHgjAqSN9pyCPtPMQbW
eNODBPPvwzW1XBUI8R5A6bbKpq0B5kl3rAjPf6p/d+BLpnKzfjCwmvY2lnLMDHH5imF74fuaQi6N
oCaTgWJRtyvwcJOJa0kmPtPdVb58HEwW797vrgrIzZ/ynzCQVgxvTi1wHWWebzKank+bgzWpcYRD
p+QxYBFOHmRx6k8NSs/t/Utu0dTy5Ver0dIeQ6eTNQtI28B206fj/3T5nW4SIPoQ28z8aVxrmg2P
R+/QXxUd5JX1i9NkngQMFcPITY1YkppKemLW9XWhH/qAML5rddW6nElkEm+8+XZmncOM8FC5PKs4
+lx1oeyEOcbTbuUVh2LYL21ICgnW/kqoTekF6seuS9vyZq98bwmrr9F3Hp180sSRvXPxdQo+4Nsr
9iE1BkhJD1toE5/0Ko9SeaF2b6lbw49GcEPFVjL7dJwuQBSny/aHh35YPGPjBSRH9mXd+dfpiUZo
jdfmf6Oco95ie5PwVuetRdYLk0rwSaYphb+MyXbkSOII15Fl63MIssxJlGnlz2a1cYstq9co81Nk
JenzU9Hhie/rLFHPtsNQQisXYxXB+ZqWMcAKCUc+//CAORTF6xwCKVySJQZ7+PTZ1YUQ2ykN0d9S
TyJVuwRBF5hIOKgXnNeZsJhwpFT56bIGhW1Lk5itYa2uQxrPQ+assSOqE/+kCTSo2dn07DdT1fpz
soeAxOBWnDEiiJVCPOT/a+Kl9TVEXYfpA7m/ZDEJRDfdvQfSWqY0ai4445V5ad2LsCGMO9jTpgpY
di6JnrwW73SlkQJz0revU65WqPBzhPk8Fc5b/EfOs07SCf2wKe0vWZa8rNTqX8s/9cVgeZ1wCyHP
mHSRCEdkffzV+6fspANJCKoSlAx75pYEOTaipbm4UuvJ1/R13U3iWXFIvrwDYnatTkHip9W8+7bZ
+D96t1QsBYUzSHeLKWfHzBUnV1VdgcTGtysIYv2yUsvOf+2/VcPdAzADvMQSU4olnL5HuLjzZKO5
A3twvqhWoNP4U7VRwjv6z9//y2oy1jMsgeNTaxLLOcAncgNcev1Uobc5jXZFak8GFWan3Yodtf6J
P3WR4V+PUbj3zxP2xL4X2RlL51iRYT+mG7j2GllsKvrWTqrQOsreMcOCflgTdtMMKK84kax09C4H
blD9EyX5Vy4LEU9qvYKoWB3Ib7JGmwSOh8GrN+QfFfb5lEvdNb+7GH7owexde9KitJ9L+ATZ+zWv
Yt/EBnNygcXZ/p2i+yxZ+muyip5HLCNOZ56vAFuKZyxs13Cx8qYtkkPRmfrQ8JmYVFO7f0+y3+Pp
990TZG0kFxWVeFcWYqsDyZbpsAboJmAiISIl7Ll8xnoUoKn+yHzu/Gm9wORtrck3Nr7X7KvwyRIt
Ay6Iy2zbnzaX5hY5MX9Ukw3BaQHS3CqLsdcvZo0AkjQ4QhQWMZJLm5uagKHvACRQLiElS1F32RUi
b2NP5Ts3iI6KwOwTsoViXglQwz4uswcTIQvbAWGlhXSasBB6xnVJ4HC7NMwi5Ejm7VIP8e5yQjHQ
RouORwhYhUMYLcJsuPiuGc3FcJSylABpOMjeIUpUThVMJ1DEy0Ujc5ikj4YdywdCXLQXOWeJRiLm
nOCKcBi2knC8upXYDXcVfvKCkdXhfOsKkEZdzF4BY+K07LKDtsSVdy6h7BxedlQffSHWBdSpiSEw
zqMf0kMfZ9NZid6CdQZzwv74EDeGbNJaSxlQ76uX523wmqB/NjOgq/cLP0Sh/wGQ7mA83RS/vkTa
EKoucOdbTJrH/L9MehYenICMw5IlWJvLt+6Yzto70ggr6hkwGGG6gcJDP3GhWGVzpCv/jbifdONd
rstNTF0P//rZswze8s2MJMdIOjSyFKwyxw05Mo/5KpFFkqE8ANoMfHEvD31yNXUddwGxI6rQAq5x
FyfYn7HxueZvgYV5wLv6SKMbgb1EFIkhKW/cpwDal5NkYQp5CJL4KfttSU47whzg653+QtNYhfCn
hB4OyzKPG6RQU2KWwNr6/ziwvMMpIATWZoIGPKDs4EvdMaDfLqJqPCqBScLGf7qNVDCVDYZXlpmo
4yjnLn6UQ5MZGjWdk9VeDYj0wNLDid5HOokWvyNTqPuTBOCdQnLm1DszK9kQt6nF6S58v8A1+qfK
n1kXrpHPg/Jky0CwxXM1IUqAkTX4MjVbkQ9v/gi/d+r2v5DQKcOxJX6TW8Mr08AiToQAP0g0xOGK
AuyCmoIBcjQaPYuD1rfYrZTP8cpxY4JUJc/wM8i9nWY3mQJT1nBJScc/P/crLO7NMVPEnsfynm2H
R/C25KmYRY7rRtKK3NldKPLt4Tw3XpEZTBTFNdTxsr13opngkabP+cbfMeGFkGq5oHQHGi0iSqMl
tu3KdgyqG2tw5Q4fqFwMPYCHAZ/6uGxWOLwgS0gLdlfYi/hQQabClhRMNqz5v4yDUmqlhln1lENK
xYEVzBeX1QekB9fHv3OMXK+0zlNf+68zs+je7AJLbePMe2SgyaLQGEBhHQVB8rcKFnoa5ZPwQbJF
naPYY1mVfWrp6pPe3wJpHbphZkJnClDZh5dp64/LCVSPsa4r4LrEz9QmZ8bAtsGGGYopqyIg9vmY
au9pirojG4RDfNhcbiRY2LZMkcXOScxWfhs5I9yW+2LJ/OIE1MFBhnkr6HIUEBT8IjyB3WZng4GY
IGrF+4R8gAE9nWxHvChMIpdEhhyB/JwIe9AHpLvO6BtHRBm5YVTBctMta16jBO0l+gVtp8JqZqh5
iKT0tzxzZ4SyulVbzuXYz++xvxOsIWmJL+PODa4RWkOU/iUhjPoPKfmG1w7WqKaWg9AFFWSJSUB0
ZwQBOHgLY+ukh6zf3J8oyAUK/sDrkSoVKIPwcJ1lHBmFoO1bqpG2Yqx2jEcpHbmQovCHDztSLZfO
+YvVWmzZnupuGb1nW3mqUmBali1cKgceMttotjE+qYMe8SRePW0p4isJGpz82Wl0TEptWo65DIwG
msxQ13lb12k7UTg6EfujUHs424hBnWPm3OhFsK5ZuB/asC2Q7Xy/ePGg2KRvORYiPXkGxFMSd11R
2uZJuwvSawvxUycx24ad42raSwJGojSCj0ihG1oJiCOxpXP869kn37NmJN48ZZwsXs43xL/WgAq/
O7TzR3Aks+cWTav4iJLBtwOS/gpzy/GW2LBoebgNKQolTIyiT1nbNjCq2VCZDnKU4tjpEnQpMgW8
ViX/rFKoNBWTRx+4yob7coyQisDeyJ/kbnBpgwCPQxeeDUS4MKnsKmw5XYmv/0EE/PQ0PMeoS7Oo
FmT4fZ7bNbsbML4oeV0h1kLdGgEqRLet0AwOiR4y8nGStHVgnQhHejthhyZR05vFDgQKERZL/ncT
fW+EFmqL4KzP6Vtu1RdGpBABuXiqxi8vEsqmBebrW+0k66Shi8vpFUabRk7cfpNwOS9GmqF5tDIc
bPAzJDigBIeZeGkDcfT4L0wjjN40H5SdgYG6KiOUURYqnWQEBtdajQ0hNjohk/81STE0W5gym4FY
+oJ47DDRafNRy/js41L7YCi9F6OSksk/7mEhZaNFk0lhlmpJSVYobtQZJ+OfJ1BVH3Ol8lMh71RL
irZ/tnADMOxtGc+zQH5nbAD5Jc8hLUBosuXn6IlCmqTR+PNB/gPG+rcdHPg6N/QHmBhxM3jRh49H
hfyr1Ewjaq6VpOoKHKM0hJIWsUMhDZZrvrEgmpoPq/qTy5MwPwBYZgxmUBV0ws5EhRtp4ESCLlMQ
0TwWQykjy76oJFwAxawkDZ+FotOiHkLs9++ujNtd+bSjqe3i+qghGkLt7XLpzyb4dyUjNSkKgTsM
VrTtn4QJVmwFCF/U1JXpieYBAjqWpVkFkEPD0JXdreQEfP+8XanhxEWHp50BiBmt0XA7tlusTEle
x6OSksmUvAtx+t6xUb8RId791VG0mCJ7venSjzKYmppGv2guokarmjtjHF0drObxmDStus2K4NfQ
41hp9ZbSLtupZ8Xb/RvjHhR8YSU+0/ZmRtO3k33gQOshrAAFTdlqD3dSaQxo7vr/BnqkVSCFqGmf
ogwtfg8GZ29cOhn1xoZOFGZK9VQFCWXSkkqnQuYp0LPI+2rbdBT5JxXgCFfZgvYIbraShDliBKdk
qRUd5t9cLo2XpuB3ggKvM2Ac3pghKtUyl5VyUXy0/L2+dvoLIBzWoRbAiv1zSmqYqFRhrD+BzmEe
hwlfItnM7lRsQna4mwrL00kaHYlEAqSHmVIq8kqm/sCEggXdO6wuS4PpeJucRunmEsQTssmOc+N/
72ubPG4nUU4o/tSsPv5bNj2XoEict2YOy38Blxrz/MEa+GtycYg+CFQ+PeQyqEegV5EsPzXBRS/y
+71vZfz/dl3ULvXFuxrBvX6dfdfww6ruEFpmLGRSwtkaprnISG4/w4ki100/RYhUEBHT3iZRvcK6
3p/MsQF8Zm5ncig4uozalz+UMg7WufrgeHyeT68CqydX9UnRJ3dmY3O8r7scRuoEhdzPC01aN798
pXQSt7vE90ucn+4+EUmI+q002J8n711qT4Kcw4cd/gFccTCf3NDq4Ka58HuUnaapNasGPBvCbxh/
JnHJDMDSSLOiOs07eRsQemTysex+eUUw+C+k85kliW9m6OTIPen6Hf2k6TwTGT4vnppBqZGq4EPd
gKZl4oBnxY0lk8Q7LnNovBS5XPbYAZAdCPv9pTRYn8FhTFoX5Tcf8bv1MI6KeAFN6qfWFFHjy+PR
m0Gh4h1woBnnTXn2xWKJZnp3pr2owGxuJioh6xS6ThHGr0iZNBRt0JmutHp63D9cUeKaxxNfJ9A8
wE7JLgtsjOMLaqiBFFzTQa/WoIx+ijgp/hBCfmEJFsvpIiu5RY6aKp1yf2s76ojltkaRos1R1/V/
T1ODZnr9nIAnRccO9zFpViWHnPu6UWaeWEpey9zOS9/a8mQFp7fv9I/9FxWZJZ4JO+WIUDct74av
4Cl+soZhBD8P7zqeFgNBqMN+QQWZ2uhELtoTAzN8MgqhF9Bk6I2VNekcUCDGq1VSnNSO9yyH89mp
qQgrz3e+GIQLUAMAR/huOpj1kS4PwnkIDhiUX8Xzp6axCM/tEUBgpsva0zuprU4etcoARuZIGHbL
Z3YJAqvI0ZT4/sUMARNzCKl8geJdwOrLRD1pwbsmwHKyrXY4FQu8jPqn4JEz6nP/x823TMvO1k35
cww2rZe6Tq2n7FUXItvh1R0uxuyesDHKxkfhKoZZQ8vWnklcyNri6oJPgYQ8E032PC3ykqHzQq2B
qED6hYEja0oMCMEeK2o7lC34ETmGIHkkbc2Z1ewJzB+CGmbbVHHv+OXjpRaafNNQws/WA8KIv0lP
vP/XCmlybIc9Q+DadVe91O8cr2mHkdOSCbDnBU1dLyHVjXwaKsN78FFJQfBp45nilOfsxlGUE8Sh
d5tzuqqp1HxfcCnyoGAaeAYuARav+kKoMUp7G5Wq2a6r+hCCogGgKRfHUUPUtg74CvSfiDdiDFHM
EH2TXyhsAwkdFtgp+ifctDQmXeXPZu7DqhEPn0K9IHNhtkWWowBBOqwMJh4FDp2fngl6rK6jHWY5
Qnfh3SGUlvcKpAOIkOrvt2uK7q9eLBuEg47t+gPRafZ+N2MG/rrkzQw+cpi8oOxtUngVx5HjUWEt
+FoU4gKuYkpy4bLWeMEANx3qyY67SC1+9uQX6szyUuKHwv9HkzqMlmd/mMY/Ah4Uqed3PocoE7K+
LihfcUC9vhtyHiHW+q+BXI1iRv1PF4sAdcOflAM75NQJ5dblEFnKjtplXYfiOzwA+HJi5AXu78j0
mFmWGwPekDjmhC3nedrLAvq6IJw2av0rWebPeyZZtnaTN2qJSPl59dlV0/ji+s9OcYBh5rEvEku1
j1XB+Ga+qaCirr2N5ta+vydP33iVppEEKW2CId4e2kvsLTTkCJUBnzMahQJlzpIwGk8KZo5356CL
kjQyx+hfTTheCL14fztw1mYArv3IUaEQ2RDgn6/OMZJ6UXX15ZnTnEF6kJEF9tdZA6OQHu4Go2sd
SwNN7Fihmgj9rkpruqxKvDDXITq07jdKK7wOrOHgfCbdZxKwVOnUJ+STN2A9PdBKqDBcISty8LLA
6FgSnR//cM3bsgtSOKb9XwtOVYWZB6bKp3u/R4G2pyajYgkDSDYGkx67GXF6XrE/hoCIXER4j0is
gi/vX7lBmzC84tGJJOlE7FfuouzjjohICAg/rndkGSTPN+AfB7hR42Lh+omPp0gMLgQ8IXwfY6gk
SikfHJKOkfxU2fDQ4pscFQt5miy9XeP5Ff7K5oOh4oKQpwYDq+9C7pi8zlffo4xjM2D2o3xleTZ/
BTKaZfcwkwOLQpSn4hvZkDcRQogbAS3IBGcp0oQcZ8e00rg8K7Zo9fnYGk4JgTx0n3Gc9BAyUlim
MQaEKwXlTd7NdJRPuzX49XxUD8WMJzAnhG49Yz0OlYPHDPZ/bTv2Yco5jJTnap23JygcOy5dgILV
Vkg4TBUwWKd7qAGlwnTdWfWVlVlvf/6Ivfmd17M6KW6Mj0tbT7j9859m9cO+ItK3uzfWuzteR+yB
iVc5k0nLM8D+6MjdFCA3u++OZAqO3obQewpVREWBDDmxdiaRGAyX5uD8ir6jytyD0saVqvHg9edn
XXtY8UbwAfLZHOgptl0395XJm/+bY8qQqXlB+ObxFv4Gu98imVCSErAWRuUVGQm4ZhGZ/n0BtAjn
NxkEwaIErd7CBkNQ3+J2uIA5hTd6Tg7ZR+R59yDqp+HjR3thYDOxVJFbGDXYUoYXmot47yI9xzsX
nR5W85F3MLP04i1nopdENpUIerd5nvK6EsE19f9ZAC0n7JnMSRZwcJE/LrPdXpm4e2+eh5F2Wv66
/OU+/0JcHEvTs8I74b4/uF0hRD6hwrB7NBkCKUw/9/OJfymyhT+3rvFMVBF/j9YbVMfuT4E+OlwP
/2M+97lZSRETqUu400u+7a+1WbPMCJeduHNBb87BdkxIaqiZExdqp0tEimOnQ15RdjYL8NtmFMjd
60HtLuxI4IoShWJKHluSgjm9c53L2+CxQ2alWv7/pc4zHIA8//RmZYVeAhfImdGZoWN/XFj1AWpV
wsG91yODqojZ3QUcFN0AouMSKrh61VmxT+25UzVLc/T3cMS7skkE0j2vS7sPJscR/ES2Iu4znZQj
zYx20cTpK5xjpGAMurwAah6ti6tYHPMIarJD1AQcWYmr7CPUefg2XDZY5cduOKeMspQf1TH9CisJ
GnenUyjaEq27zENh+NSskbzaZ5+GhqqRcIaO+4Q9F1p+HRBQg8cSGqJP7lj1Ipk++fzwbFzcGZY4
dItcjD1IFAkyuvUJWiKLFIYkd+dwmA0wTZDbuTBYAnWsNuGsOXJRuV2nSrOtuAx/mQtbycyUP0vU
3ZW9Bt76TmKhI2twUi/R8KfEuRSw5ifr0jEJk8aq/yUZTYcYQlfuDENbfkMNcZ1tr7sC1J5JIU09
huUroilna5dXIPl9l2hBBhPvnzszM5fB3cAVVTzNR90LX2shifLsVZ3Lgh9BxM1M3Nm4AiDWkeN9
fo/R6nsuLypwJk0u8Z5JH5JTSvD+Pg8QusxrajYnpKNzyu7R3lNiFocYsqx8xuGXFrBTGkwjJH/p
dFtOyZIxXAgQ0Kj8tO/DM7os9BsBDuN4A9deybThm0q3ZoXJrq7+j8jjeENhkAuvQjwaSdX29Urn
hJ/oAXkMxzVHSeV4CTZLTp0NUwXKuXy7Bx//uKC82TvOXbidGcWVj8QeFwUbe7zzBgsANoe4FlyG
ReOn2TmEsEj7a1HJrORGjiq37Z1AcdTg0B00siL13xLCWI4KgU+w5neSBk0zux6qKVQ7BQU+ZqTX
nXwqNuH07OLDKHf9oLTc1aN9+WXXzTLjvMHAENxuHV0EU9Sq2RoywMiOQ1xMgfjhW4cIDBY1/Fpd
20BgN+jwClT9917g7s+LbnebFvKE7S4tjobroTe0I1WvUSAFefSligHiVco8JfTmwJr1FpRYBpE7
XvXqEpQFpbjkqz0quJsglLw+SfIWQDVoWUuF0yg7/CJNAnzEfu7l2J7ZyKg1FTlkpVQLgSSFDZCl
uSKALfiZgRopkisV09omko3FsWbeujq38kbWew7l/NPsSJdrP1o1/LzlEf06V6313uD4KZDqIJrE
akOB5HVt4fjuK+GuTnFQeXUjFNXc4C/y4vJUOSu/cHy3cz6Z8Yorw63iucrV5k0rO1DdGqP1vYKy
AhZlgnn1XpOzidEEZtMubR50ibizmM3GPCjoKFTmEni9wnEsHel74gGx8fLocnq6oTWkw34xUcE7
jn10wXsU7uUvfYmkHKxk/0QEHMfconHwdbjm6Zw//vPrCso4r07U3DtjB/6fp916Benn/oWCmhJr
vCvHPiG9yHluO97s+F4URI7S4J/EjLbHX6P3Jx3xlT/WS4Wp8gkTz0pNKoy45TBir773E/4pUtk1
wm0Ht2UO1awC5Uf4oucMUGCake8sqoTFaEPOc392UVsEBdiN23eB6jNusvLnAw1YIXoKo2vq6yfY
kQSqPRsBvVQQpwkWLsaAVqghZBQlxBpZiRG0Pk1ddCIoodnZ28936cG67CwuHguNzphEEPmU+58g
oSLdM0YDd4ABnDkYFceQz9V6a/W1qvlq00QzQ88efx3lkgeksHR5tKoiKvLCewgls0p36X9/5iGg
Z0bk5XOgrtHdMddrfHUSYZFSZdjEDfuhdMh5THI3OMuPE/TwLDOMTCI9RkT4BLZ1gS5GNB0qAP/R
VE7HVwsX4JuHVbfapr8QPVVzbEUZVToMGsEoTrUKMpT/OGBAQHUQKAK18z6EQqm0uLgCtY2XW3iT
UT3o6pJobh9XP7WeucjE4sx3SiDeqG6HvXFkfDC16U2zQcYsHMw1kmCsoHfhFpqnc8bUpVV8mTM2
+hln6td+hmHyeUtN/4AI0YLzOm6/dJvp9W0BmeDuxUHhXHcqFiCm6XqCSgiUx679+NFCoedBYFil
4P0+kftZdJbVAVU3VoIVizosRFOH+A+nR7Ogv1lJCruk4cOEgCOJa0WMF6M41Q8sZEuVeS/fygHN
y6tI5ZCasWM3+eTqO/NHRt+RK/295VUmG9hDK3+NoZV5lrtK+osFB5EPO2IeJ4dL0dcxXJb1EwjB
I+TMNyK6KKLy1X9mJXMp3Ta9wk1vv6Tmv1zSMKaNtszcGtRd3TvqU1dwEWDoS3fZIrIIkW/8dt4s
7Qv2/nGspH8Xr+wc8xEYv2XJMcrOrBVJ/rGV/6ZRY+6WTT939n2EFqIY/hNYxSIVRazV6qTohaD9
f3Uad3CzUm0Zmk0TXQJBRhOtMTkaM9DdR22n3Lk7GmnrPG+awV+SeX5kHT6KKvBB9W/2trY5PLQt
pEwnMurtB+s3hcbi7shC/2ZPc00S+SmYVk9EWAXYmutSGeanXCtJCt9zyi6d8v/g9+t9pYt3HZ78
DnmpK87yOZnEjrx4w+ZVkXJlnupKBW7mzcE6nTcu0bliAHtoQQapOwzNApbmhsJh4L8wcCkYbJ9/
usrm9sYbrwRqVbo1/fEX1p/OrBcPr5OHLyg0HgwdpJzDdtyEgp4Bblv7hDfskBFteS8+zUraSR6D
sNwzLGKwM2Y8gBmf8byd4DFoNBGhKTf+z9uFG/cltrwadQ64RFYera3rS5SeyLd0q7xqG30l71P/
gG6+p8UZ1ZGeTCUkhrU8W2sTc9TEKvoyk3hcEjqG8udWMnlgwGrMG4MOixlH0822YavGIDmk11BR
uIvOqRhJHR2uV3hlPJ4ixQfuUpVXZzHO7p0I+HeIaxnFwjXHof8ObViGHJVXw4OQX9Lp8w6Ejwq1
7yVc2UefMDu/SBFtqGb81UbzUmIHgX7bnoPKi16Uv0bju+WngYQXpXjoqPSSH35JhK+5gjmHsVHL
v+o8+oN9ce3fmgLEKC1oPp2/VGcIsOHoAjNJQZUjBbrJVfxq8g41/1d/VgB4LbLPZ/JMUAVQLXl8
HnwEiZSGo+h8reYYz0zgmzlVRc/xfoDQI1kKojXkDwrVd0hlqC7qiMO3ZqQAFsXK8ztUIspl93oz
uXYuIsIyb5KJ28tiTtPIUYBf7s0x3lzupOCERB3y5hCVfJmixQOHAhxE3FS96TKgrmTJzhcl8im7
c+aM5cMd6+KZf3OvrZcI/IeZ0pgOlmGJ9QDZiPG38dgbAC3rVWsz5Kml4S4oBH8ZR820i93gh5Yl
ZckWG3GnFmH0ldnaSR4jfca2tf4MVdH9WKDYIKQwUtumh2rrxZpBixMI2i8UXNiDfgVCaRS/Z4Sc
yIC7e8AZrjvLqRMBD1WlUEhrSI2phP3rHUCkFjyWOI3LEZXtAmQlz+mQPP0epfFLcUimzLfbnloq
Sckm4KWtbm7etZjOJC5z47UlLTBEc52J8bCeU7xHiUEGAvGXuPEX/DEZBRnw7N5NxCkV/y7lJdfG
lNWlb80FrzI1LsIPNgJVHHryDJ1gAbPE7GO+6vuxM+picOanb8KeuhPqiZYQsvFOJhFI3TQKnY8e
PGyjVFiO0Qx61pdo0SzOtQ536kfA+puCCmjCiKir7pUEFf0NsBvTRIauwXzJdOEXoVYTFCa4K/uF
JbjUOT/KjI96hs7nVG8CiHpHAQrbmHnsv9izd9O1u6+5LurXShfijGEVi9tbcCLFD8HxjVfhO6GU
OxAEurAQNotDi2ch97jWWjTpRG/C3iPxIsAjRcGgI/tgOfvOM6FkyRhKm844LcJul/sLnKQiQ8wR
OHOOPgXpeNPky/znOErpFUApZxPr8paNvF2PeEGB8WBIIIBefCHywgkGmbXZAPDtj6GXInl30zvy
ZMp6d0KWFIALyQw+4dRmuH+GL+onlre8WK3SkxVWOKDlQMuCJw/Lc60knUQ28sZqDCPgp4yx2MEi
O6wgR4oIPfPUSdhgXI6IQyLpdimEPBuHuOcq4OJg0lBGPYceSl7oSwJFsJv6c+6Ta9Nl2I4GyC9T
+nOb4EhP4cPGo3dLo5KjvRxyepXDL9GSnwMqCm1jeGrvg1YDANvIJb5MlKSJcct9mvvCR/tiby0A
7mlgu+TDL5QexTI405k52rUzbFcKojptPZIG4E7Dlsa+QK9d8y4k4kOidGa8N+SVPPT/LQcN81nQ
pBDKbrN/JoOKtPB3YpDsFTk9l6jinokOwWurURCChILuNr8tBTvUHLDZ2VA9x92OJ12fGk7xaya6
koaDSzF86Fw0RZrF1Qgc+Oqr17dZSCN+REHjgVembpSowifw1YEUIEl8W62OU3WTydYlx4Qvk7hi
8GPweDWQDGQoyLe+LfchVCND3Er3M07dlGMnyahBYRJoW3mYxBweubpwoUA/ZqK5fBZrROi9BZ00
X5tHkREqtkIw8b8ucm4Sr5oemRo1JcxvTNv7L2xt5OLrvBWYejrdDTyZtEdVZ2zitkM/U3EMxWwZ
3/TMfBXdNh8gxQrsgaC9Eg/sJ/LcG1rOINnyqUjwAQTKWJIh4daBuEXYkJc0w6K0Uclu0kVYcBk/
ZjWnvY0phA7s8r5prIcvA67Td+KDphxOKmagN6NyTBMIiewj0/ir4RnFROoVc8OfoOiFV5BGtw+z
o7TLZgLfaLX73HeEJ3mPw1GYqYUP0zy96KL6kGTl/HvNJmaYp51lxjsChljOJR3z1fH/+3NaChnI
F1jr+40J4InM/bXrXopzPj7W6gnM8oscU+s5zGV44UDQdkl8TvhaxPleu42LQcmjDAgkZQG/7/GU
wxPA2czye6tu/ud9fQpbPoJlMvLqNOVvL/mfS4IoPUyVoM58p/0RMF7/XhrXKOk20tH+pBbBudOG
XyEUHYyzdwNBK+xHmTc2NdgcmQsjGOeEn2qiS1bivjwPSJOT3Z2EvABYIBDE/4x1zj1ELd6FtesW
Jaih1HSx542O5MuQyONpNX8etqlqf5L9h1ZeO/zefvo+pH7VCvwVGqIRTr6+jZf35pMD+KpOi1yn
WH9O/05CqCFtKu6Lw9AANh07Kwp0Y4Mw8ncdxOYnwfEYzob8uyMDJ/qg9VCjBYJqq3bRf4JQJ6Xm
Us9wwEZULV2r7aphHb83+5C4Eepl2ybSjGSyz2A9ReDRlI8PrQKzKAh77VJM7ssOJlrCHvsAh6WP
zm2OLq7Uys6esFTYAWJjMXVCNyMuYt9iaI9r7qwiCnacM9xwCDazdlh+PhXcm9oWR5+4G0uKFudE
wOG3vhGEeDF/WFpoYfpeE+GVIw646VbR80t9rDVNo8hDNFjMIRhzVL8JeqQfH5U3XmnF1DgbeCjc
jeJcJMrOol9GtbdHSTRAMu1rmyLb6t5Qj/LRYdr4MBbw7Fz4Ij0Jk8e/TQ7U814HROkOTRuMsdzq
YIaXAh+xRqN3suDhK3oPaLVS2sqYOJNiKc6/hwit6IR7UQEt3+nDViy84JKjRyLBIZK3iSXVAuyx
cedygMhpg2gVhNIysCB3M6O4J8gLmsLJD9lt3Ctvwp7P+kLF9/UFNzWqORTWKLlZQRw+q4pVPd0f
KnsQJWeGBvzTAaPKt7E7g3XLsr0iM9rcXt+gKF5g8IP+DfiqT5nZqAIna4TaJQQm/rncYIY8s4ih
bneaXSquo4A5ALvx5LTHK50+OHcSvbgp5gJzLyeNlyUE6rqlajebBoVSzMTbFy8+VWyaHgSU0C+Z
I7Nq0gzc8/y95Wyu9/QrXWsF0sbGRZZraj5m5jLy7lVZp2ZEjG6b7zKZLpg2Cjl2cCCOkIOfc7tV
JH7/prZAqeCTph+sv1qZBBb9prxRJoJE2QPW+ldQdsfwN9USIFwj1E1Yc98wb3XRfLKP58w1Q73f
mIAzldllnYhUALejqepxZYUNMAe4CiVHUzMg6yR0icSE/qoPr0dgbcyTTadomdPEHYJ14w1/DOry
uxyr6lrSelXul7chRoqXNLedAV73rYa8VaR7r8Zj8nK1sNTW0zLcxm+f9qkzzeOoF4jCCl9bcoc9
nvcXtSMM5Pu/eoZkVh4PWlZCBGno7n0En8SvHfl/Sh/WGJMoJeOsE/1bCcfR+Pb9K7+snm3xaZSl
itpRj35ddznSMqjwirP3y5F0/+daKifW/3kuMdmh5QBI7vFd9VqUqvSOq4Q6e3m8A53Rma2EAccv
KQMt+Sr0dtGwURx0z7qycuGyj0O6Zr9yVgacK1gcqmO+1/KafTbuDd1gsbuSOlfvz1sfkQ6rUjqq
kKUBMhSe6+pyur+ardP9+AmA64XD4N8Tao27ghMI8xJHeEzqZqXmQxAHwTmezcqNxZv3RpgM/ADB
nBvvhPYI0dFhreojLyzN67C1OuTBorP78wjSbW0FW8UmJf0xuRn6pUeTJim6x3pJON0Pq1z11D1J
1FeYbcoJXVNZ04u5fN52ja/jWObMcT/Jukv+dN7+woBu5TciMBRauVVbVPn7PT9R2wHwziXLfQA1
+11v2XuesAsmxQnUAhxPUTkZ40DobgsXpi48PD5gCFN2yWOuLQh9beIzhU3aQBVOHu7ILFR28j9r
/4grb2CNbRrXV2+SeGjVnNjWLA5rsRlqzWmpAsSYHhcrj4ir5Yd8mi84R8g96mHoHABx6xmzO+vz
+yoQRgSE/mftKnRp4ZqAXe4EUVqAGZ9vr6S2sAkTBO3bVubwKgVHVnWHrmmxT8vuH+e9NCJaTMFT
kPP7eTcdPfmB3iTkftRqaWvsguuIi2okZ/rgsqSJviJap4RminynLF3Y3EYg3spigjKZB3B6Uatw
f7tH2CV5HZ+H8pKPAg/dBvLxVxGYUVtFpgupwp76aWafnD0YyLRsyRnf6R0e0zMnW8LMKc9C3blK
dwAT4weOlUd1SbqRjelaa9u5UUV+5BXw9HUUmEitDXR/zTIN+6gEdOUpRjlgmTbstNNMLwRD4VlK
M6G9CII2dkNjEWupOIVXcyMZxPRNLn8fo8pU55HTUjH7DbRoTQ/CAjJ49KMHr55jJ087U9EtsnfL
dYFiaIE3AAwCZ0grhDYWjRp7Us2/Gq1rFmbJKCjO92kJz6LbuT5FQ3rY4i7o+xdOF7oBAeGOPdIG
d0fYON29Fgps+xdDc/8wRtrgtCO523WvgjqfV1InLkmXXikRnLb1Nd9fQRCATy0fp1mRDd0R8hvj
AeIoQ4iwnPuAO4L18ocfozXJPXxEQdgE4wdmZeNZK1sANahyHDX9SI3eoB/CUsPjZ3D9YiIaRi0F
OXQegvt6dzddc9gEsDgn7RvdzLeakH30zmMYU1Mceja8eEMcwoyEoDRBSqtORRDyeSmGkBzRNLop
dlvqw79eyzCsjlXAQHr7ldp+eET6jgcHj/rhDToVLItKOJOnxR+K4dpSGJtql6o364yEyqiX5nsv
H4MSnxO02jWvqoDaC5GsTFWMKpW7FL9P1pdtAiejl+tCRm0Qgc6l5sZROqlIGDHoj/PeGbjJMTYH
VxsVnmDNIfQ7gnV8O8vnpdighMcFmxJbBeOUEbP6y0QhyYbr7OOukIrdGFGtXth3T19zfMpB3M0q
I0hdH/W+kD22hnU0opDACmIcgMxZoGRVfSmg7PAarXwAFmT3BkEl4pc6ruO4XxVQlFOg1PO4BUl3
0UORwRjeZ9OZSk0RY8Yr9t7C9C8v87B6c7frlFUX02FwAAfIeJfZInr5cfp14S30J4l4ud87y1KX
dUXVRImUjvHzu1oZfFficZ8MG+ybzzjPg5BPQIGqUOKsGBAxbGFopUmwz0OziePzstAltOrYHbwi
fvcZI8UNeJdn1hM+nevpDJ8Vbt1HST0GP+KKvMU4xG1SOkPuN62Txw1vIWrFO51kAT96Y7nHN/0Y
aUX5K2lg3yn27xLTE3/yiGxhlXLIHUmKKqgmDmpUTtwLV1i555VeNeTljrzhGovPpc+Yl9k3CBgw
YhPTPm+mKswEMo1vEmjYTorNEWXmpWlcjLK2N5hkfNOt+dcU02rvND2EurqB9I4FE1KUbj+ciCSS
RpczyRfSZOfBlfxxpzhMOLdyrlabNX4w796Zt5LzFUGcxSCIo8aKWuvciopr4BbeVTiSaWqBj4A2
LmF88QWPHUl3XexIzisxQvtP0OWnSgf+hu4MGvUM6wt0g9RYNapmdWFnSCO4pxQarBI6Sax4A6nJ
yAUmhVMh7wez4GpeaUqH4jtYPjR2GHLXRPxBTWDTaZtM4o33TFU1lHwRNnDvrKKPtMcXHCeELXLR
If0RnQZaqcGTCNsUUxDodPnKkTRBtol4Pq+Y0uBfZUjDT5FaSSgaRqtSIJPrXzt3mlUeFBsD7Atc
qLFZYHkJSPgrPYENQztK34hAUKMzyK4KISbHZdJ+40VpDq4MoZYs1xAJPsVAjpkmscpIp35gnz2M
S4FFBgYJxEPAW2OCJU24ZeEKB+oDuq0kzsES+RO9zhBMME7rtEWtv+RrI2zZwL/pyin4XVFv5QFS
fy7vw6wr1Zp4PDIybXUVN/dSuPE29LNowEA4gtyxU5o/QIJMQ57+PBStL1PGhONGDGMvFI+Jd6vP
pF/LzQltf5z/gdG+r6RvMJ/y9aECEYOp9+zUPzdhZKEAkGj2UVB9guSzrzeLV0gwwA3NOrTlEDD8
QdV/fG/9FeJPJFTpPgiZABLyzt6U0LemJ6zxcilwtXIOyeEF2v9b8ne+6hWvuid0ShLhpvBKcihZ
UbTvAh6Lry3GW6AhrMaACOu6DUgySyfd0UXRS3MGbHX7IdD7Oydptkweg/IsUMm6KOPTw8Qp2bwy
scfBdsFhsDW3FpxyYmouATjdNdWlzkIhDNe6o836hYPiZ3xy+tifJibxgyCeooQQid0hXc2i3+cJ
KamrjFPi7zH8dbafVcE3JclRJ1Olv1tT5Kyed2rRwtDb2QxVp2zCFk/8jXThbB/FdL2Zui8zlb+R
dV0+u9MYy2NRuqqIEkOTnLy8kM3tal4hsGfxvVKUg7ephoWSpqKJlulGVzT/D9qtGu6fO9scnYFC
4Zmfdez32YTsICM/uYPpLb2bdRzCiEBqnkyKG9yg/5shlUNVVV/FnhxWNwzAU9fqlSO50/wny41x
3Fj93KoLStLQEQdcL3iP9ju0TOslmb5sywpTHvT0Wgpx75vn899tUqm/3E4HSIwf3rsKf8RvO2hc
J4Jp9UhtQwlQwEGLNI0oTj4ONPIvTYafQRLGb9FGGA0AFS9RSkij2pHCT7yZE/aMfiKVYYFpgw0x
lviDVWIk5wZbQlyOj1bXcAtAoTLmcxu5YfDQKklNnFxpJkXhcSBFlNJ0qJ5HQmmim3cIXxjfnKr/
7F//VvRrclaVN4QD56OFQxgnnlr7bDRqOcu6PGAKeUF+T+W7Cbq6b9cYRVxvSSaN31R/lgAfz3yI
wmcG05fFVRKVJ7mDZmbfnZUyqXEZ3D0P/rTNi3u6/eQzb1LOeO76NFQ7Ue1Em7QEhCzICwD/sMZU
rCTXsrJ3zKHS/PwVygrSoDNbq20gDwA5VeIKYP/PVdcJjp1sJ9rXLXH+P3k+2L8u+UjaN6m4FVaN
260an07u7Y8YdevSKa/djCNTCo055K8fsLnSfTZls7TzJkqBb0RMcn59ykJ5zMLlp3nB6sUs4Q3H
218L4gvld23Zi9DdvKJ4Kf1PVD3ODDp6FuqhDIsmAxP/9eKHwdlyi3lpsqSVF5sS85P39fgaSWVG
hc7gbSZpPEaTlvo/vloONh9CjYMUBm6VdJcexVG42LuzUZSpr2Cn4aff3AHXArruIA3g/0kwPYrE
k23zTYS/FOiRYNQVyJmmpkR+wShqRU3onlbic6snEB7VDp50gavnisnIpc8RQkUIxLK3ESpeMvut
7FXbnw5uJ4k70FpPTk8JJVaArhoZNqo0bt4jeJP9ECaow8L2m2+DOvXIpaF9o5g3Y6s0wN3UTChQ
khYtfXdz10UYhe9SeXX/duruetKOeXjnbMLOtHioXJPjMCyzRgX8YlnxBq1HPEqF5zzmWtONuXE9
SUbORg/uauLXdRrBEVFtpdaEX50Lzl+9MART5LmwyEsBbiLBUrsglFcalwjDBk39b42C3bkL2W81
JM9oq/jNRjC33kqIDIxAdkBVtgzGSWEpd8vUA66O7M4RN17jsfv+wlcV8lreTjPqANRaqGPTk1ty
orQS2JYXghnmmhboT8S/dpp0qixwHsJA2XRXSMMCiRCCXbuFPWY/M4w/UXGBi31Zddp6/fcMXik5
wSbXBxP3rOaOwzr739uHgUNNk/NT16X6JdB5BkOe6SyS+nxz7ZzzLf1B65PDv7FfJO5MyAv3CZAP
7RkrYdmluh58ZPRHT8iPzDGo0K2iVaKpvGr4Q6niGXtRSdqUeCP3PATGOrBQyOUNxK2k5X6BunM4
JUx+5Naiks0KSuNgrbEMLjuMtb62UQprkmPwsBEs1m2pY1xPTGzr87Ow5jJimUIrR6Gb+MX0XJvP
SL89NAnpjeJwB6dxndwl3xBxfjA+5O0G2m1wYtFCeLDEE9JFCsOJHwQ1/0VoCnEBMmsVztbg7f8E
uO/PouMTcpK17bHeP+Y6BSTdd47k9aQuwlNeZkLaZ/y/bGEdy+1/F/pThCXKdaI+RqOfmG2FmXgM
R92XU3cp2LL0BKzOIZlVdNtq/Ng+V4X2OuW42orgDVK45O3gEpLKUCG0qlVSXAsgoHN3Ypl1rGMt
6J6eAHl5vkxK80TJrzLOJpY6JOrlf6FBYLmpke4Kvnq99QHEfQZMbKA28os5w7FFvlAjZEKY2XDr
5hPhi9bbUSLjsAaU3nFcLS4wLqqvqncHa+Zer4Y6KZDCslbfj0/bder2vxB5NbDkCC2rvJdmB/5n
4YHVgRqWPee6Rv3kAn9S/9+y+ygnaWP75aoockV7QSBk9+gX64MmdnMNfLOw1MT4/mxqYSYwjEkI
R/IHZBpj95mh2BvEaG4VEWisCLIfkjt2CpXJAnKczbn8L5jNMHrDCDSvj1jvRdRvw3M3X+B4ryWx
x6spxjdLo9WbKj6rg43HkVqhXGTKBbBxK1M57czTBs1YrIpccxu2gNMKt4y04wtG/YPRuvrS3BIg
6Ci0H3ok00xJ7D7DkeMkA/dyGl2lGKUdGLQ+G1b4E75mgykOFNkT3f2YVP4tQ4f19vZW4MJOF2WS
2ACEqJwBRQxvAqvQcpB8V329k5nRtZAJoUNyvxkNEiLdOYR1WJflsBk6mAYplDrXRx4ZlLMJxUSp
IR/GezsH8MAyl9BQhK5XDKDI/kRdsIXrwfStZ83AheZNksOg+mst8SvYzl7LrLmT/d2taY5e0biP
p9jzUe1ENaiRQhgxZ2EfPK+++cC15+9qGICG1N/u5AoZbuE/5yHtOGQKNiq5uWkLWEz/Fn37wilN
W3J6vywB/ZoATVDC87WKfAQuYHjUOt7fn5m5fYDHCwHc1vPg5LTTf1L2r34Q66kxfAU4oSXxlNvL
LQBNFRCq3rW/SR5xLSLTn6igeb5En27b0VPzCPRQOpqQkD7KQ9O+Lyx/dgxiMzw66oy1cmqB2h1O
+DBPOZb+Ys0YRKs9REXCBaabHzJDijxsD/pONExVmEDN/Lkqhgy39EAQt3Vm623KWo2FFBlq/+hb
G2Epl30M4z6TDdT/QCzdTdDiGU18oZ2jtWJAupBRBRgzvjOdTr0Szc3G3YLE/yNcYmk9YF1AOs16
MIKk+xmBSHOorPjmEMWDVf+StAKt+QAN/eTbPFJB608T5Tl9MwHznHCPPcJRlXwwMY1hGLbx4FzI
HLOlsiuoIu0R+eRhggNFBpG0ui6mYupG8Hq2Au5UZIVnKt+1MHsjA5qLcc5yqQ3XIeOArVRcJ2h5
jKWFcJa4qYktCAdeJiSOcK3/HADz6XVeUpV2dNrxtphhNbMVJAAvdEnF0F6QHcVjeNma1wSq1eJe
fO9Y5hx7rB6FAr5+iC3AF44VgemxkJnlF166+8bx4CPcyXvvN/RbU5SwsnNoRRLVJa13+ElyTr4s
Ysu73gOhrq43UsMjIlxlHLSLL+y/oL2RwCK/mCwzL341KoQhHSUgV1TerHr9nWFtfsHqAPDAeO1Q
bDpOo/nmn9a/DZNRT2beA09tEyDu+FjNYQcnfRYyhxKqwdWYfVICCW5Vs3bw6Ix59ZPblNGisHT8
avAgg7kDIpUr9nnIhg8UpxZe/ltsfUhihVxAobbGOLAbPG58Gx8GSdKvFdUSNtBMQ9A3Zv/Vfw8J
253xPPG0yqiZiZhGFd0TFekr7f7zgxOjsSltTV03UuyG5JTQ0nRFJU/yROxWBfoC6aSwY24rRGzS
w2aixoYTuf0dcHl8c6IIhYRmtFF4iQ+8w5Ghth/REzhajniAk1WxbXhxaAUyZB+MkZZbLX2P3szv
V1RIqdNk0bMkYbXtlznLxdwEe1eGhGkGS/k/ATo7za7yElpeemaUhufFTgXzyc2Uinjpy38A+vvt
K5tcu+zmgSYxv8wRR8JYi2EAVoMw3T3MAlx0aQuuIexu3fnZi8HU1AB3CS22Cr/jx5+XDKOfI5NV
hRknhKLV9FgJGrWAtNTBMUQp/lVsMggVkSasF0yrjqBD7yfRrBnuQ0ASvqvog6VcZImok/GWjmXm
eYM5bfbBWkIRufBDmU7A34itsEZtbR6M0N5dPpgKHXSBSUbk+7aRE6StGWHLc8+9xp6U0fSGU5FP
xt1mG+v3bkd1G1aAENHi7l5Bm5ItgW8XeaDXjp4bKJWqSTEy5S6B/tJl4Zn18Oo+uq7HSZnmgdQd
KkL7cJmWzKZKwsQjuGmAlI+XiAnxIb3KNZMQv2G0yCOAFjLimz+m3Lba+XMrzuebSq8nI4vcmM05
ZNi242KXChNFaJ0byAvd3qQBRdxABgsRpk58UI61ocepyFP7X3VwKYh29iQ2Vo7bYxsoEKRaL6uq
EZNPDDpucBU3sZQz1JVy06/DH9guuKd80fq477pAI3B0a6ZluvYgfZ943YQW2ASUVm+e+e1cVIaz
IN9NAkrCsK9yXzvCsRwxfplSwG93PBtEVL8JV7pZ5jMLDg4+8UA0AmhvycLEC5uAyjKOymdHMNKy
bllKHEOO9abRr6v9NGOwgQbnpVl2tWN6Mzhn9qE8dpzqZHOn6RHrGUJ01AeDgOMbIv32UJ5DtQtC
iytCLMxduegIT+DR8hobtc9cVrUxRbhCWgQl761YxcW9ykUnayS6+eVp9JnxozEagaYiUFJPYjGD
ZOr+iH454zMMOxTlvWAH5w+cwpbuYG3k5e4S2JFMmbxrvRV+jxOYMeIXvxVhohZo+n6fX9IBG2Lo
MP9LpYeLEHqRf4RcwETOHXQdHJ/2jwAv38YKDCYWGevpceVM6j/uEeETO2iowP1D4r5LdZ0mpEw4
9equwaeAG/gPj3xOW/ai7gSqj9V4d2aJQjQDth50wPfBrKMX3FFQ9Q2c9uHaafXLFvj5IPVMfOWk
X4WHTImxtZxauEK3YFcPioVF43nio/j8ATBz6HYLdlfjL9x2MZ3C2VQVRDsQtrk7YK6jmgHe3QeF
eiN32FoYzBZASZs5M2Zjou098O9XWpwR6aEthBuYYJuteMafLOX+PD1q3n9EhdStJ3Wh7gmiWq1V
7fvtMtSUB2cwwntbuVpixH8IIQcaqgrcuTlfA61aH8xXbhE5Z2LgZL0yoIElQMrgeAY4tuATuXim
TtfO+KAIC0HCcjeKagf5eSWJziastsSj8XoNUhL/xWpzW3oBLqaSUc6uhOxwuFrAh3DlK8wVj/VK
cOvSQQ0fbsJ3MFGyLAE5ytQXU/biEQyqWpaEybtMYznU9grcAyiNQsEFUzoGhVxnOR0EJ6s5qVod
wyyE6jTIKU9mql/JKG0oZxRgJcR8VbJGnt0A1ZrBCBajHuI2TPk5FvTmFvBXkysDEC8bLvMCwTxu
PhuWZ3LvicKgKvnZ5lOTfavBPH0sAPMDrza+Gze1UwyYQRUQDkgO4TCHcHtIww5MsFxSCThQxa+b
cx0SKC3CLim1LieOnDi/WEbJ2z7+3+PnqiHRNSTo/IfWq75MfTx6stJU+Kcjhn2I9KRlpkXSU6tf
R0LHpcVxAWcC/NuWi7dIdVl3AQn88NDxIYLrIfuv09Jlw9mh7SwGRR+YHorgl0OauAP8lJDPklBP
h1NjqwDzQ6DBmgC3cyzO02icB8rcHnlUUTDQ/n/wbwTrKy7VIOLF801IBEfdw+RY9LUhoBzqaKMl
EwphM2w9da9M3qhTNu7eNFIPg7VWcRLUw2GqRw4N2IHSF8Pf1V6mwNmx4oXNj3o4CsMEEXDixjpH
kxJEsOJQMbFR/Qvd+NfPuwyivaDZ5X9KZW3x29M5SAWOg05D+4Gvz6eKN1n7yObOkdi352PlKy4x
W+pthzJfhWtjdzowNTwGv593rdrmnJuCDDUUgC7Gm8uy6cilMf6w+hxqcNzjhplnQPFg0mIQPta9
3KC5mMCWw0aLGI/j49cRho6yV9OlSN5RW4NXtOdtFlR/3bLxOFfnBYPparR3nUOht6GE6NHfwkdH
ZBM4Q59lVigWfU4ZT0EKitT+lue+RU6q2+Nqgr5OkJFCAlfCSXX5lrWZp+Zaq14nVhIxzrdzixL7
962Z0+WqDMdw0JcsbiO1r9QqGMoQ7WuGYIKN4N5Ze+m3hQ+DuPx/N0FU78wNIVZsNQ+Hh9j9BRyY
4NTzQ5bna7n2hVa8cqw0uL/iMZoJn58IXSQIIpnH+X0CkuXJyKEiTCM8wNErIpvheS7fdJYr2csM
+FnbrSOl1wlvT2BTGJ1q5Wo/jU+cqy/D5+njLexrgxU9B8znlJQN0/E/GlkdNK+7DlRye8DKbHNb
XXwoW5/Lv5ZfR3wvqMfk/GHzGEXteWz4yFw4aXLICs7PWd6725wpVo7ZfH1uERRjlaxBqzRT9mBH
uAu5CTgzl+UUm3bErtsBkS53d4FXLvvCznR9+lo34vXV2FQuunsh+Y03iuG/1kuBc6Y+ZffSr+tg
mCOTnyG1J4hSadqtGh3rVq9tTvx4Slk6V/to58GCFRiSQ4RvjhjzSV5jmYoOuYgDBpCKMdaxvWat
UNkpGcn3ReLcARiohBv7+fQPFguA9vv9xAWAMnjhZLCUEYo0SmdkGzj1ggF1GLyqNh4kiGfddgSS
LBOZ3FBtrMLHO0xE5pQGYLwlAhuRNRpov624TDh6NZko1xCGsj6k1hS29J6Iy1EL+1Bwxhf1ym7j
yh49XZH2l3KlVfKcmkNDE/ioLS4syAbJ4vjZj+S2k7CjoBtpUr2cs7Fp9vT+WPVbbCDnrxztV7XT
blYB/L/uWjeDWZqBqk+rgVx2s8EnOYn1IukhzcHY//UKd3VdXtfIwd2BmxQIHEhDr+YGyTMsFaSE
WcZUl+JZUnmDJMjS5pzRNem2qs8eDZbYgN/TVdd3vuypR2RMo803qbT+wWZHdFnnDvkdcKUFKhCi
QQyD3/cF6PMJWiOSF/9YDsjvyeUmo2jrN4Y+a+uVyxKYtQA/29HHH0YhdpzVRA4YvhrBFGmkvz63
J+W4yU1qDRsP+ZA5cplIHFUQTaNLIeHeR1/WC3JGYurHipAIygxYFdZ2DwZ50nYqTduEGl90hSJT
td+d6H3a1WKZOzDAlDFCElVHh3yUudDLURvwaCL/KjzR6XBBDMZDpKPYlbFF++UbgZWoYROv1G61
3F3s2n5GpVlTS3VvZ5PcbhH74DkKMXbTY5mSrDTrg5wYdovJhGDhTyogiizDbCyC51OVqoHxPDXW
NsNi4h5f3ca1YjvF1u7VhB/az9dmrFZJDoSNHeQ+e/uZVWwFJ0NTJH9tgt2Orqg2L+LVP+4tLOoq
39S9tM+KvdWHEg7+QwO1keZbdtzuFEKWfPtQMbz9YFU4w9R6e8G8hoc94XwqOErRkmWkPRU7ZtXT
crE5HfWhYMD2ucZXbsIJIkztAplkRguHVq50URZeqr4Y1Ar1zdBv5qssIoU0XJvsbGKCbc9n4T7v
uRA+fKwU18gKfmxD4meK2Q03f9DA0NR7zQtyvlgF7W7z8Pu/nx9/XbV+41qlAeyIpC0Yyu0MlHeU
t5ku/fftUIgXZoyFxSZV3xK6oCfVnZ6DyXWqOFWKrMSr0zAPWOpx/4lSqAa6whuzkdBDKAUVhWky
mVCkCMSH5/M6F84rhg4BBcrh3wv/Gy/UUBx0M5//vqEkm47ZvbW8ay/TjGWt/xwVo+bqL3x+uUXB
uwcHVTFa5+yhlHauN3BDhnFPKkh0iyjYarEK0ibCXNkPsW7BdrzHL92TrTKM42XWBZO0+buFrdMY
t1VNLI3vgOviI83yK+jj3xxezA2s7F89aXaoLCrCFvWJ8AiJ30JL4vD6FyIHNCkfLaWNvG/64i4V
9Dj5rad3Kka4Q4ITK43k+2pfYqX5TiKIoHUaui+YJtaNPAe4WIeYtzNSjZc+7L3LTAIIw/UV8diC
nGVPH67xzOybYhhyRhRAuxvmQxrJehoO4weCdxdWYHY4TBl52AjAeJ1iMWO42Nk3UNj/qyq1Gmli
FHpEqxkpQycl7juCQCBBGs7KR11SundW2WWvKjqePRaQPAhBG8l3f5PUqX3gYy8qhZDR0JvsGamn
iq5S562Kb3eyqsZS+6tAqtwY61tstCZahr7FvNYErUJqUfZx1zpGP4SB4ANfl/IeT4QM6bJDkKY+
6gPdNz96dOpaSkBoZ5uVJDr56MF0/RljrHwDW7vQeLKCXDT1aBz3q0NQRr6A4k6i9Y+fyQeuQgLz
nYZnV+oWJgjRkOm0LKLs7L9iWX8GKH5hf0y0Q2vSMS6QmXusjvj3Tw3mMoIP44vJN7u6aRw04JTk
6pZyyzw57OdO2iPoLn0xND+MLaJIEpc5EyiiTAyh5pjqpkI7UuHhy4mpl8acwAw6jK3M7K+jJX52
Z0vAKDVk8r/YMjTt74N+Ec0aentJ7W804DvMboDySILsKVZ9rL5chzeiJovJKAueC0wBGTyh0+9E
J17uQIPBQY43/jt+z7zzDKj0dKfGIKSsVu/DwCALUie+T2Ry+2YUgBZIVXbg/zvfZFi/u6HnSVlD
hpCv2cBQsinYTD2ji19BI/AY9QTdbeIUTceacTXDt/gkgrazHKUDOkLbMrBxUz5sgygcT5h196sa
5rRYzhAjlHKrScdPnJYGZtsV+6RfZtPZBbgifaHXfYYsRRUAGbqL5ZeDLzRXaW6+RBnp4YwKudmn
/2QCANcnguAZgw2hgp1CG9E2ITtfTaqFMjbqMT9lGSr7NldV8mnkMdpZvNDaa94yQ/LeO1A631Nz
0wmZ3so2MdpcW+9MuSO/1Bk9Cz6dNSp9eCb0CyAPAQMoJetJOKoCCZ0UZBfQOWuFILkQy3C4HasA
Z0mAnZx4+Pe9laM1vRh5ZX2RY9Yk3pJIJo4spbeW+0eoOeXEVgenceeqAMkDG1ZJjqf3hEDLvpNy
lRv5lWV74YkFgXnDhuuB+fKHtl5aN8gtwEYxTcvp9lGNGYsXRThA21tXSmZKcDu8gEPl8cSJXnzZ
bUAo3V3xvctaCpF8WrabfseFpX8iORks2y55bbLwm+CnNidp5k+k2d5pbiBTJ44/PqIGbeGhSivg
T5BVCAkMeo20kYrGRB2V86frZS/6E9wyio/AfDNpvW4cAWn8TJU9gdzmOxdwYu1is3zu1uvVYzTr
+v3lg660L+KoEhYcKjFGeoUETTXoS0AxgXx/atixtVuR/ApHDeXAUe73kAsR5tJvy69RpgCX9iPX
OEIzN0sM6guK68eOpBHQ1C/kAOWFobhq5tb3rBgX0gMs+xx8w/zQ0ICGKGniN+3Fm60AWxJ1k2Hn
j0DgyWtyQgpBNcq85oJTFBfYBkcYHNHaBtyJFd8v8mFNzodwdVQbr25Smf9MFeyo6lDu8FcH5UbP
NFq4jaEJby34GueNBCj0VTJEtN5o80Y2dfFW5e7+UI8q+yinSA2Q8UUPyCv0sBE2kJwovjIzj25d
J4mkBCqZ2YZLrRWQ9AmEfsXcOLCMhZivXxL0fkLtTz5AMzROS0tRChTzbXg3om1Cq50ZV/lJeGXy
DOXN9cJj3uNFJnsLGWSNbWqjIBV0LAPLEYFTxG6LeaZ58LCW4de6n95wWPf0jjyOYC2tNhmMZmoG
+c/91BSeaOYqSXyJDQDexJ4QaffsHdvqzz/fVNfDW/bIs9l4OCrkcQuwLDLp/BXLxla9AnQmNVU6
sBr7IVeZ+6Ql8Jk1ruoIKqr6rbyc8ukkxeJt6DPD6oS0fEcQNfO0Bw5wDQY5UnP849tgXTKOQNsi
SAc5G9Zh3s2w6OXM3UJMAtyI/8RGqkzq696ROpJ97nLGRG5OacEWHHBcexxXxuggG4gIscuhYuRX
ksv5vp/bt8NgFKyjHJ8WONdE9dpJlH1EGSJ44K18tAfi4LrJMbTELIGjUrCBJcibvIwSrsKxCipf
HcZGNLvqMDcdBXTS1foB2tjzDR66lc7SQFvZZdCFP74Xes9OeXccmPkTvMzTG2xzcU4R4I7HvcZz
YhKN0QyxQgp0qlKBzSO9+e1+0ygsIEpz3MwoSOKfj3quLnT8gt3uTJderOABHT55aLbiv/s6SkHV
fAa++79Z+Sn+XJI//9rjjL5MMy7Xxoy/kZt1hJ75CSsbFNr4kqePuH2/SNhdSvIGQgweWsksMexU
O/6X/Jo123rarwOXSgmG1TgVOJPRMXKPVDmOtPxSURiILs9QbB7c6iStD4dRPk32xNYZcK+OSBYH
gu5taZZhvixZx9ernoEMSw/TV9uLcT9KyeVyTI0/J9qpwH8lOaAebNJWIZZziMoUoj8uiarsg5pu
ITdi22QAvO7LWEATJzJ2Rz8nVO6weqcylj6klhxbTLMnknR1/x72aMSAnCEDgQ/lpzE8xIeDBf92
i0SXrpm177elWSllocXgONRcFB+wyreuio06yzqlI1nmLU55YcGPpCHt5jU9GPIe1bjlYWq7EGsa
nnyxu2DxJLMhkbGwr1ucBCHHHs3r0JQpZZEn5pMDLqbT7Ez2Oqgv5SKstwujLmwkZQ3xOJA69Jjf
kClFAxUzVPRRDnCVV+zfupzgtwgRCw8MAIUOOj3CQGKdkZgc9NRAJEQE2wWVfQgV7z5plAmF17hV
2A3k0vpq+f/vwN5R1bA5VOx1hQz6UoVKYbjkaWvAPpgSG41AkYjJNScjks2668PPUHNly7+49Die
7mUGZ8cJ661c6Ll0ENMWHsB7S3/OGibE8jXfauQKA9y4bNlfn8qBhwwXvzZttSIBX+uoTqt8bQYb
DgRBa+VPYMP/UGvBbabO1O9CGRGcwDcPn7ZOiMxu+nNxJfc86dLRhIcrjedPdIdRdHw3LTWP+b8t
YQUIDgXUnUQcgmXXPK2ELDjU9WFO2Cwa2HWAp7EwoN28fEFqiUxNsVDnnQBeJr1Tz/MlGjhclngx
HKqqsTSCc530e5JvvUl6qHD9fQd127i2gHy5FVQjQnhmOpq7uefQtJ8cuDBZlOcnqh+K3iEb6sMp
jYEqpf0ktVzfR2oYfHmfgt0xR/2ZPev10M6+2pNwA8k9yBjZY4todDBew6z8QoaFkLAseFsOro44
jEDIN2KZbzFvNbc3p6gStNZemwgTVUQ+2tDrGHwi3iZmbt/L1mOmC/EqGYDA8iFwM6AC34Vbw/NV
KeYXuXIbd7BBKwsm0TPlAfSZxGPkGSxC6UbyRh/cfiu0qxZFeEkkKNpSm8hF07j0m3I9hjVFrvwW
SNAfNQA+BilnX1QENw/qhpr1HTTIF00L/+NvYrkeqN9pxGRK1XwG7lpEyBrAKtDyoBpJUOE8zQoy
Ys5Q2yagALr8kSvUzaaMEiaAH1Ef7dKVHB4dAfqMJmm4rzDbIc012fiqGYXssuVQsimPLYfntPL4
9JN7GUH7jJtuXg0fomZ/yAY2T2X+z0Cum+XVfLigCJoKuXA8xDDoJeH7DwDVYtnIy+R9ZtK+rDpK
yERmmZgDMOipS+BZQex1Ynu2RAW7g3JrBp5aTNjW6tSTeHJFlfjjqj15SRJETIjoSqVsTbNtg17i
vEZAO68ZW9LMs6GZvqFkdmboPNkG7dDbeQc4jv2mQclHCPJ6ckQ6UyxnI6yfWIbBbejwcnfqjx5u
Pl8KIoPw/OBtlMMeLbgek9vXQ1lgljR2Df6B6swkCuVswxFWLBZ8vEBKC3a0mwUVXCBp9btQyc0p
yiU7dl4IGdTJQy/OHsOewJrxi4PjU7mulWnnLt4PisiJ7wRV8nTO9GORag7o3kNg1mXc5ZXPK+rG
0wnnKQLNEyRGSoS1Yq0ebsoI1O4YhQqcG5shBstV9jaLL2ZhwI70k9ojntQM4PeimV2/LNLarQYS
p1nO1yoUI8ngJUGzsAo2dhYZJxobM5OKn15VCOe2+vxAM14VfiVFqVp7Y09is+4/Ue5g68X/q9kZ
f+gsW0JcHvmVzk5vs0orOLCtDfszLnYAgRfZkKvAwwBqns0mKCbNsVCOyYV0VhZUTrIoXsubvnrK
GKRB75DtKzh/4qPcQXBb/On5TBamougQwKq/XnEsUgGwOuyickAh9Dwi8BzoL5UL4FlGrqvaBeTl
s9qvKsq78qyqpc+vQUYZI3izO3efdeQgrOK0lEE9YodTG9SeMeWOYekvECaNknpSazMDWsnKlGJA
i9AHuWJPbwz9C88TkJe1JDJOCQAUXQ790d/qEoaASRPhXIkG0hWRxiM/GJrxJwaHs0zsXfzC+wCs
KOfSNQcwaSNc3Q6lnj87xuRrgMBz1xr8+HVpAQ6PxiXPjcEw+x1DhhsCyVsJNweRszBDiKxFOyjG
7BkiTlFtlf3uDsMGdPRgr6gO0VTQGGztbJKWzYCBPpZbZWALYbHD+2mDsSAbyDe8iN59SJJnXnFY
1nYMC6y2bTJYj+ein8KlVuvOws7qxjuQwkfnft5gx7DVnSpIFS+CpdJKaFcnSLGUX2xfbFHpGKjV
H5LvzB44nT41pr4HJOlFtJBtpvI/AUzMb8T1+u+2sR19sUzh0EL21LiQ3//P4u0/bpjSxHEStCSF
7xxf/dzcVCDpAsGmTi2Gbw0+WWrq0LZBS4AWI+IRo6TkGvTABeTDpuM/6XhGrIrULQgLlUCeFq2K
/+X63y9Y0T3vYdJ8d2lu1iyRojCxQGAJ8O0AVnGft8UDJjX1L4jE/REiEANIHNEHx1HzjNzicCMt
2tztzemeLEkCKZHhx01KPzTuXaB6GIrFCpcG3c8Giz8imqBGDofMQgMTUvYqELp5oDYLsX/7TOnQ
IGLMRL2LKsHMbfKRqfssBYzio+oSocdBlAI13pyUrk8GBjdbikckUPgcKxD98FyUHD1YlchuoodU
9IGEQhfdL1Xvx3Jr00EfJUFBtIS5c6zh5ZP8Ia7hHrXetMEycyg+IhG0xcwp+aCY0ya4A52EKTGe
yQ9XuQG0LADR9zG4SeYXH/pejopRFZzvo81elLn98XqvR9jxDrV7acOq9NibNOqKYTDf+4nUZ8xE
KXI6OWS3prwqdX8oIi3OVsTXlN011+/M24IJ0xR20Gmfd+dTytp79aC+N5YFlwtansx2mY9fQqhH
QokH5SUJno6ww+NZNRJJKCl9o59Mx6L33JRWDQd3KDpLKoXGg6RoaUoOusJuF1zWfrgfYlMpml+L
SnbGcEs7YBv/UOrmuWHA2fFPvJtpu1qlmjhCsdK7S9/efScVJlNPtrPbHivUai3xl+MgjVQliJwl
fmN7B8FnVgw4FpgGMyjr0ZNWHdzwd9/42KhCB2BHk4MMqoreiZqJO3cyc89qX+lkrrp/gIkt0eko
/9u5nTtFWxJxMXvaf+tlg5Er6WLiGeHUHmtU2WUS8IkuPwkXPY2fRdSkVuXOnPedHeUsvMrRFqpI
cWUKIn3AuuQQ2Cm1B2i7v3OzTA8TetXWxId46ng2HzMea5/TpGS4QqP47dJC9HdHnd18cO7GI6Je
BmoU105aDlDFqYyR5xWOsHxMxJg8hMmrNlbMoueHYNCWdiNXJquanonR9RgQpYlZJDGqCcLyCDe9
c5cmvN9xzMjbexkzWXWOLjneamPVkRG5b8X49uaYkP10THsseS8oYCzYdpfFBvlgmwmIW5SVPRWK
fto7tMjgtd5pOPFjEQVApA57B4KE/vFd9HTd8jXnKny+13+c1zc5WDgJe91uUG/nvA2PZbwOYyg+
xODwC7cCtem/sl80ssqpI7BsTnN04NfyMa9tmQqNE5Ne/zNbPr6FPV7Mvb/9zIiPIdx3beYrz7DZ
YPkCytVQW42a53rouZBfwNymYAW9bvVe6z9eQurvYnWE52z+7lzffTmM0XJUo5Mbl17719i0kXhQ
9DYy70LstRglAY2XUVUqngJiGR2eKTd3T+p6FHW2BqYYe0kIL/80to7bZstfXsZ25Vtzo4/pN+7e
OXbmgNtkVkEBHCf0BemxAnzAqgGLbFQjGjI3ul9R98wQi/0LOZDyyH4Cpf4xgUh4LujzsCjpiyGC
Jkc72EZnvRjIDOL+tsB06oCzyGHUc1RJIQ9FtKbngRTwkx43RfGl0rqykCz09pJ3ZIZHCYovO7bJ
/BaY/821owolIcViJaT8JwRVu2tCedHtTkrO2mxxdyPXCnRFqDEEHKGeEpyijW5Cr9X7YMXbyMu2
CZ4xxZW01PYrQ3UGZAXTN75mH4C3y44mNpcOraQMSJWEjuu7RhD4sxd+jrEMgHm/dxlTmJYZJ6r9
uUOIc3yqEk99ocI+mz1/qAKHqjfVVAHPqJvUAAD7agaDpPqCnybrpDfghlgFgkGH+Eudj2Qro4/v
IeVYRTQFu2tChxhU+Rr99n05lFEzIkMuNc/BZxM4SM2uEe26xqny7TctTlMHBWyeaf8ikfB3X8pZ
CqTBmaNcbHek7yrHvZkM9AmYKAZqZIN14bSa6fu2YJTjJ6bhTBAGdoktDB8dE4yh+JYUK+bib/KK
Y3yDJFkF1o1MzaeA4yuGn3sZgNBpxTCNfN9dtoOHRUYfeu9n7qrciIPm9fkY+SZEyXmEkKotTiPz
5J1LUDBu9TlzNOa8tC1dJedogBlYKgcAJKxZYGZE/HLaNiSULVDBJiGdqCN2ybUqw206ZhrdiVR/
Jhp0hPOZwfH2FNuXAA0hXS49XsJkGqhOS9aMoe4kiBZRYYpmlbeqrktQal3m8g8IzL4/xnDQzMqT
Y7b1Lr0B6YjGDEWjcMRDrwcmk0sn1enzXtFA2jD9nDEFBeOgRfhL9G6MFNnidSjNMPNtZX/x8C2Y
H/c05XANJZVn3aDxhz9IwcbEZRP75VWU1z91MLosK9zF78npSLU3M8fOa07mLqOFv2wVkLlKRXM4
lbGgYDtG8Q7EHunopoMpR1wJ0IID48O54F/6UhVeZwFgyY0vJs/iIBssfzBCYxh9iQpLL7WnMmrn
9u6RCr5MiVBFi/Z1BDJZqxCrBrhJYUfz5hkCK+ClEpsWdCt7gUutr7EQXj5xd0iHf/+iv4XToIlC
pK5AdxZunYclfDtnOso6VOctde2oggCn518IKbRtJnlzMMkxNOoIRHfLFWN04++lwZGDy1V6YXkl
PaxLCCTMjJ3153SsaGBjHchkUppm7seTp7QJ6iRCTcz3dJyCUL1BjgNJ/DU3zwLNwUx8NT2jjBtz
yKwMq13Q3LigpJBb3DkZbAEJ+ott8gRZoQI3icTwd0Wwqw8M8kw9lk4l0BrJIJuxGT9U3ts/LMSy
1Rh54HzgZd9pYEPL3P+SYA28zaL9SZY45aLPuhSMdVAku7N2cZZDDD/ZX3w9FRQaAbSmOpyMVI2l
kapgas+HUylfI3LOztnJETtS21U8xMVPKBzVOlVmXwIfUzdqczqEvE2hh4JrvNmAVQEmN1tbxrtg
/14lLktAt3Hllsb80nhDB0x7a8v8zfEgPfU7y2yt5XOF8zQjtrksAGYEgFmQF4wovmu7EP8pAuBq
cD2kznK3hAhlthdzYJX2NOQpjnJg5rLLatUu0E16W7bP9jo9j6azHTifYMyYENBbj6ci5kaJaogz
Usp89+W+5/6g15zVWP8bgttPZ0rHpqgIjTjrfk0Wg9g0MQfHc8S2PykGRvr0fnHHYbhxWrxifD2i
jGwiPfOMxR8lJZY0fiSzNFXtzqz/cUyts/v6yYsBJZCcsqtRu4SwhKLBtnsQnMXmAgwCzQzBS9Q2
O00MSFaBtmDm23tRC+35884xI5lJlubEuQdN41QFIDaODBLNb5Gbi+cvBe2clZrQb192GRvP+lmz
27EblPVKvN92AcOEBfsSD4bW1+MaDJLgCx+kcG4SzxEIkqrSULtFYfUqEYSMLN/tdqi5WJvruVG5
monC6vaytDhUA/MtT2DRt0vO84eaN3aw4zcsiJknvj8MZSzPn2Kbytjs9tAlzW5YFHYzdUh0AZPp
ldOYJDPPqtCnx8705tKi5EYiu2qDkioMF7FWKFwOKjGYqHWVYrUCqAXAHD0Vdy8F8kcoRStarzFI
+wNq1k/6y2LjkCLvUXZYrE/lngtuhbz/fyxekqw/50FMP7tjUhGxrPZHCwaFkrCoJMbaYjKQFvM1
Bo7ZKfHYbXT5sZ9sqf6PgcFcExV4f5QAyJ95YfBTQqXbz6WO81gqnQHf+rAT0RSyeBVW/OT+FWxx
x3O1B9tq/hno5zgIKmIClLvzGmXFaCIj1ciS/Pevso7SJ4C7kVwV4RT2zbIXX3oohDd23KXO3Dcg
twDvraNPgdEA+C2HtSfU/FB6I8vPNNzXvLoMMtlK9nWZp76IZOz88YTgHuQrPMs1x7JaTu5wOhYR
xHt6It/wpwKLI+62RSBn3Dbvsh2HKMQjPCf3XENIhbZ6gYA0TpXl+kS+Q16pOg1T3pjRu/H7eFEn
dIce8xPF3Jc02OZI0jOMEe33HJI8ppCaNgUEHK3kd3wt4vlzE0qTz794/UnJivwPjk2M2NMu6k/y
IXZr1cj4DCvSPmXMMH8YxX1SjoaOHQ6My8BIB+/wjh/wWIK5Fa2S0oT8z0ozhZlj2ST4ilpUA95T
1sdkNDOOsXtpNUPlhfWeEV9heBHw8vkuC1Vd/CIqnWhGwgG6ypUE/n1+vThuN3Bxpj1URN4+FJ70
zh+I0VvMHIlDgzYBtkWP7L4us0XubO+s/IFcvwwp6YEwC7AoSV6yaBgo2laG+YG6MCQXK4gb2eKo
fmXb3d+fwR/JUX/rLDXmfz1nXNZARlcYLt1Z9uUC3ov/R+MlMtntgFKvmsC1ZttXRJtrT59wOoCU
1HdTPsRl8ms1kgpUMaI88UPyNbpJuIIw3v5RGSxcH0vKAXkXcPkOa2/pK3QM27cmR6BvushyquAa
vCwdIh/axSxoFow7iz7/nOAV1/zbl+TaRPfSmVUZFeemsURkdZ5pumLkymt8I9U0LYwbH8DaRttM
2RCS5J29FrvZSMtJGrPilgJRYQRXZd8gh+ep59LOUWlW0sbjZ8GDhT+tLUCSShYgR9BDcuWPKchJ
+c9PMN+dkxPCDbZ8SsmCJI/p1/VztmqVbJMolmGQxtCg9hbWfodp13yIrvJhlKB+wR7v5eBSuc5Q
D2W8+UEMcWK/J1dvkaTidpPlP27bC43lyxcAqYCu3W4wwMI4V4ZtREg2ryL4Ve8GOTgFdwAI5fPV
5pF95ejMb93rpaXPEpJXtCAyCEViOYylo4+u0ljirEBB/aeaDhlFiQXOD1KQFcs9kNJDYkwcANhE
kf1ymLMZdAt/73T5JFzO7Atn7YmqlbZoG9R7mA1N2O0sJNjR3UopFcIBmKrT3dIfQQg/NMAmNuFJ
+SAhcU2dM3az738OtfMgrSUkeUTaY/iakHZPYRWOCFLP0fe6lr802ibxcNlYE33jTRvo+UiGqrCz
efOGNeEP3JziQiu1d4JNL8WIwxncNCfr8m74FY/zxngQIzjoBiKuYHkegoe/4He6v8FdIYAf2fff
s+p3Dr6sY6wbAkA3CmJZLsa5Kl2NaFBkk+J/R4aiYwILAbT6/ndOsrSYKuCNMxkAOUo+4gI9Aq6N
KgUpExi54i3dJtjabMwThWm98DWCICCRDiA0HxNtViEFLoJRmHLYHQ+wzcQHMk7PW4inP11+x+IN
4sCC82ror6+C2OUjwq+cU5rcRLVO42DIyrSY9LKiQYCMrD2SFULAdJ40WEIBUj9klL75sl848/H8
lRc+IwnVQA8owPu8i4s1zGhjOBRGO3sgI7W+rnFaAWCZqK/3a2Qe8tYt1WHcIyamHvwdLN3oXTjc
PU2P4WpeBKJp3gm/hBDj3/YxRQ/Tcb0EZ+4oqO4O+n9BjiPWozgJriTReXlCEQjXOnk1ycUUJZiF
+TQTWpOOFiEDIrOIVeUECQ09uxztGkD2q0MMuh+PIiyeuPydUm+l9Wr5y07CfD9Dl42ko2JyVR8o
cnIHKKsOEdLwKxPBpTFD6Ls+/peq8o5PbIFABCuX2Rb4Tykv3ypmb6+RY7DB4Gsb04pbONlOMp1g
sCwPKqneGPGBN+KOGX0PSwc63BWpBsFDPV/7zmxNkPEE1bTauREoRgHNO5R6V9RUj036pGX14PBu
sNbsicWjVPqFGdqcbtZvlJ37rGzv/khQvEqbBxc4rBBHVXODa5nMqok9v2p+d45+XBvSD9wxCCy3
FQiJluQhleZz8nRWIiXY++qI6xuTpqArLvMD6BFA5M4zUlUYBhS/OlcXA/h+/dCsjjnAR2a0UF7S
Mr7OlAD3A8+ZAOJBbJS0pCdMPv0a+LGSIxBwvpJG/wtLf0Gx94hHuAm2h6Ruh2rHuZ926PpacKni
1mMFNJRxZmUaQl9N5CK0oSc7rbJS7qrfQSbascVo23x5s5ZtPnhyx5bXBsM0TTiP5Y3jn+go6NQ3
lWuquxSjzT/lDsqAXfEE0JjON0DSObos+1ezNKvlPGHv36XcD6fnMcldt31nGd1MIwZ2QLQyylPz
FpeH6z5rLso196egIwDwdAegD8l8P+ZkHnz0C53YCWhkToDfMY5CvglY7pQYlQ+VdJNGRy77B8f8
CYqw6OWcysiHl1Ve3gp0kH58+/5dfN/sU4C1LlH1rbE2gE7mXoaeWjSZM48CORzfptz1CBPfOiQo
1MyPEWltMCBsU5fGEyHE2RkK0aMthXDTgKehe+QEIvAJAdYyDkmeG6WLrz0YZRJOZbm/ote6oRRQ
nBMhoBIWXO14Ducq2MHzeoLbAknLsOkIlXOrsmWB8zJn9pWpoXqDe/lJdOr/m+tABbxNaOJIbqqZ
r5Q6sJlkT3mhybRoF4yGkTUppuUbTIGJq2OZyrabwAIHlSRKrtI796gI/qPZXUOycrfMTc1GDMoH
yRMrLLKkP1muSTvTQKaDPjNkfJSg0A6+pqz+6kQnZaaHat05A5tRLObtGKTHuJq6AjMS/du+6Xnp
AkFO0s5GY5x/3NeZFbHHpHvdYCOmaEZjOJHK4SPgRX98oc0EZQrEXq5VKnhqxIBlPy89eXxEP0YR
0VaX5zFCf0QdtjbrYbfAchVNhKNZqOLpG33nzFsefWV+mUP23H8ph9ut3HsZ19HGEP/g3hAZFt2o
l5ddI+T75c3eogZZiAx4B1o9v6DzWm1Sk2L7kQGdfAVnd+VEZPlm9mnmAxLxN4DimAUWMQRBkJWR
mmZ1Yv4Fd8skrieiD1rgVML0E/QnMySJvusMLlaCHkKRna2vnbPRTsGvqS24RZc4J96sEj+jGfwn
vxxDCf0FwRpVzm0b5Dpu0c9W9dI62nHG+A3kdhf5kS/rnyXf1Q81+R0D3IkDJu5F+TzlZLVv777k
+xYzBo8Z/90pLlbE8G4pjrGK2hcb2GF3FyYMoE7+HTljkYkx+YMGwaSyTNmr7zKEjFsiYQGZQB11
eGI/NHw+QGt2aHJMDni80+YTjHj4k4stByC+fUIYCFToTZiK+DIigOEO8uyLuZRo4mxwvkK1Lge1
kchRo6xoTqOqoqhQQieDO4sqUb6zVsfSQe9c0YTSlFrKv0iRAhgCP7Orp6sdhuj1HJ5JxpQ5FDNd
xvpUUI70HS4momPfPQNFHjHwUC+MuPkrdeQIZ/hPPKR8jSb12DcWU/3NO2fhlaob3iIKUxA1LDVw
5CEwdBTiO4eWB4ZRkt3Almj4uPEB6BUI2zfzr+t70WgYxMfWBE7gepOg0pJWuWy8+2Mxq/QZAO3y
JfwJIUDcy9ftyYhprIYz1CLAJUtFjCJY9chuJU1G/WWxHpQ5dG8fh9wZC+N0Z2EkdTTTnMj5q8MY
u9bAEaB3M0u+S9L7MCf+d7Vcb9N3Zs/fi3gNcJCdOBZc/g3sJ32jgDlJiuOIpP45ZeKLBIkzwCg+
SgeT/eahFsuQb0/hT9cJZF6Vgpg8vLIiF8yNaxzRzlYI8tbnme6+J/3S8K4KQmu5GkmouUo1daZY
IVwXNK3U1lh6RrxkjynHMqDl2ehadwuBDOdaBQ4PzTZo5gu6JunZyzfu9m194Dp9qp2EK11XJf3u
uBZ/xAE97Ml5PvyzR3eR4IqQuDLEYNoPBlgxCQcVg+F7EiVfwSeld5ZsYCUSoWfkZz8Zp5wKtUEg
A3SXFCLMlWWsBbvKCZO73ScsKaUu0CcB98zyWSEhA1Jzn0boFmCyQm0sm5RyXTKPZ/eevD8WP8Pu
FO60gRp2x0ezwiGRooKeCNfqEVxXEWk++49qUPIo1pKAPqL2w+X2krnwNRLrE91CtsP9jRm04oBR
BxUXb4guWkZh800EB+Yjp1hY3Nz1oNXv/sN0vfFQzkFjT64BhF4pDV3TegmgDGtlgzrlDgcsQEoo
4y6osfs0QAgQD4M0qr6v/B3eLpMkSCGbCTkTy+hQd5KEUFR8UFdodCe6AhaAfkIiQNFfu9AfxOnw
dh/5MItPdHVn6UZzjrQRuDnNSdhKJlAlqW2tFIsitJG1DCkzoh0NGnqJo+kwMV6JTqLoJUlSI4a7
zTwtcHq89dxJH0tk0reyjclPEEppFvT+5x6/stXDLIpvuONlbfWRPCrR8rw00M/fq7zUl6AZCUYK
vBuKz2o1fcCRvXOyCrCc4ld7XYynVSdRTP5J+LE8ngHvwEUGbLKjnNwOdhAAafAUybXa6hnsOal+
k6elAVcxJrJjkpB7dUptz82tk2UcG8nLvakuYyt/GKVWXbGFacCN3EM9CPA2QDjOPL90Nt6du+Bj
Tk6j+/lBqQvWg1xS8T3uKJhd8g8HeeYrexVrKqsKcEAl8eAPz9/keVxvL9KblhvXfzquj28eiVhQ
N+ItCoAsH2hwqVr5Ch/ns0X1lqskabsMhvRJKIyCIdDJBaMFGyhpKFCRRf3GHJVs27sygXMiJEB3
TkiDdBpjJfbo0JqSbMei5DeCwoxV5jsWWIpb57AaEZHLlPpeSh20fei2LowekjFNpIClxSVSXZkL
11Iuzau+aaQvtOVqz8kpnDM3Q1rAQ8bDdfCS1Rameyn4Vs5gEhCwGZZG8DErqXAQRGH9zbtFkRws
XUpvbNpazH9xMQeGSXliMdzYLlliG9gpO75n4f0cqMPhsb7FNgWQ2PEDN2QY0RePAMlYy7Dgeep6
iYxaJVrOxAm4lKHyPPHVNUvayVAxOzDGOy5Fg8SzJmd6lO+CpgnQKKcaNQaTdnrQD3XHejNcPbjW
SlT5YhGmr3pxymG6abshjCWdS0VcxYW8UN60PyAz8zoiZZeXX5xk3WlBpX3Unr4lTQk+8funNmsz
gR4hiKK8BBUexGV7z+jtvTBDTLmzTon2cEMJ73nQe6UVXEHA7FEMuaEU486KdtlWMhvSKVVLs04H
w33dnguf+b6Xmc607NcNKh3chiAwReOPUWwx8qSIT8O36DqprhWtuMOLjz6gd5TAp70ZR0Dbxu8T
moCnzgcFMyjONW6Iy1f/3fZzWPmpOSfXTKbLOx5bquoaDN+rltDC7PfMUkF7BZ14iBPG+1HGyHN6
dj5IscNgdBTtTeKhwN7lhpByWODAH4vwFg+2bAKxXK6pEatBbJuDebwWN9KzZGiHv2/IvizQ5kNe
sLwRm6dYqsMTg3txgwHJ9JdoVChcKedJw1rKqP+NmteGuYm74r99MCNZo6QTbmLGWHkYyNl2N2Vx
29X+SFRo+B7KpMI988PzGDvFyIQ/w+8IVEtpylS/2pbeTUFqNutNVdJ2h3CQtDMDWX8Day3DhDUE
eAnrWalE/M0Y5Ui+dok8Ct9eAbhJkVPBB60vTgWH2KpFWkwJsEm9oNFUJk5nL2HKFzmAOt7Jye6f
E/B/IYiMYrCEDMXIcR5BsB1Jk7FBr+pS6jZCQhi7Ghvs/++SBFJi/ahT/R5ww+Zd7svTPu9XWI5U
Fcw0/F5Sxo7sqFuX/jy3xpF02kIyTuV/j2yXSbNK0Hobgo1pphl5BvEnfbeaRA4SQx8UJBquGmDF
Nwsmbc4+7PZlDUVJkfGoXx8MdIr+lSzil9AJ2Phuy6suty39a5ji3LoUJoyOxnCdA26E2FUv81i6
4M02dexdXn0IElguE6nu/DQnqhYbyWZxYuzRTrCjAPeWpakxBhxuwoWGps9GIQO4U93aCoDxwckD
Rl8sLEBfs0P8ZweWEeuOuT2hENDAPGCocTlS94hqpvWVNiVL1dxerOFfuILDRq5S6XpaVn2Q/tCO
SSkN0bT/k3T9oa8XMf/Lhz0ZtRtPgUrrBdzoTRRSf7YVVWagvM7qvk2RBQISlRG4tXeE66zFCV3I
/9P5yLJDlOkqZfQ5UrepgC8mXdMUZNEbZPKJMz1/KfnxIgYoLOFlQEf7o0MDPjn5BFT/jNEGnuQq
zoCbC5iyfsRjsKz/paR7FTZNp7iLwyyNOiXipuufUrAqDoS1rFxBhMDFY+XOBu1cVPVOCQL0gRxt
moppwVFdTn74LjXC2cowUBGacNcTYDT7lO3aUzwhZYzHeZYxyAHgXM49gCuVi74WEQSgfaHo8SDr
6Lylanew1QQi+linoATfO1GFSqyZepZjjpj/7O+ho8sEJTeWn0Qe6UX2tlRbxIzGGASChCSofQI9
sx800Qs/5hdGEiK5xtQy1cPPknXLnrODg56olWGtqJjXvSKqAfdH8py11q6NchnDmGUkr0NTWNrn
39BdQ1sQboOW+drNII5aPWcd8ykEFCwIczcyT1uD8f4Gbn+QgpmT/qHu+MMFrqXw8/BWsYNAddHF
k4+6pUiWGMCQKY8K5VbFScGeM3aEJ+24PUWFKh1ed7lSLdKNCsbLlsUmM0/cXRZGXXvswtFP2Qq9
gLvmOWCIjNo63fDGjvt5N8vkNYbZcWOebQbh/QNgveXPKM+QuDEoUEwxkj617d1mnEOirQPevK+6
PvsLPz86mNqmP+nZzTbdH1AQNe+hki2iIDESGIxPSM6KqTXtiF5zfLXCvAbD4mgImPi3LswOWzZn
6nLRMx58HgtUVc16EfcednBx9K2Mc6HmcFFm52tF7bQqOGTmptww2jsGzoktOBv0k/02h3wQQVqM
vZZYxKy0Gyg+6fzyMdbPrXiN1vlCBrmzzjoRtkxahOfXYP3Nmm4bL5MMpJum+1eKBas5LqZerKol
fkGAPvDjYtjgDI1oJntWT9tMuTs5JC6k/n/awN3X9Sz4f93kGbaixDKazKlZA4X1cyCpOcEj2GyP
cLqYhmbjaFSvafojGEB/gdYqXSkELoSf3F2PTc5pw+JA01+3MnLV7xd87eNWJzTJdmQK3DGBj1gG
OI2rcX7Azmw7cZv85jKUnh2raIeGekM0SWsOl4+le0o5/iKtruKT+edsacqbl5f13CHE/abShv4R
qkBQRBfqZX9GzrNuR1IcZcaVPmNy+9YTxOjUWTI2mkva6dg///hM6fdy4tBOPuSuzL7H5y9mpYyq
tT3xE7oWHR7T8ea5b3vM/KEUNRmCWRSaQvyRDgVYXO+7BZ4i5ndj2yCZkmj1H7Un4vTyCC+CN0I4
CHUxCeVns5nyfbR+YsOiEWlj2N/PRd6tow7LzPFIogugvW9gM/kHIoZdA028qCxpj/WX+kZ8jq/c
u8WKC9aob1pHLRwxClDy8/ufIqItRAiRg+JY+VJ8Zx72M2ifYls84dgOIOkV9Rkv5OFOikoIZSn4
VJUguIJYbzpJHmR4QgwJO8zRFw/5GqqYsEqtP/Rk22FBIyeORgQCB5Tr6uGQ+vgoZ7KoTeGuwGtF
eF8zyswQd1mG70Je8bHduPoNs6vDlW4HlDcwcxAzA3JL87t1Vbl6idPCmrHC3sefnxknVh8mlqfA
1sejrXwCGfLYXVXAGVfG490akKVcYWIlWrQG91TLCCJfNUGKwEwVGHKoiSwe8ZVguSv5GhUI0kQ9
kYGaHmnn46aT89WH0/TaX8N3E+CKS65WagCfq55JIjJM5d60lv6uxRMFueT/fDuBnbWEsePwigc5
Oj2Jyr593870CFKt9u/FYrKIkAdpqplpRdhOg4r26XS2ccmc9jTiEPlw0QCQikKej7+vqVI2WMcF
m4DJCkiK9SZdTfrWGkye9+98h/eW2/vecwKm2tR/tX0g/DexHo4gDE50XFoZIYEDEJ56H9rvi7OY
YjEz+rMxQDGGDNMfJQ7OsrSS+Y7sY4zQjeaD86ry9Ssld+jWia+ejAD7s/gNx9Z2aKOpeCQDV49V
OYM9W/KtJbkX9Efsw4RM82F0lqnZyLIFaDKQ28eusCUTablzeEu52P+8jl7K1aG/b9s0g42IbLKe
YW5ywMiLEDhOLK6SUBNq3b80Z6i0wyH62wGWPpokRCqYcOaETGz6Kt5cuC8AKtesM/tYpA2rGPsy
49bA1cHRJ5kn1U/+mDBbWpyd2gPvaMcKGtOxJaaXT6FFAWR922RJW+AUq5K+AWWVICgXwth5qjto
wp8F0qN+XpvS3yDB00cWAIsLTltbehoASXNKn9L8tsuAeWdBo4+szsT67Yty7WNKlB4shg8ORJJm
OP7ctXefweDoePd/srhojcsmYjIxm4ZAYH/VwM1H5JdmY+g8eE4NVfGXtRS2BA7EcrjNzd/AOxhx
R9rhotKvOafuve/TIZlXatAK72onzwaNcJPQpcadoPnBX8rZR2z+4ZnS3Zpgv+ULEgleyIflHWvu
WW6Ms1RZxydV2FHUsObTKvxfZjJFj8T+AffwQyS41esf7+8+5cU/aHD2zVrglxaP4xdJpd9bGMa8
vw26dpwzb+5wLHOQbz7jlDqnW3xNdoApLOmAh6ApkOA9OAIghfWg/j34LyH80GKOudpgFh53XNgG
6W2ZIpedKkuQktzANw5fFYYHgiB7EuQoar0M5ETvwzs1OPou3o6SclRCQ2XFZHLOz51mCHe6dr1n
aENQkVnO/+Pa8P6ibJI9F77INGSe2HiEXph3T2HNWF9FplG2HhE998QPIm2qTtVcSBkyIB0Nq+7t
JXtQw+rveDPZEtC9oFyHGkvNZB0NbJ3Lw3h80u36Xwqtq1jxKlfgE949p5JfBR3jh0ClwwhJdOar
RLXnOcBRuu1VflWmP1EldpaBOpR0AobqRWxvSd2JwrLdvJBOetlnhoRahAzgBd8YmOVadzU+FiAo
LWYLm9PJk2qUIbddu3OJsRzOfGvGGEOGy5HjqX5uqJJVQJ5hlxZNVMWyZWKd6aVnzSmLMj5d1xoT
z3aZ7pap6Bn6Dt8FWQ812MdL2Qf5Z9BFjE6LPaVmLeiCkCthZGbcOmS7kExyqVeFNFVtOYmoE1Vu
T1gxe0n6w9zq362+Bn/OFlbqGbmvS8QQEC8YEnqA+gWLD8xr68YdLZUf41kzJkP0PpKhxiXpENPL
vQ+wjzJivD14EID3vf7q1eAYj/5tR4LHcwdhnEcwMlexaZE/kERpvDd+j0fAqP7p4x+mL3bEjeV7
xheHtE3F7k0SV8BC5UDHC+o/m/yQ1SWQkW04FPBVLMqAuzdzm4u7rgAUkJjlJuEhF2OWtybWOxSD
ko1UBr29VzT4hWKeAJzCp6X1XsR1RbttHbubK+X01sRHR5o9aCrkTr84Zghx8zX4G/ao/8j3igmV
WEXwKv9Sg5SHs4SAV30yUAnz9YqC3O+cMKjnIDZJ48KeEUvySt3SgRwCmwcKRLzlVcvNRMehS4eY
XvwjqxrSxgJYG4pnxhcwr8F/ztBjVsISE3eFO8UqDSYh/m0OpGMvwNC/2xdNJM11LFtHbUXSBSj7
nEm7xdw38kFo6in5Kdhq4xXaFv9aB26FicRyP0LF/Pc2/Y3chZH//jKp5iWmHfQ5kiY/9Na7NMd5
64POXynE6ytyhO/oh+a/yXoIZkM4xziqRxeqRkVEKW6fLZViUs1NyrAHiPli3fwY/FaOTPtAY7Aj
hB6fynPcgux0gSaMIXH4Qt5L3fUlhYc0DlqT/s85RUVmYwG4zL8JW+GXYSgF+AF10Yi2VS4MVn+A
UU6RqoeqwMsIS2uN/uAHqzmH3AlqMAy8Fkq1uxeM/WpGmxEOIAqbUzaUbVsKGVaiozWAdr6yjFGB
Kim9L3x0736GtCNHCcHZa78eSjTbVW9O+hJZ6YYlvJaTdEWuRGhz3OJX3Ux7eZQiqwpaZRNEvYPO
vumoabctPPzssWn39+S5Mge03Db0tIGa5O5YEu8x9FWjuNH/Wy0YRvE+VYDuKk1oFoN2PBWkLCvZ
RcC+xLNCT8YJC2yi/4eKlaNvEl42dR6nUe0xFif9lSwHv9iW9ZwKSvEplfTli5H75bs5a4rPRmuK
bnsfM4/GhhSmIX2UVW2ps6B6u0RLmUBT6cXpZBF3aASpAmoDCBwUOpP8U1MBNnNnRP+rjnhKixJA
Gy3LH5t1CIQRi2sXNMLwf2Jj9MS7vr8aLkzirY1xe+k+SJc9mqTnrp04EfyIBWx4F2wz+paYpoCs
pMz4LjBQDYDHjKKIHYD+LbAVlHlL6X4l50RcMX0+nl4xCvitpWj3mX/oHMFUSeUZKgH7QFZnQxIc
VQTeczUrIZIZZV7ApXBEXqJaWlS1tjdsPWJnj8kktJVEvDMeVCIXt4Sc3mTVbmdKWHlBgPkfEMjY
YtiYIkHRxDzsqVe8GApfCQKUEXKxgdU0lvwMPfTH6G9SB5gSQFSKjb6uHiK32meoVVN4q60TrDDR
BvupKKRrXXhDcckiNteCGMbw8tp7XXQWxwfW71aRF5jThJUeaPuf5tfJKHjH7puq0UjOqf2uUdPr
QM3m8LAQnDFghx0BY2KKX97vMAaqH1xAVd+UVCu4hQUgYQY9g0o7nxclbI078v95lmGCeQ4n3lu5
feFNb7DoLtUMw5809QpqaIyyfzNkZLxdDfX3n6skRou7DBxGYbyBikKzriefTTtXq9QHIRDI0Z0Y
xD2u1W9tt2hWbQ3tegOQjxAyE2AO5+2Y0IWcaB0F8NSyQF8nlm6mrov0jOErRH2gsnLOpZcNJm/i
W+aVyQfBub5/qr5j7q9rIQ1/t7u8y9qYu40HD5pSKom0VnGrOi4n9VN6FR5qjfubZK+JmwDv2BrS
6cMMaYMV9bYyyvrN0Oy15hjaP3Vnm7OaomLGrbWy51RZe7qvTGEAlob7mpDKxE9BHcC/8c3vyu8l
+oNj74hK6sBB2Bm7ueWTSJ+1mWZLW6Ht9OJ6DqMYfDKZHzc5/0do4pwkta6inhKwCtK8c3llPt9J
keOhxfGrQp4i0SmjmUYkRRwSGM5Dhf/bBZief73qZgSeCBIkocqYce2vmqiUFANq0xfz0bMWbb5k
VhgRVkTeDqmV9WD+jTZTmPZVw+15KVSNkhDAPBkCqxPgub8ssqqvg2qO2o1/aFZyjPHcVuShi4ia
gzVuZOMgI4kY0nkXskZhRBT9QCO1QWaMtRv8k4oLW0AuAPIiG8w7vYtsxtBfD2Bev1bUeGgBmZs6
AjtPy/RS2hni5k1mLFVuzc5Dy4C35rDpzGimP1P660B8V2Nw9k7c6+fW8e81//c2NHFBKigWO/EC
KWpX+honjKuX75WoIsn/eq1Dt0IsRjah9J2rSAWprs1YYIuCV12xy6A+fB+AoT5WCpL5ECA9RJi8
t/ClLU5HZpWppin2yfzLu5iI14lIOWamMiYoOQIop4F22qTB5spsQ7N0o4M1N1m2NuHleiVi/O2W
gxYt8o7yIKKC5Do2b9zgMm6hj+e1gKngBffAqYTampFrWIRfrI/iih39q7BDXOgGLhFSlLDJqgQJ
C09rC45OUYNKbWA8ZYDGowPnaOuVOSEw6uzma2sPN1FpZFYVk+yaddKvL4Vp5YTJs5uAFyL15ppx
/q8ijQjSFtT+22TbQb7LPNaRcyRqvbURmbusZsWQLVWsYBX0RGZ9nLjw9VWfL02nIYBvUbEs2jFJ
2Gi+YKN4dAYu7mBRvmVXk7ofD2ZGY9gSOfPJ2acszNR7Ckw8fv7yzp5EbDGAnl8zWb52lgTMV7ky
DGBhHI2gL+5fsStywVNxmb7kovtB2uLS/siBJeACcQ8SIBv2R5auRe1FdiKcT47OnGfMfNKr2hZT
ToTSF2mltHbjFzfpX2nMaKxlyXb7s9zxHlEJZdurb1Y8utMNHicYg7tkmhapbrcWghw17bmQ+M99
OGt2lsHvdUWGHUkDA6zLGprPLC3IX3UblHCfBDregtfiLEXLB7Aa5LvZPlxb9vAJtK7TgLtHbS8J
wocXNZouVY0OnGUnY3yT/UevUfsAZN5T1rQezWM4IHR4swBCNSjJYs95gOikwX37MlaqRQHcueSk
t1koEXsiIITmFJn+HXKL1SvAeoSnpMypXd670ikaWRGUu6xL5aS00F+ihfvv49y37WtQssH79zPi
tGEUapgJ91kN0Uz5pKQEX5Q6yS3V7e8pFk1KxQ8YksVsBI7CZHbDRpiLnqelgfzGrcw7+uUMG85W
KdulgxE/lal+GwaY0n35NY/gjwEoHEa2Ljbjz+aVoX5YIN6QMDA2btZojMORTkoqh6ukE5yMsXty
qBA+eys0dGj+37KjeJgyUwClJYCaG+Ke8leBOGU9IvvWK5HCSka4Wl8eOk294+DgzYOfPFx6srjH
5VxH508t89rQtm1WFD7COkL5jWL+2S3PHLsOPLnLb+HsCeHHLCpOTdcF0knbWF18K3qOfQtbvzIL
TCNNKisIWH+7bT5ijMxoULF8FDusn6bzo5Uivcejh0v28jQ1ZopUx8TYyrfalGBNb89E/Y+xssSI
F0K1zRoc5TXhn/5scP8L7j3CxQpAkA5zbj5hbBXJdmAdqZO/5lEaegi1AbpJeEIrI5Zgu0SjdZ/n
3EXF7FdDlEDHWRuJJv4MezaclsjELekMlmv501AajJklmUY73D7qkKmxE7dJ38bVktQ+qy+NWtCS
H8hl0ClMIFhplenZbJkGOJzxUGvm7LQYz9wIvESgb8P9fVHt5obwhmzRVQuzSaCxJIy5bDSFrHpP
Uj29LPdhys63EanFobQbnTz0diG2F93PDoo8oSAlgCK+tTXMhX5hkGahTYLuBdR0i5ttREtkBuTQ
DIRb50JPOW+CudmPwYFjFNot/HUrDV/Ob0kio5X0m+D5d2q1V/AWUpv6GRsFUjvXX1KJ87g3/U+I
ODJd9EqGriISgfsHR1Gp092hknrCWAc6TY8cVBZhihi5IkbooullouKheOyKN3Kei8dEV8FcTpp0
d5mtp7RrXM+GPVcPecD8E2h+GaKrNwhnQu8CKi22XVioVnPI0t7Bx/gjHs8A6V9pLCsGfsFEUlSt
kny/cpcm5z1eSHDNss04UhSHElmTepKm7W93rdoPHqBGAa4z3bAh0HGHiY3sQs5LbM0CAzB/AEey
C3xEgtJTRADArchOC4BPTQfcQIklzrQ5bakuV8Q+vgrWPssX+CEFbyqo48s6XleI3FD4QqppToi+
JNDqAAbkC8fXQznAppq6z7Vy7EB04JjQ+OI3SNo3swKRBJv4LtO6/HFJ1IrdSTSc6NPQReVuBn6+
CkEFJv15mU4NB4iKdmRq25KYwZu6cqBRxaNLiaPazQKxnz/dxYQwCJZ+Fmq1s8KA9/n21/eIu3aV
LkZQJKqGwHZX+ATatPIZ4OQHcQU9DfQa67zWnfc+zyN9k6MKLdpyW6pc2Ia3rOevPc2n6hEsx3FS
2x1+Jmpf5rKZaQVEshfVhs7OHzh8j4jmJbgygGNXXnIKMADMHuYHpcF1Vtrm/OiCUOWC2HKXCOWD
v2z1TZLWAsVtrCQr1ecz66qC53kU9vrMTHoaYsYsuqMx+X7MkMyGhWzeXcDAWSRb/KhQiZnN1BNY
VJ2VuuAvtowy8FV+X2V43+uu1qcKVsAq0od5kkcDUe2A0rS1hQSXbqa+JzbEu2tPsVCvqDdlzzwU
wU8Nfz2wZ74a0lZKVh0l4aVQuT0GraNwAG4AtgRrQLYMwSR8tWWTXLPGUP/I+ZGBnhzvCj4/oBta
tJuVvgJTLgzw/TyXyHOJFkOkF88AmI2udyXTeSYUpyTxhQNZ5Zn/STj8OByBro53ADe6SVyjE0It
xTj3HVhImiWUPHMczy+FJk124K0+G4EwIePXn3z1FKaCAB/FBnBLeLPzUHQSMl/frZXl6a810LmX
f9ej3gvstltJsTz87SK2mA1xjQsPLfoejuIanWHop19BZ5I3uwN3RB25Ls3rCQwVvAe/YeiipyDU
KFC2eHduk2FyX+XinH5UpAYpGdYJeuDF2X3wFI8ZDFPd8YIPnMFtec+MblPSpLRoK/hmg2YiYDpp
oHhNIHEcvy7FuR9VcoFCyEpLhkWxbscsPH69octWteLYRBqftB3xedxYTAlqQSSAde2kO2NTZJ2T
sJCua7GXyu4+TYzZ7F7H8qG2NluHt0VlYpY1ojvlrd7TI/OFm4R00xjTL54AXHpIzbFCr8l+Wwby
yy0DRdzMhA8lQmRpMyLLkwhU+ss+tRUKMa/D6/RFpGUuTulfgOcJY8Zlkq1O6obYZkBobMyJIe2k
MmNLbMjoMkUSzq9IPZpx2SdGxp9XCpUL6Pco29VmMIz2008elQKLvqA822C9+cY3llLgvcbC+3Fc
cYVPv3iJhcmNddEwQEC4MzXLoSHMt1xIVT6KM9hsM/cML/UA9JjfJU1F7z83PJem8bL4qKNwYwgk
7kfXucT+zM1SUsfk8FOa42KOWV1bq5QpDCFMwlSY52IQrJZv3SK63nbOP23axLrTabHBmnerVuhc
5OsES0riK7IoqhmNT4LfORe1+fuCqcbL67hAuN0ttuZ8JPMA1kXcos1AEmv3hs5qOtP4YqE/TsgS
Zr9TmJ0oXNQq3742MHEKSWFQLKYNgNAGbyBqFmQ6MPw6rRD9yJ5/yIYPFka9Utjh/oI9R/5z43sG
mTzq+XnZHbaYOPumeDLyUxbFkRSo8J5oOCOocSECRpA0CZbQ44wEwizGACaMIDEIorBNPfC2VwfB
eMQ6vng6H+3NqEVB1FUIWR79zq07FBaZMX5Tcpd6/echZSFmEITSxuQK9TNFXHe+SPUZfeC8TRaa
79OTEyiBwIr6Sb01lS15v9uBDLHZtPGzSbZq5CFD57IvoC5cMqjpwL8mXUzlhjoVlg7R3lgKZAgY
f8xwFeekhs5v6T8Q4J0BB6EQ4MEF2zt/80o7mbuDLvvvBrSZPRKJxAFY0cp4nKCX3kWafEoUrqXz
YEwjAvITpuQyqhM9RoB3XRR6kYp/GnjdjoFMST/S+nVkbGJ476WUEbX5COM7kDCVCMFHsApc9PDZ
VGRTMk5p6rSaRfQ6//Uf9L4aGRMeYw6nTH65UCB8N4wHqcIo/Ka1pCqb6u0U57HwvbNM/0KKhWfT
yhzONY3uqThHMwcYudFoAZilE4NfGOKIV7ncTsoeLDweEflOh8/vo+P1kId7VyFkEeslEpjVwyoE
4OdZ/dUBO11aTYqdf+oPYvPmxvCBHt47YgEXT1Jfe84l/nkMtk0+Ss98SHrBzUuos1K3Fzx/7XFA
LCqYiMa6lqkVEHBqiWFpFN+8/QwiRz4/aLzL3TH6lbAatQajRqM/ey9L7Zfq6Sp6H0hSuFKKY0GI
N76oRjzHaEuOe4we49r6kZOdd22IrWup3D9SY52yEs/w622OM7CLU1L0skGUjDw8ehjDKDtQn/ac
GIxxiyhuSMY2hqQnqsw+KL1EfCCs8AIAFj704lRKGvOKvNwZPDrsYabv1ioT4v1jcqDhUF95wXgS
MBCboUO86eFyBCkDshftynWVrOvo2L+xmJJxwVQZt/2yfsh0hun31OcYIVz/t/u384j0L9IyNQ5j
P7mdd5ZwLHKFyOqEIpV0A1w6fhn0scdgO3Eg+Z11hxoPsAPqRu2rADxixWsOx4Xgz/LkfdZgYqB3
wT9LpFr7dn+QVvRDlCiGeceOZ5+6AE0SuwzkcfvSJrpUZtPTziID2BUZAfJ9+vPICX8jtwREtNXO
T1vud5Y/PZ16kifzwWjtCuzVMZMCk82ywt8mO8BSue0ornKs3yecRkGski7BWGFy0hYLch4VKrPG
pxDamPYgTuCDQOZgSWlRzmdB0RSPGortLMW22v2mWhQ4sNhh20bZWStTFEJGROKJlONr+ETp7vg+
dtTDJJLTTbgku3NVZWFBAyOL5CY+phVfCxE5z6JPn65hRSofCXhWI/AruZQKjEh5lR9ADoT0jjXu
3L74bf8GMRFr2zSJ8I5VLkn9U8Zo8xMWQbrJivwJm04wiNMVkgaMKvs5EOgoXRQPRoItrKg9DcWF
8kK0IiJhgR5v4VpNK7gCUUEOpLuNIubj7yYNtlJDnPz91cuMoF/NFtdseSDVylJJfnaHDRDAVvah
qznTz+a9XQVhPaZriLBJwvmYuKADPMwgrTsj62lHzOLKNVK1ek+0zhJ3TGWLjJRkay49FtMYWW7+
lPujZ9gmsTSEDfdKRdAxEtPX0ch/oBJ0FbgAits9RbcTH9WylH6ATzIixOF35wiF4yieQm7MBhY7
NanQjmw/c5MWFncWijZZLVr+EuRAce2zSaljdYxGw/ob2SZ6GtOoHX+z4BnT1aQXRDqda07XzdZW
jKkt+tZsxJi2EdZNgF2gK0OK+XCZj/kTOMAzO/59UqLq0w3MSYFpsEXIiLueL1uK5fAkBPswCcM3
DMVWcR5y0Z57r0hDY2wTJqBTnCwticq98wGfcL3uFJaoNl+nQlHvoQofYWho1KcARS8Zh0jhbeFD
QSlBuRH6aeL+i2FmRNiLg3IHqz0N/yj80OI24wBsRl8FryjDNmohWb7VZqDOXy8zsjHskviryiy5
FtRMw1fpSMBcBGXsziFxmyiTX/ertk4vZ2sfR2G0Lgw1XWk4kJqfO3Qt9cyTs+7os2KUuir+GCaD
wzivC2SmlKyrAP3qhxuM7pjEk+hmKC5MCfeTvpCAXemZrlble+RXn854qOhNLTbOm5xwKk9PZmG6
twhf0U5Ryd8nhIqracpx6E+g2wArivPs/nlY9Nc4Pg6zh+UTmANfHJKNOD68fNS3/nesnBbQydNZ
ael5CorXTosyZjCgIxn6HhAo+d4w/170eFnqMMxE4e4leRk8bAj41KihHBAdRk7/MXZ4raQLOHAR
jPcyKLsd3UCl0hnyu9NScqI6OuJVxHiYOpo9DOgEMoTPYMbnA6Cf1TAXPYzvQyovyQXhpf37EEnz
Q0dhFh+dv9EcmRb0AjaM7Y6pHeT1Uk7u/W09/JIaqplYpvbfYmo3k5iIjw54nVm7f95WR47g8CNK
NJgAeGdLSGpyMG3XauibxbrqlwOYaecDocQVHWfcrkMtgtgXWeu6qhowgNV2aAmyy5yYHlOxr928
m8Gcj8GqILAhVWo0mEJWobKeT5xx3sGEZuU0+vf1pT9JCXhNHGTMdJmufVGW1U6KF64XUlT4TINl
fgGAl2JRmB+cde5fljSm7AZgpJTqSo2zhgnsej1VDRJQJ9yPDXUPE5WC1I9QDmxVU1mxKYYVlROW
8wJiY0cdA96P5wFdZ0CZDsylTcl4SX+2k9hJiV8VlLny1RyvtXzJTiTl7uiGt+XiA6GKnkpHvIQE
mbj/fDcUZU93bmZay0wfH+H5J65EI7cMCtkaVbZ4zqweEyronO8K5hWh6UEj/CKf6nYciZyBmWJE
H7qNb2xASGH3WeWTgdF0yxH1y2pte0KBA6UAgxNbr/bWYIOt3JyDWyX7HRbTrzz5GChNzSlfJMV8
cVhxEcjRIoourqDEGzcebC06DWEu69hHpKjOFovLft9WDJIqf3Eqxgj9YC/iXbZngXKWG838OLTD
Jy0GTljQgWEdIbNZQliibpHS0W30K0k0IXuEgHThBt3U3DbuqwwcRd+bQgpkD+zDZQJ0Cz+i1V0Z
ef0r/jq0ShWVOLxDWnAQsQBvzZPEhR4nHBlki/HTETKBBplvcifK6drTYPmJFyrEVLNnEzbbjAaL
TNtUioyNH5pwQ8OpS1DB4LlkrlwxpyGjwDD77f+R50zlzygbImTsWZO7TeB0A3lxi0i49XqOVdKc
qGp8x3Fer3IQeon/0XzQx3DJZzFppN/4bL1//Qe5u9b3t8Ak9NUvR8gs6Bs2JwaVYr9o3W38wRz5
i6rehKVuCFNt6df6bO4pnY84IxPEUCN3I1xbAbcafb65gy4ctJjhh5GLs0QkX+Emhp1fVg0qvpzH
rkdbkeVkcyfATY7pFW40q7//n+addZx5z5qcNHZOho3SfpPVt+n5S2Sl7U6Wxnvo0gyESoWsiTUL
bp3rll42zo7u0cUexiq9G9OT9wv3/xqrhkqjdPmSv61JlfHGdaVDJyl2nxlly8+17xVxRvmgg4rE
w5Jwo1ajF9ZnejpSO5mGY39uDAlL+h/KUKyTLXhyTu0g78Iuhefm+eg7Tt2kibup2loPXtWec9bG
sbIEGmN/MHBEOjcCsuSWOeKq57V0vvdUUTvX2ozPXgKh437YQC46Uh0j8mpDHoXodfqq/FRvn3EV
mMsx5xKKXqgvGk9OKxPemDqQUvVvM5RdVWf4VZ4+EZdlexclRZGcd6DS/n6vlZzptIVj2+2A8L/e
esttizgNjFkeYB23KaOO7okPcfnQrOONbDABwtSKZ2vRoJuiaIhLHxzbowz7VKzkcCiPSJXY5/Za
pjWEkHRTIc0U+G+aJcbP0m7rPZm6sVg+I++rx8v4DV3Cv0W5S5ncrK0AMt2v+YBXCvnSZjM6QISn
zjc9/TB4OGIIVVKYS9b8immuD8mRyjsbnw6ksZalYIjmzcBBXKsmCYuYP6XQPMFwRRgf9rpjeIrH
8DaAdSzlPTVk8qZII6KrPkmrJo7EaqR8h37UC4oHBlqH2EZIfzFqIEcNazwUH0//vclTYnWCuNTp
teFTuYGuHOc1IHkDfDtIYCXorLSYAp20IsejwtgkcLWAFtqxHkV8nmlT2G5FWRFVSUfBDtYOoLk1
IBfO0BHN1t5vkCHXy2d7v6o0Oq7WwW2fOSV9/5+DdpEpcUnaKDFY4DeAsvBPmm8sK6lBXJT+4yxr
TZO5boW8RqsnUay/x4syXtIeH5l6BPZdQidVyzP1Wl77poiPSBJ9WckFAYwMXQFkLXAce6wIIun8
/OkaVpZfzDoZFwypGdok5s/H4Yk7AA0zwIzEvMjDk1E4OgKSI0pwgqgxELVNu/0xohC/io20JeG8
Ye8omQzz2Ld4/l7ltYgoOr6zKA2FmHzxv/Cw5IZ7whuQakcl5GHn5IURdoY3vzBkWSQ1VkotzI0P
ZhtEKndPjqI1O1clQ07LsxwaawP373dgQosmEb88SC5W53PDEpGV1EWE0hkF8OcG7PSdwJk7YV81
JJAFAT/JN1EM25Yv6yM1LKt9xf7sdu06IpSZqeoFE2VpHe4osEVH5GJEhGf7FKLkFFmucGCNzMUg
tRq4/y098S2T+pNO8bvd/g3TfZDluVUhQejfuHzAq0+psyHEvucm1dSLIJHIKwkAV07bPN0/SPRF
8RzkzxLWQgejFovzHbN/wKhQ8c6X3cotybFE05zd8iJCPpiBgdpkHbUXxRxHwtxuIp3rMTI52DBo
f/FjZQfutwwJfRe9qt8ybG2gFP5+LTuotOh+blCdaJTKdQwsK3thDs8NDs+AV0jJ8ohf/E9E2mKs
EpsCckVpJSS+lBfyX22rnW8XvaT7eVJ76fgss4IT0/gKZwBY1iX3o8IQ53lZuCyjaRYALkimN7Hw
4EfDgpMwLFVXYiUcf/c7J9WyoAOtbL1epsfI1123A/S0HHWafxwmXR5ZdpjXkQBXn+XX2F7/DG/J
pfJJhrj5AyREBimSutM8+bhkDPTn7tVy5bILCW9EphCAvUMf/KV2qeX83+mi+ZmTTOYoiPbIe1+y
eoRGon3ZaxCasjLWsDUiMMLioCEy33xgeW9iaNrQ8aHTAT0oPAqSyHC0iUd6vveewqJS976A0RH0
zqk59kiNJVWUBS3zbhCWlOkybM6+8vci9ogXkp5W/9TAIU/4QtIB8BOhUSuUpAOl3h+K0bVNHL3i
LuGCgpL1bS8KHAUByWdjHl2fanySg5C+6n7Fk1XCUGDe9bXQFzx1VhCXhRrX/eend2zvK0Zl9Ac9
3va3PNf2BdgXrGQKpLhCbEF9uICWMKSqDfcBLi1t1qdLweu1dExJgE1xujz3huCU4kM5xZAel9VX
DSIN5Kang5jTsrNZaFG7HCY2sulbaia/s5TEUyAjjL+VdvZBKd8VNt23pyzyRw9PrGmkwvkBhEhH
p2nji7anKbpu1RzT9vWQpXIWhFoudkGEOYxSomyS8wPMHw12enPdOJo9jJ7qWqTTrhtv6x4J18BB
FBMGA3AhJNe09Pm3iBAFYBp5RS4dGMGD3e6w1YbS+hy9IYFfcL+Y/6Kk7U+sLObpKS0FhCvz6m3c
AcZsSVKipDqzYmuW5U1D+8r23mLbdWadF3rRZ23xcwg2DKFgLmAgPUV5OUeJTB/IyTSuQSG1k3t+
MK1wJ69V/GQjHndGxKPrwATd7tDDQ+F4ELbi163uWOoGkKxcFgu6TCp3NWfcMXLbTTucllzkDwoF
i5AESisvgqPZcl//2QalXN9x7Cxu1yv3pFyEdudgjYcyRwCq3iFsz6VnxSlyaIk2FXVXT/mgwl28
R5N7ELgsq10Ox2yWiYGjU7tgiHQ8b2cbRHO2665n3ygB2jlZ3fnRarIRGPODISzlRcFpVN7N8l4U
OhSNrFdALzxJNcgFXiMYcJXqGITqdUzEyPtnIMV0cX+iufDgBTMV8WVN7d/0NvrOr7KapRzsR9Nn
1vqk+OhVBcnOsILtEjG0tiOz/OY7roeK1peKlcI6neWl+qfXKCvaJo8h/tyKO1mM3jnBwakr1yW3
5qfFuWhhQAql0gPbQ8aY8RU8+aIFD2XOasD4yWib8W8jRdsWSNz4c0e+Uu7LW/PGp9CCtVPVXDiH
5Sc9r1pmJQIqlN0C9Kr2dXuPzMSCPdczDzZHUE9rdK17QgMQOKS4YPIPgfISBdOZCr7BHeCfa3c2
kqwrWAgXjoGxZwswJVOrs78KIm56Blr2QdHp4eyP/MA9EJ8S5ClAtLfpbYAqTXwgZ4A+pQGEZhFL
ZGQ/dodqfY4tGFdRwkfqpI1D1yRJykFuJi6Lh1DJ9knuNSDDVOPLuH4yLLQ1jqIaYPlYtgJv9iPW
Uqr8/qhxipwj01M30rRZ96AwQVZVuPBEHTIJAKbMZdiXxmfUXPqpAEf8zOviCP0cOdQUMFjQjGvG
cqloN/q/AKMJqmiSz9aW0uYx6GuRxwAG2TvohqbEhpRoq3Ku+Rv8+n8xOd1zAKlPLhBRI9JLIQSh
3W6Fzve3/Fbm6ptjjL2MDqtKrWk2EKndbzqt6a5oJtzpvTtNjdbIWhIqUV4IcFSZXMw6w0glgj8/
vWuc3HFCV4jGf7SJpZO/Z9NoBgMt9CYklQefvDrdex4M1umkSCKWN9vWX72krMYpMS1jQpYQUwM9
cqGYCA30XRslHWsFx4EWKjcMlTkVcmVS7uqHNGr0sh2leY4v+ErjnQOZ4sLt1AhUEGrrazXi5CYr
VcnjIDTi2zb1QG9boC2m3fY1khxrIdg5czwWlt9vCtQDzmiCc2Dre2egopHBFNsBNo6Lb0pHPmeX
Bg/iPmLzpRITf02+6My1s+8hSumijZoyRItn6lSOcwPZbM6tQfSwp0WYijMYvM5eYeXU22f+SyWv
lTU6toIcFZPISyGOpii9nXi3e/fG3W29L4XfRq7cZKpbreVLrhDjq7+UUxAJ4yGyQwExKiJHP5DH
zgrOI70YnXrByXjDnUsERkivrGPP4F+SNliou5/Dojbocc/kotyugYGdJKDkhpxcA9k6JuwB95mX
kdyY0k0OGoCmK5dIHADMMovOCJBj8PgA+6o5BKU8vhRgCMpP3Kxwa8Pan2QOuDW5fKEwl2PY+mOx
iQQAKX+cj1GX68FHrA4K3+LfQU2hthgrU5/cHle6dG8P+Iub+Y8XHLyZdZawrPrrBMgNvVVnQPEX
ErVvbppuxiSfI/LqJkVakrbPjoulNYgfc5mINhi9KKPAj1i/dfjn71oDkdrnrIApZGNRJNc/fWf3
N7LeaRgPNyiJYfW9HiYYHs5LOF4V6kF0UgjQKJP25uolot1JC1hgxIrhoH5gXeqK4W5eM3MGvC+H
prSbw5NUo9pqZEq3ahRYE8u8o/2LdRbcy0hX3dzyuKvU9IabaYnH1gJV50GRyrKwqw0t6rajZuT4
cStqKTsuo3X8jbTSUEfgccVpyswjORcvx/fWen+U2KhmmIURMQDvJjDoHXL9kWnxSOIJc2ZnYoN+
v6Df5BdUxp8lKCIuwMX3z8rFcsUttK/A+jjZ92Duhdhv4dxUTIF2MSmY27cnFS5uC23U9rL9Qbtn
vW4y5ZBjInNDuv7EChzP51+3fjiYJjcBWiMyWAAlK30UMP6KpTrTq5tTVZScuPvwvf8pyDNbKZ7S
6DI8XXKxsosw6AGcDtmGE6MD8+ppeOhutnTQbe0ERyUIr4LV0Gs7RQik4GuPbOuctbHhLnFEAq7W
YqQ3NtvRt1fBzxiH/HXb9uGI7t3kjgJH0P9iByoMyMV82d6FRi5lj++krCZq/2voFzgJjqNLz732
srS8CqItB4ACWrFqOZ7KwlJJqtIkO/ZWej95/7UcuEt2rJt8yZQXLIpHGNDIcHKGEDF0X2ZnQUEu
mEiBHqJwiQzGbZYXieBDPKHxfd2A1IhUYS6gjPu3qoKffQmCmiaI2UnX+as1coFc31KXn3Xwe2Oy
RgBIQ9z7YJvdh61HXtQUyu+MG9WLLngl0iiUQrzxvbH1w1r/iDnnyxs7Je8t1LGENJhn3eDIi/p1
B5q1VzJNDyvpsXM/elnoO6WZ1f7U+9pPPsxg7fCKIkVgE2PMXvD2zfuNp4oCRUF08Azmq7oBj+6d
Cj22gal3EcALbQPEVpzvqmuEJJMJNiIbq56Q3klo85tAfFkcd5qWjBP2wYZLPISHb5qw8jrAfMIz
LaNcCGhKRrwSdQ8hocPHuTmQuJ7f8WGavnWrQjW4WBWL0acOUCR495ZMBODs3UWjKgVAq4J66gM6
OdBQ/E49wUDiIoedEN3w8SaTGMW1bQyBTv9gJ17el+Y4kliBNMJRFqhS/15wLPVdoc1iBZ/yXgU+
MhrNyKCx3Sn+dA6EFFTRmbXy3JQB4PJ3LZBOeZr+a3TRM2vzyQI3L2srVHkeCV/3HbRyyvQSe4qG
aQPGWUOYda6Gt33xbVmupWSgHv7wY998Uc+ypEXN1eHa2JJQZj89sAyBoOwYsJJC0xCnXMNB7J/5
2eVXxQkECNmpWImyGAJWrdrntyrh0A7aeFqPJIiILMPEmjakGy9NnVz/8LyVj7M2XR4xjYZUGUDs
aKxtnxJGCv8z8bUUy1w1OUum9Wn00505ZPF/7w4IwVGy5y0VSL+dW64/n3U9yeAZ99fi3CLbr+1/
ID81ATnqmJoOf/imbyPJW+W5LpwWou9ez1E6wTNk1HxKffIJm4Us2glXHLnYQyjO3TZwl6cWufLH
S261hKiXI+G5ThPufzLUskJ0fDE2raKmQPeY/+1ecxUb+4nhKvwUDsSNcKtN+PNDox+tTYh5vLvI
flIwNMEmlEQq4iPfgL5YsLFFCvEwKwWwzVa/RvoBwhRdOqXQ3TOQqPsxIEfc4cs+kmqYSDWRMfnY
ozvJd7nxZYGiOqBLhRJl3FBNGIu4ARwdL6ZOGaoY0b+T8qJHfAAsxlI8zappJ4AuneXrbpaaFvak
8puKiqoKdh/d2r6p0ODV1/z/7++uUduoECTtttApK4k5PRWWRTrf0RtCjmY/tnb3aHmbEo87nE6s
t9iPSWnE0jWyaHDlWFZqNKp16f00egyMXzo/5PQtT/6b6VHqyqEv1q+UleBHipvTKxXPGpO+9L+8
JOGVF4TRbWOKBA8zqwNHSzOIGCJoWEzESnJpehLHcp+yvfKdkq7hE/OBEAmuPekAR4HXJg0TaEZr
OiYZz4nuE5M/wC1RZOkH8WL9tYiobZOyn9fAokx++evsXvN7AL2BRnUZoQfPmZGvZ9gpyaR0m0H8
cVVSzrcK5fQk3WgbmZjr7gyDaoRlPY391GoZ1hs4VyD8mzjCJ4k618qvd0q3Sr5Im2hbgXUXvIsj
+yG/f9jsqMn/9sip+NIQZsNyjH2FkcXK6P64ZcG5gsTTPPLCaao3ywnCBSmsvFvdd9xvtLCR30Uv
0Vb50xOF+DcF7dD1hKaiw9sYuVRhXD5fAuzs7Kv0Y9/8TxBa/V9tDq4z6Fa6M0gvr6kR9HI0gJGh
GJC6Gujnsxh72omPPd5tm/QoNVVCs92zOcYskkUwq7NrDgQbxwKOYIQ63oqj0585s5NyEUaRHfPO
Y+IFoh2Zhd6ofL2gsDu4d1ZJWQEtHv7Pq/k79EfsXjhLv/uoXVO2EoE1ZIzYRQzWavwN7dCnByUs
GJZ6dr3sxeoxw9PlZ3K9j0VXO+99Y6HYX+C/Ope82zRcfdu30oeKslKDZl/m1sHeS+bT6TIc78Fi
z3trkemXJ1KHuDJ63Brq4/zQKEdnIZAl5O2gc5/gccpzeRK0bqQL8xA4Yl+1mtRsTMcaYRhkJtYm
2EN3e/6AkPawQ9b2y3hkxJbUKgmA/QIokvgQdXDp8Ps9MiUVHUHDoTliGOdP1UqJB4J76JGjq7OH
83yHdzZ4UTYUSf/NVDb2v0HnkH2Xo10dUVFVh0Vz29Yu5+qFZSrY4VfVUcpSuipIR4R5oBFIY3C9
pvD3ykJg4MF4MUCDzj4XrTbm+y3oEvHcIKZskCbjFfZ8KXBDZi4io7DYCKSTesh1oBurNjb7Gv6n
zsTTx0OWbe7vTtGKvs+fJWYdtPHG5NkW0ECsnnnFmAG5p86KIbaFnuXrrh2W1oOf+f8jgKlApQw1
5sSM6dD8QJ3lSlFQi5wqervOrW4lyjMaXnwOpjjtIogJm8WgjcxyaZpiGR3aUltc4v6/Hfvxq6Xo
EqoUliiFoaGH6reOgKPtpaVGy+MJv+jehS2P5wTPUm2/65+qYuk21haIBWIf1UGkJpd2ssSKqWS2
i3BsYUzqIQlLyl704uNT1I2I5T4N36J6DS1dfcmDySzfofolaM3lVUoTxdJej4aUqKckRBUF9rV/
b9DSt5nJevVGiHzIRwQHdP2Z2F7eFHP//NSp/llAIq7RNd21Lm59twh021UcgCl26pUCu2T978pR
xQlMPTahejHRv8v2YWG8AWXnEqZCnfDmLs/y5Okg7KAU/ZYqpa5EiKqvNkUz7eWu+AKdq024tCN4
e2W75ixm6x0vSwx+rQso4IxyuIv20bjOoN+jPlnZ5nUbF9obRu42bHkzX3/4zSwLdhO/2nm6n8Gt
HX9OIm90SYberHJ4z0tdq8ZhIOHZXZWZGu1zqzJcrJfcqBpzhRKkiwyicpdgqqRaTLUuwWnxMrj7
4YhTCOZ3z7+8KwNT/k53SuhEixXWjk468AFWiC4epfFmBGmIVIEoaaatW4AQ6SqrP+kekqU2Sr/3
zpJnufZFo6G872x8u46hngKpL29tvrdmsqqfC2FIvoo0NfGK0QNAxukbEUYMi2pLFvQ2boStMV6b
8D1vQKi0cc9NzQV7eVRb6a/h4GrtpKmYYzDF3TaD00VM8TQBxCCxUpSBkDXbydd2T+hqZJUg4ksm
EYiuV6AhQ9wvriopUNnNXWM/77wSBUqlX4YJ2UCKdm85UIh5SkaPGgtRdEXV4qtwKTG9whb18iF2
TCH3wOtVNM98ia/spMjEr9rh4ZMkjKExRPnGLF5jzgXLcwEsuKd/6S1jA2MkvuNEgzUVbXVkuOtA
mkxYV7ocnH4VBDANHt7D3rMkp0L0icurp52OKvhHDHhRI+tEmt/FC5syL4iOLD/cQurFWXsgTm0c
bb8sFr0pNExNyVljON8Si6RYRzUxrUtytq6humxwnBoo/ztPrwQcsjzORg/P/zKZDcG6a66JgD5B
xnKl/+h2lZlFLJDrvMwQFUIsxjgtX38gFoWKl2cGq1QzajHdAEmB88zZ1YhqUCqVaqqhTPwyLWLn
fTeZIPkySd9A02EEgQpASGYybI9+5QB+roZGEQwxq4IYov3Jx+tIOqymDQLBdsNEwzNQMRXfvSYg
ozq1yIGqJTz3lDfLEKu7CvgSzACKgwF/SLMGj+foi9ZqyQ9QdwWHWGg8v9/9VytrHBGekRh3ptsu
6ofkrgLxr+M72bIPoXCyax+Ds1Jm+ROVE7vVGYnLP5hHVWERA1qpf08QPEXd4ofONN8AIHcZdYOg
F+ezbBRSwuQpJb4Czzgtj6XwZLJ/1VKz+OLo2cyq+Yz3Y1vDg3DKXRVTRSowulsmeF73/dIxazbS
OIxl4cQCkPyyQjjkt//y3ywRpWj+2H2U9QtnLBCQnv0lFkweZZP4PitLFxTavtD/1bF992fGrLRw
DkhnQGEIGGFc1puUKQqIA6tFGuCYGczzZw9lHY8FgxxGRR3SjNxUIe2DMV7nW2b4eeiS3lWGckRq
OxseGXBVRDLfPHAlh33zVgEx8KMeQwTuP5L+JuBBL09JtFjXC6TO5fXvrBq34ayWZt+CO+yR8k6f
xmGg6hY+xS9KChQlZsCSkkPP8V0PmtV/ifoiZBe9IAlirE1CENNW4sz+xXaDHtQM7jxrBWm8tqAS
l6wH3vgatxVy72Qyr05OWVEaik4GNG1PjCebgUAQBRdPBQwJCmndzQgZUH9RThIKKpPzDVjUyzu0
fp3ZWWQ9MeZtaI88YlduvXMAd/+XsFA9pNHAt/Hk+soks1j2gOV1pUH61WIg+gRjhQO38X0+u7ZG
2R9p/sRB+n01nqDcT3E6tLNaIfllMW3spHvMzj/s77frgEcXuq+OvBlzXERG9HOqFMRN8gy700Lu
MjFAPeiM9OwCR+tefKhYYrgxGC7RwHOqDsBu5N3Y2K3RrSxfdfuzKIZSYsTUyJjKRHJr75aFv/IS
PRimdjZ0/kh5mnN31LRsDIgOnM4LAKEmv7pjQPaIRK2fBdzp6WLGL/6MgAzdxXwVDBC50YAHb2YY
SVX+6LRDKt68gjJfz6I1raZ86h1b253bdnHP14LGhungqrK7daIm5ZjlG9sTu8PcYyvXHojhf7MK
F3kMDDbxz1V16fFh3nTg5COR/hosUC/XZM+mFc52VKfUgWZUMQu+zWtWU4cgOIo1+9qbH/HpU4mC
D85w2owfhIVMTukaHfrdVDHewi+l/sboNpQ2OL9RGvdWBr+B5j3YDvN2DpXLVMV2vGnn116eRBTj
28c5b4qXd6EPQLJBsnHKk9jBZFrkEXbCY/J6Bw1c7CPA2hKR0LZrY3TqQnJd5MY377miCP3KK0ne
d664ma32mH3I7ebWNSwfjvEo4WeHPrwToTGRR3tPWfB9Xf3wYmeL7TVSWSUSnuZkyZ3SdpA8I8mj
tiAJDeAgj2Ol1qWl6iswnhGKm/cJq/yh4xp9R3e52THzhR61+ukOoLo6SLqnsweKlR0pfGxWV+G+
rF00D2YxmigymiYPCQ5pXkyuM+Q+7KOJc4D2/RybTpsiRJPp7y9cr9ehWsWYf43ocHrJwRE8X10P
31VNc/0sIRZkV5BAGZbB6tSrf1n360rzYKPKEaSXPMdBsbETsJIpzmeB5n1L83iDVjRgSrl112/q
A/p7co8W6hbZiUlqiiUzQE7iXAPLP3P/eVToIsa22cTnDOrNvrxsDf2ps97cJZXwy7ePxCaZfUvi
1ru2NHXdNlygtcnodESophyXdrkCuYOSYjviPLFk4TTU88HYlCzT0up7lOx2MhkVh7IwW0R3eEml
0YwTA7vR6dAA35G4sgaevMLIxJQi777bIBN3OsVe6qXCHi0YmWeWocm9inMKdR2VFSfpsXEfdEku
NLwME+d65rV2AJ0+hVPW0tqM1hIqzOGkf8XZY4fn4kSqOS2Q6Q672IpOHDx3ggp4B5+dNHLc8L/q
jCdKFTs3DCVVhp13nVGN9pOqURqet5bfejIuUkw1YPSdR7MtD4B6AHRmDxfZ61n5r00vqo2UPsPM
dD5waDAONlhyPkvMDwtaq3eR6PU+6gvU/tt2sqewBXVa4P/Xz1y5PoxWUaX1VdAGTjnAia5nYLfR
99GODlzSfsSpqdEVJT77Z8/UO5tceI8iB+1JyVr9s5as+wUEidPim0h3fpMVzkFybSMVgKSCkDcP
l3Y1lwV394G7Zx5g3sqY0yubyy3FQ0MSSmjtfPRqDgV5gKv3IY1zan6ZKhWmyjnmXjeTz0tGRwi/
opMLl2vBE8GPJFSjnZ3ZWx1fwmt/puOP7Xm25xtz/OyfDoqUKUaw31DDpgElT1/rpe0DkI6FN5ij
hwEBKSZ6cx8OtXUJSwpgFhZbpQtEC6MSjdpkyL4/PjPFCoNplwEGMypBKzfUl8Ii5dhfkeDOYE2f
wYbNdmnSnCITAZSE1XYwbrtY+SZYPHUby0nbTKAnvXNY5YUhnsyfEjMy3y0nqjThFqvcymW4nHgd
WGxHvxUDwCldlPUneOF8jIlUnzxtkeofbuecu2KTGqyg6ytBm4rCU7palPLyhYpDJeSKQrJy8VM6
USW9Bi34bYbuJwK1Dn+M6nvawGmAdUxIKzrqy01oqj5/ZPHR08VfzUdWJH3ccio8xkZKzW49wIdf
OJrE555sHOJYauDgJYZKdmRLw3XEA6vKssm3FtDZl8oB1f/Bi2rmQSNMa45FcWE/y9W9Adli8/WD
/4UAoyp2NsDPSUNpSikaFZK0DGzg7tND+31ozC1rW90lTwqLjHvjPN0g8hJFhKsGx/pVRi1XSTgJ
Es+iG0/eub8LgAX05eOAHErwS09Dxw3Yf9HrcH3ApRu3Xeiy8ttBgKaXIIFiGkIquif6Inm52ZfT
PtLvxKyr5ZgavrY1/WXQcy697g9ECzsi7x7UBkFpYla1ZAuXYWuDpEk2Co2lFE+idT4TAjO+4+Ob
5lADPWF4pWfb+9DVZjQk67Q7QDQIb7JuPL2jQV1i8dWx5mPV0bb87BP8KmS+oAE36qvNKOEwikgU
v+J2kDB5K7vckGV4WrswYrvQRh3czTx4on/dsaYRiiuQYO9Q+EKo9kTYL8wUUucpzmcNB1KrQDlP
8/42ccMhqXvC+anrvJ02XT+MmsBF8jBu7+6EMCn28JlYeP83OJsdSyusAD85AqfUsRZOfXQxKBUB
JQWoD9p9P7tJpyKz5eLg50hLrpT/bAl93fAVnGDObwQqXbRyrBaP+kYE7Mm000ZjYeWT+nZEn9fN
dXiEe2HsKXNginOoX6JTZA36RnNGDkw9RWJDDDEEZl1n+87eCzWwLON9OFL7r+gbQp02pkWMatr8
pHv27RACAex1k/WIdr74Fry3DM+/U4UClYD4t0ZT9SrcZC3AIQY9Ch6Li9Xmc7XXGgJSQlXEax15
gt0xKAqgaSfm0/0bRHkIDIWK2WKwAfEIjfQhlv6aBzapBLNPB0ac2N0MpzNzWgpXRZZhglANLhaT
5X4miKO2sZtSlpZg4nj3GBVRxrg8L4dQMmrshsZ15lDeGXNHKhLEEwjAbTD0eyQ2Bl2yPJ+8PBjz
BaeQCfWFc486sZDE++wlv1b2xlYdIOJcSruEVMBMV0LSL+ugOiTQkZqZ1m7PhXXK8GN2MSJxLG7s
dnczS2v75+lxZMBOKyn/4pK71cOrKJEiojmVzgfHM/vCiz77OuXyzO107sA3wnUEMkVEZRrruNG2
xuJ6PHWlY0flsoz1YwlVCFM1Tjd7uv7R70lg2isWW8k1+hXuujoLevk2vRiosAdMQ6zdMu50ryMH
1VEEOio0l9b5LbAO01HjOwgpO+Fbr0aA8hhntRzTMcneFraGLNkh4WlHYJE54jhbN1SfCX6qSetr
Q/Qh2EqfUxx4eC+h61lMSVwZoPFAIcifJwo4aMrhZ0GWrwka3mzCT+1zewYZH8DSOzjDVWV3YBlD
x+jlM6cvsLGWKZd65BtSUZU+0B7QgQmGGLIZh/Gi2UFjdJruQwc7dbpBREsXgnmgTOjkidvduJ+b
55KnZLmFH5tEnH51VkRNwc9bA06pYHWp5EnlB6dHhth+8rhQMI0xTX3j2wrhDeva+gvZFbTcOigQ
9Hp2ay45Alwd0glSnK8153HDxYpZsiPdJq77GYkRB1OEFExQxxiMxhosaYbg/TDhU+6U03C366/G
Ly5OW2RrtUzrfBpgIuvUBKlMoni1GksWf+UW0q0bMBrhgg4KXlyH21glZXxp+dcTEQUuK2px3/QG
WaRSOpPJ83cztjGeB7fjHLBV89Fz3OvtWt5GrKs9W3IUPzO17VFOK/DKivdr6amlpU5DaLyB5FqT
8izQDRAd9rWd23+ylZqPrZMhTtM3+r0pNa/Yd+r00nK4IH+Oe5DIc60TI5YoabK+I0BelPPFON0K
FUJ/lUlScgWvKYD5GSOuWK7MbFnLJv5/nxwrddPI6C06OXDscLQ+6Z3iv2HyyZnFP7f5vAcXLr47
MF1tTLJw0J56boemMi4tbsj5J83BrseST7EREIs7kI257SLbzqabRnwHXEfM/YNi9xyfl5yc3d+J
cuNNOvfuEN1RsxB6MGOHJoR7LAQYJQNbG8oQ9GGXGWTzXRlkNUAlwH6dpSZ8el5jbiARlVJLSN9n
kN6oBSF1NkJlNNLO0EnE8akplXO3kMRJqTnq4QL9k9pBCOc7iff62EPBkCTQ/SQKD2sgFtSCQeOu
0GbZMUJQ/jpA/P3iMnuBS8XttdubF/2o/BVDd6k8IWxwYo7ofA8O50unczitYoC04F/H3K5bWpQ5
U6wXICfuzWiOhn9EkJZws6b91S4q2GTuKJVEr2TQxkoecJkXKci11EImy5cSPKWszcLvnWllmZNJ
flv2yqpbWPZVhddUTQIWmLbE9W0XrPcNmuZAc6CPq1QU07kcoQXH1z2eGURMnH2YzMC5A+Dr8QKR
21TF88EQmsyOewUBZe+hIcPLBtb+ie+8XNlEGMfMDMm9Md84cVi0wv2NUULOiJMEf/yhaR5o/s0N
+wf1Mjz13OghQgh3sOgSykHjP+bLAuKqEMbHmQvr0JdMmK9jKyfpxxOJR5KcbYdDXUpVhdGSJARM
K0gsmnGkMTBWQucPrpUR3fKeoEXFkO0rr6M8LG1m1ksmwD2GtOn5aI0aS/s3a2GngvzDs1fO/mBZ
ZdFw/ysSWuFXRqosG4x+RCHGuSALh/iA4aGr2cAuZYp7v0IWANJJ24RyxjPrISSf1+Si/TDtNTzr
yG5hxDPPcG6BYseUv29DJdQIGLmKPmFEyae/JsGXklKpbfRPJSSmIM0Kj+FGp3gg0D09axoWuot7
QrawmyyKSmDdQyiRSXKLJKO5TLueBDxtZ6UhUH85e8f1gEFITqGKTRxsmwhl+Yr/KlFVsIrRdlhc
bRZ/qbV/UZAmZQJTyE0n/tO52dZODqP/I0WGcsIVsn9YVD3IlBsQ2Pjx61WimLvuM4NycSV+OVuC
nYlL6SaZQnBuHwBYngX54gExgY6mFKgqGEk8T2LQmykkWZIi9mK1CRD0PCHjaDA6A95wGDblki1K
Znj8rmTT5dA2ySlyF9nhOPIfskfwNHaS22yePnEpckvHTiv9JJWXqKbSO7/+T7e+Zc4Uu81dqIoN
GMkHQyL0NtOFxEUij/lH47CITSzKNN1CB73D4G08AsRW/aFbQQR6BYSr4wf+q0rsRGTTPIndCUHq
KE1lJza5liaM5JNUq2sjSRgYaG0qde+HpgQKYRXLfqyMditpw6cPm8HeGQk5s2K9Wti/WTck3dVL
YLjn2GQybI2iuIiF70c3ZcE2PT20Zv7cJs2gRzloowSQumtkdbD1ttuz92C5mym96IqMhbwEgLqk
b7piSMEegy3TjGmUs0KXEL1vWpSV78tG4h+CuflbsMPe6hNRHcAzxR84qQcD0RzsLbYQj3gUGkPe
NFfMoqu6R6QbnUBKPpcVqz+qI9k7kL39w7Nbfl+s5qSA8iN4NGmE49VkorerDaeJDT7F0TdQjpoa
M66xpIjXWckYseuBMKHnoZL0a7xnpEEUh4CJ3pHQS49maknpW5ybyZeE0d6KnSiZRMyIhHNBg72H
ouOYORwP8oLZF1MNh0kAtMDhGEn9xTQ4nvY1ObLmGPqlMlx4tOFk77+x6RJUpOCrf1kZqaZiVK15
GleOspUW1NzLzwVNHQHX1swNEUE3Br9aE56YOXi+UW5B0cddHeUxSF/TahvnqWjq8Zq0rktAsoNA
7Am++fDjxtbzCFT/cA3mFAmwl6l15WV6un4dVYmtGns+at+IAtwHjp9Jp2fpBi7SfC1nh636/Wxr
ZpMkKYh+FFS1sGp6K5DrhozAA/OXUF+SeR1Uek7vg164MVkIWGQkDLYTt7OhvpP+1XddrmZA3JnQ
FQQdXN6tGXI6aCevlUEKlV7t5g1jfLioXWWXcYt+mclwmwzCoMZxgtjRQI5NBB9b7shSkbMfEqbS
9ZJnXrr04bfT1X0Q6r8iTjHlreOiezyp56BMa1O43S1SBpG/bJIe4jtVFezBa89DTE5JhtcnfMUf
d8cUPJe4oiWBjnQQ8viA/aObs3QfkeDm08ySCKwmH60b4QPy3gf6FGDSthYYAxkCpSEQpZSK9/Ks
0sBnAV6yhiHw3kNY7X8IOdaKagC2J2dywclsbeux7f6BGvCTHowxsiMSJprRVluxbj1oyzQD5099
uHShyvtY6y3IMH7/B/3gIXUZxcRUmBzFk/m2fjTjQsLSNDTibsy3e2InAbTP9Lfmh71qJL5HIN1i
zqpm3f+TIJQccdRIqgqVCZYOsuI7DQnQgs/UwrixZeKkGvqOzLY+o/gvGMbtm8BaztfLxKdqkXoU
8/FWxrvaSDHkJjU+XE+FmZgYSd7bS/1Flkwfm8JUCj+e+UHUT9O3b/iklzGNUAVwNRTH9mZZjDu4
BJrXt8NIq9LxlEZTyJuXB1J9MLffPS/KsYx2zz2YySkzu+qNRJDHg33jgQxr82avqgf40sGg/htH
xBia2fgoWo5UgPrPEYqJSjWO1dhZNFxjrVRKS9FgM5+GvSk2Nubb7rTNj+6vEJguAc9o1FxNyj5G
WFWp46P1373gtoKpESUNOISDdud9ZzidhJ18AeESnB4GmXYgHgCxxKFRJEL9GtLhQAc/jmqZJ5hv
Znej1jWu0Vb4KcAsD4UsVHDFd+LHLr2j+qHF7QnwqgesHPOZI1q0FI1YLu6Ci/R0eZEvbTL+N9fL
42hS4037Bv3oUjob2jx1sVjOkc8oqG2+Oz1itsmczZp+16HN3wUPyzRbqXLM+cYTSWKY6EhRW9Zr
MtUO4I99r25OC82edZ1iAPGAA16lkEashokWHyzCCYX14NZGx2KYAQtAbGd6CJZk7NNJN7V1F7Jf
lvmqgDXhKYreKoWNfpH91tIX2av3vnSSkS5y0r5XYIMzw08/oDe2eA+WUCsjIjiuySepph16ZVh2
M674o8W1pHTnZw4/ID0cQV3S22cwRL3IHsSnQB/WQtvJmc2bo5YRDDYBvHLfiAu16IX9iMGYFqZl
+VBZDquPaptT0/6HThzDpTW5sgP/pksxv2BAfmNtD7g/DVL/oqDQDuDw/Uj8zoY87LzUqJvEUgek
TpjvTtmbEfOavue9AiRD+onEd6h7ItQEqsyHT0KgzjT9+YTO43eGkwROPHg4CLYIxP+gVbUHYril
Oegtz6hBaCo1JgKv/zow8MJ7wAgmr12eCShVdXrsCnzTkKqulWZ5Ca0PRpC9T2J4lm1EEbLbrlw5
htkQDJgjICY5tBODHmdWTalJLHtCkSTxMVpOqv5YWjqTyfXP+quoKT4+lRHMFqEhrgsFE+oAEm6Y
9Z5f9KAlg0TmpgUCrFImlmRQdZCqDg2JQwA+Iv3YF+QVFGMIojcqWbRWwMWNwyBSSCd8djl6y27F
3WQxogIGenVy4He4kna1YpV9bWtwgxowL93zCMuN8YA+n3WTVhuiQqMMaeljhItes2hnqu2ATq/2
Mqb3N1S9bMFegkYihEmfTE543fa2Guia8NGecnGqIjot+r/C7LCBqfhsSao/6Prr1sALS1gVKwcB
KHENr5lxU3XsFq4AVv3LJptCBfpCpR0b7QngzwymddSWtaHQw51n9lI0XbB/jl7fWeVOJI48exfd
l5C1FnHi3PO/NtCwsJgwgIGtPdpm317aysT+oonYE4IcyaBuHzOf/PghkfqQG2W0Hq+I2PeTUKdr
olcSpkZeU15950lJ7PEPObmCJ+dkzqfqdyUAfuL5aSDbvmndtfUdtt2fYeS/nbyGSLWLMVFgKB19
MmSaxRHGF6uBtNcKHO/cLInK4ZCbVt2E5HEWzTHOCPIl38nMUJCGC2UGkdFWrwbbssoZCr2rQSxx
2+evkkaAX8HuKCpEhsQqZTGvmT2NkK+OvYRtYyJur75foioM6O2Zl/tR20UvIPC2tXoWlKDYyaSB
KXbKk0iuUXG/kW//T7JGVi4y9LA8v70gYj7hZGdJtCO094iraNEjofsiCho/RJGlDjN/kC42X5YT
zVyNfJZKjVtfOLIVz/SeAzbT9aTXk3ZRer6xqOwOIdMnlRjHqbQCApn3mDd+hSHnhtHA87eFFtpx
ZIK3aVxxe+sI4Lqa5ctzEErSm83X0mo6rnttVVwK3ZPItO4MjpJ2mIhAJCCtpEMtJPg0RS+Pif3a
BuYS5oBsvIDYzklkR+jrwDn/vYq4l+ob07jSXeqI+PmyABQac74EM2ky8gRlYIHhja4Ru83qCIKV
2JAM88HQD8B5zbP/1KanH2yXwDKh5b8x7/6QH21s0QdKeMR9NAwhK0UL6QkIkGE/IkRiNKCFGwVO
rBbJ8tXziB9l/WgPHquRxpY9mjjuSbsyX/3pSZX4B2g/jyrdGW4clXeUCDmc7egrUSXRy6urwMWC
h6gS/K3AAzV+3iCfNXKW7+8ZasFFldBSr/foc9jAdaGrvqtySFZol8B2K3IqTqkOAiO6g17qp0pj
EMiKU4EOMth7jUJDGAn7Lv3yGa9XtCRKXyMjgoMbDlthhyaordBDFPt9KKYAJxZn/XE0iKHlH69W
f69PMxiCqaAiSfbzkfwzNgHKEDybOGHmyJS31IxKlFjiE4sSkYz9WkB8GlBByivz52oJG7ESkVN7
iDtoj0hzDhF7Cz1Y9aEdP1CGSjWGW58n1Q18drSsBvuZlhHD4zGq34ZtfHBorq8rbqPjqMTxY3N5
/zHAsIvqPmyeXLQIU3bKAyGAC8yf9CxHYVQHKV8S0VsyFKUzSz0TIOFIa4npsQt5Ty0ZkmSZw124
NghXPsqikbJOywaIwqV6I1lgYeolAadab4CZqC2s1V1f54VCVYwuYKoyI4L8dyig/FSR1IjRE1YR
8PqC/jI7lmx/tg2D/mMZt4UXV1WAIKO1wpeJRYo2wLK125Lopcjns8wbMZd7X5r+YlzditjUNXi8
elSHvbufpl15wnLwxqL0ojuuUpLYXLzWzaZkD1a3PESy4xtNo7LLViglfNXHtiXUb8IA3gYoC9Xf
a2QJI4fl+teueRkx3X537hJEV9LFEhv31TyUEzu7rLUr1ymEdOcsatOgfBL0dqghiPIhQA/I6HOX
v25M5iifeAq586DxkZcDJiunqxwSq+XMV3mNXpn7M8AGcZgwSTTFpeEXVlb2eUYOszzTeZ6hAeis
ACbBVmmAZTaKSJLP/iKomc9Do3TrJGQvUpH0oeMXwpyE8A5r6VCT4GrDhoZCg+KVokTodHpinU0T
S7FljWHp7CPGUzpAwxZQ4Vzglg+mK+GUP/gFdqKksUMa64lr5I6g2k5TRivQkMasyDSKEKAgyZ/V
Q5LIyN/5TmUTdLp/2aAiGxi4A5JrQ7jmD99KxOr/m62SZE1pCVRxnskdmF13Z+Ulzo9w6Ya0pHLH
iT7Q8DIBJhegyxDmUgOKhqrrMoXSM9utOZziCd61kTMh7LRXYwhcfOweDVIw9FoU5/9BYCfvZq7x
PDPUJp75OWPTjEcX+PtwO6TPYOkOmKPM/1rtdCpq3/2/7v7sHqziD38vzfXugEgGvGJYVHcfoAsK
tVYNb3CynyOne7t8rPsbTGdd/VtlrKNHawpRAemFx5Gmxj1FA5JS1gPP9uicDdjaruw+0SBJmqGY
dpO7sbPdFU37+3XIcpBJAemWc8ukXBbrNZyZF4gW6Ise5viYMVWk1eavuMEd5I+CfmdjZBvcvoAb
vLHyiIMdD55shmMJUn3jaZ7BvU1wSKCRtbITmG+QIvTgFyhMjgxt7h68jp7zks0a4qJ7RyZr01hH
70xPTjHbsuqLZHRYWsJNoDzrrK6ByapZQDf681487RY2jBCgobsGSoakVx/8pWw+MtJA5PpzP3D1
widu607jja68CGIYt2ZLBVpPlGEOYEx8VLUcbnithfkKdAaf7/a30BRHz+kYRhAhYk6nOiqwrJf6
yt0XBNaf4ZnSc5K9ZqLFbkWFoDMLl7foV88RvAh7n+ON5VfhdhW0VAT/1Whoan78dMlB2oR4rhJ7
Sd0Ds0klq0/6GIlzFtSJbb1NLZgm7gMOhis9SVB3i90xED/mv3nbe1/1GqhQ8ZeqxAWlGvVJZfOO
JHi4UwbWfr2q+9yogSoyOAJfqP46toYYgi4FfNlUsO93EsYilFGFYJuf/mcov/MeZhKgb8m+2sMY
Q7w7ZgGuNZ3Fwvk0mtvUBZGW2XaFTmG8+z9IhVpSJQ+WEEm8zn7yihKdtuTZcYSJp3JrK0ezpqJT
nbExWDKxDmWx/lv7f/0v3pxQIvAmowRewFsuaufXtQJi2ooc80SFvNR+HXQ5ogMuVCA8DhCcFvO6
XrpaXj6nZe1juk6zMrDHJa5WF1hbsc86agyqdhNiA4WnzhbIlLeFwXGm+jke6qfhUeoEmB2RQjZ5
xoIR9WqLLK+8U2YMeFwaZGIazi5QqsW9n6vRFqwjQaOip/Pi1KRyYmHGoxfOX8TSItTNAdpyxN9k
97ek24QuTSpGDOddd7faREoXPt76R7UgITJdEntOcklnTBvnrrnb4epD5sGyGEL8Ck05kjtTTMCz
EuqNRM+FJcyaqIkDqzWpBcyp2Stw7C4Ma6OTHp6aSXwpfNnEjqC+8CodCnlKmmta/zFwi+1uMmBb
UQCygGagUvncL5W1GJiKp2ZxX36/foLzA6fnPFLfyQkkqvMBGX19HAHs1X4Q3x7RzSRL9pzHtoeW
PwDV+z238Ua9Zlet2cJpc9lSnOmyaQSmg1QPG0yxVNTpw/HgOKGEahLycRvyb2MCB6v+dDrXBYqP
pMe8lX5aIQuTy3WC6BNA10VJ3uP95Q5eSm/OM17nvBbyKMEZT3H7kM+66mmSQKXM0OsLZ8YsPMme
BzwZx8Woia1UIh7C34Uhrwgr2FHy0cb5Y2X4SZfnf4VgV0UyZiv5lYszN5mbuH02AyzQyvDElzRH
Xo+7eg0LxWfXN5silRWV5ZPbCLsKj+U5tlGjV18NOgrT8GZ7LVcCBWBUZtty21Cqhbm/b7Z5ytFL
tyUd6Afj5vJ9eLgll9BLyq0L90bjJS8yjRxTaBJLxJTh1Ze1800Z6T2Hsj13EXNgoZXLfYXBpA8a
jTRddyK+PiWVGVYTR0o5gd3XMnVDnmqnywoiwVygIOoVBIoyE5IEdgeuf2wVZC+0DWy1wpZKoqYn
ngCst9wRLU6neOhKucykEyBRH4B7DRMV5Mb0Pcj4nGMfol7oH19NXzxONGIku6TtjMWN7mhONnAP
McgpPW95pq9XaPG0YsC8tR0conMtDJv+DcgdVM5IH3MDmg61seiOE68Gbuy5mDzQg5O7kV21NaFS
hW2PoQ5A4nS+40WPcGV1dvAxuZ9AMHG94e1QlA8ZOuwsdj3q3BJe5+hEjviXFb7rVYQUvHZkMd6m
xu5fFdzwHdDDR1M38BQ6vSqfrBznoNQ6pSEvd58HZ7U39Bg9b2v4dtWe9NWIM2lxqUgNWk2LtVzX
AxoPtZUqiOwn5Tb51sniHLI2qlL4Hm8y5tfHWRM8Yrbw0GH/SANcp6dNQtW7YUMrUavuFhuG7p+p
kpWek80FZT7dm9OZiUQRVPokFub3M53FWmFb/DVLGy7J1mOhE+5B7O7KF367OQwl7FG+t+K/xhNS
353jPxwHtuq16sdsCKiHwJU62znmbhOj3nI9p2Lv5Wfq4Cd4yP+Px7tYATyjwkn3HopK3eBh/LcP
tJbvocu6I1HJGABBYwt8QrpgaK3K24scFOP2ABkpUEKllGecxiyB+ZEt33iuhc7+uKY6hmI8wBdX
BK4OR5U8Q/j6S2N76Y/FYNVlJAtj8z5Aq4I6loWi5S2re0xYjlfNDZo577Z+OSjkDwb8OqCtqSY3
WCpFtzIPAuSQEKwsmPxnte3Eg/BaE5p70BAqutbfETiu2SwEOaBrHUFaq9pSX4dZ76lPoc5CWiHI
ePV4ni1OUbos4x/WjIfFmL71+T+2YGeXowtXYYmiJ5hnO69nXC3PEM5Ix4aJdYbZ6cvAJMwY3wWs
fSibRSAScPUbU6p4jXGS1shU92bmgfVZexBRXFzcnYi3JL6H6VZ3k/T+zEDx+Y+6Lo/wiX7QiZPo
eyse4/HG20GmOjuyaTl3aEmzlzZuupWOLu3/mgltLIWDUHin45lt/7cCY46THFc82sxGTFNKEe2V
qTAtU6H5NCCX+o8VymDU0NdOUNjvLBi5D2awgpSIQHdWtvrOkvsUc3PSvO+zfXHexFk8nqeqjLbX
dAoHCVB0drxlb72n+rYskV3I0bIDy42WySeLeMezacCJXl3LdoexZkr7SN7CQDiqGGDF/+qAsdgK
uy0BglHwweqziCetj64xieM/Wm8KRmnICLShrLYwiNoGOrdvLrswif/Qy+QRToLgQ1SgIdbT7eQB
0oBIpU3Rj8LRHxqhsCfFnJvg2jU/UsOjWJzTazwRO55iDoMLFXxN6kGl5Ui7KvP9qhFLN5BCU+Eb
v/Z2SrmokhxFAu83GsHvl7VRSg2LdJG0yWk4m5TOzDCRfEo8PegVhnQqoj6s1kyglDXc9Ej/owiP
B1zeqiulCDXxmHyxQBhwUf3iVmmxgUgVdtQLDUYZE652AZZFm2JWD6aD/UneHijVLR8Khwd21xyT
0WK52bfsKx/wKXZlxIMCKVG0IChd942/hCxif9nJoVeDpdtCHlUk5PrwgxmEN+T1SvXg4IFsBbsF
QJGTtQzF4psWpLkn/VqT8080r9vKCxR93IlNiz0qrtY3iD9mKimznDKYfwEWPXVQ++XhxaDj6hJ4
94OnCrMFrbmUfG5QQseMAinA5XzSkQVnU0FxsC4G9u6/lU7ZRo9gSJmryPwBiu565Ivdp1bk65my
Gk/x50A9hL/iAHTncJal174s3NxW2owu+ujcsiBvlH8rpDRlPxmdNj9a1O2eAFNepOh+/q+PMvq9
8+IcmxLeGLTZ4KfeVey/+v79RtWO1Iq+UbXkJ3b/KB3i7JlTwUs6VzYzuJmaF64z/+U0pWW3qANC
2ewDdNxTubzM1XXCS8ivW81DFuExU+M6kSVP+WFhop8fC3NId+RN7wDfiE2Cp9uiFmL0UJ6WGz+/
xhWJFMHAmGG4vCLqAx9lb0M11pyWvIyuN/5Q6cjfHf9RcWTKubIB7J7k+VgfKdaPzm8c8F2aeOVv
WEA5zbKBOPM6n9XWf1dstoPhcoCymRXAuynIeafYAbveFAftcma8CO6jWLx1jbRafko1S8PW+8Lz
jmHWdDh17aI1q/WRn9noKQSscz7LK4vUrUL72bEdg13ceUdjqtSGpmNb8qxTg5zeQ1srsuwSKZKH
O2M4UExw+aOTyEzDj16TotT9cBCgaELEPsLePzLn6dM8J5YW5JNeu/XMSZxZ/xdxS5WJ9RBxy9Hk
REVf0oPL42i3Oo2vywqkDywuV1qmxA4aNy+LKCGQeTMc9cHqZz6BBOLdEKx5pW2jkqinl0g+DXDg
wBIa/MFa4pCupO8K6I8nBJQBsh9wEOYBsZMV+MrCRWJGvYoVEMRMXh5/lipkaIIP9LqUPXod7GyS
iVZ0zRCB5GkSox6wdDUt3hfxCnZvxNhB7ME/CvYQWZqn6fyMJEIo9eakjK26wsXhKftikthCgIDn
Nxc4ZSGaT+lur1SjYVvsLylbLg61WUfKR/8mTYt5ylTE36+C2MrlAHXrjZQbDT0PJzNMUX6kChSB
m7o+UP5Hjy6a36tmEWWjUyyVBiF+ie57KRtVz/G0ij3QedHHMJhr8NXK/hAWgr+VLV/fDZYsJqpJ
xi0jawDxSyrZe0wtamzmAeDAQgcKVP/iPiT2x6qtUCOON8N96AU8ClIYHOmWWf5YzPLhogczBLBe
0/LokdvO5ndZ56Nrus7bnqqj0SuF2Gm+K8A4Krt4hUH5Wn5Iz+UWQjHwUTBX/1wunYYi4wbBhpzr
yXvkOiJo1xat7SDVEEoT/M2PwMvcJ3PNyHAW211CruKJBarVKoYHE4KMoABMybpx/V3U3GcGKfzh
G4T1XsJ0wREZhfNGL749yJC7IfaiNJtZwg1i6d8sJUnu/DujJwPGorCtfcuLOIe9TcFkIAl2zGjG
vkpAGDfQ8iaDLCO+jVEAOgk5JbzOMwmljXQQP2MXJcn96B8bLRyOV0emDmsIj66z0TqzB2Fvjfq6
Lm2OWWyycd2pVFMBoewnrqTCYc0GhOUP5JWFmHwRwl+58eJ3erc575Ujs0tpLALX5XHNPN6Dse+5
phHi/ZQLtF7e7X3ggCqEZiisxA+iT6Fx7hKFf7ifrN1YGz3orW7g3gz81Vq5P4h9nHkxT8edz/+y
yzpMpEc8y7Y1WCVT6CoyIMz2jhxqIagOoDmJmxM376SyqVLwbihaFu+3KTcWyV62A71ZHDW1jmyk
Ddpa2cpX2TyKMDapSUX9rxW9L4BbAm815uA8UoiR4xKZvkfV0DeuKRMXFpqMQ0hp/T+UVfLwnrip
LNDabHhXgDzWkP3LnkxMtA8YLhi+bLXJERLOTvRYQ1SpCP1QNvWBn4tzO4drrITxrFhy8ZDQaP87
63yinxg4QTb6cXS3wM5lrZLsAJNp1MyL6CnJHkeZFk2eyLLEM6kgJgS1i/bHfhXPFg+rnPwZ1r6f
ygyiggfBtAE3RTFtrEw0Eak93MHp/BpsqC2w4XSmdn4zUVnS7P51r2FD0dhD7qxNswwt8s2jVXzx
OWnezGnmNBcSSb4bXBbVrZHpGcR/jmrKvHLsxNhZTAsxmfPr+jQYYMZVho5b5fcYjjQz5IAcz9Od
QTw3MTaNOcub6DyjPzOtISwE4T4tq3m5xkK9bktoDQVjlEBc3t+YBkm0ERSt/CPZY+1pPlXkk/JW
SjJg568grwap7PyXmKx+4lK1ml4WlKLLJcwzncMdzLll66o2okWXMDKvMxA2oZhuQZy8PAw4pnPe
N3omCSxwnIt8DfrnSpeq590BWSy4pcesKwhGNJqQe/hKaa25rsy0oRyvCuuqxPty/Q/lM8wCqp+k
s5kRRgcWJRa6jQQJNnOM4ZYmI0Jqc6Mx6nzJeAVDSErF9KtnpuC9gfr33vGc8w3oSQnwDdeYbd+k
Z95F6bNwA4mSr7Gym2ZX5drJlhW9v+NOn2cTzVtfERXyw6KO5VAsAYyc5AEq/CSLhQcYbVvItcWb
gnoYL7VsEU/5UknVxjAtYkpbbAo14OAMGOP7FF16bvjXnavR9mHQdgFOtUbiJWZtqfnBvrLhMchw
inPT2mi2d8HQHsU0pyCywA9eaY/TVK4mIudxuLb9i/a3ZUYgZoiXVh62M+lmcT6EcNEZ6AuAiIZI
szZQT3zl9g1ESnnE/ZvO3SvFRea+1JpmXkOm+QV/a82lCiBu3gGItNWqyN3AQze0rc7TtGZTALbS
jqfQsbMBY8TZNByonpL0QeI+nFlV/sMpVKWnOjcUp/KCpqrAOMhJr73OfpbZ5kWwcgAhj3AIzaES
NNXlGqwTTFlrqBreXxktas0Oac/vEj3OoOLvWcV8nnEZm7AOGc+RdMPFMEPH3+ttsHktJ3zX5U1B
bX3pdX1dwW0KdW1TyT7uJqdLQIn3iIULrv5yUbRpPHORcT35cJxGPeqdKLB8PBUv4AIyD4ZzBfQ+
QQRyZEA3QWRIXwTLgZeMvXrBJ5RjwMg0gG2is6MevBzEUpGDFPIzN2z7eutR8VK5h8m7fMc2SzAF
s9A9UJVFOWP5lnsZeYtBIfn2ya3QBOAaxgGqUEJ65i5HfMbV3EmC75cQFqIgTyXwrPph6hymt90T
sOPhBtgkmYAvLXVTjv+MQmhnY0r58VUbw7/+UgUPlVnmAeP2GI7KZwTjbrAx7/oPeFOgE9DKlf+S
5xHwhjbwxJmL+fwYPAw5TyB231QdBlZpV9Q8qyYf4hZflqTDOXGkJCULO7af89SX/DCm4mPsDMHq
e1R+79uydq+bcMKmNxaVXRQMqGbxaLihHtTIbGElLlE2hezX0pGrs4QsuJ9L5TCauytcBFrrI/W4
wkKnL2i28vIZ/HHHvHCUNPXLX+1u/lJHWgbYeC0CoTZh960gZ/9QSx+Eqp/fyXceg7SxQA5OlJTY
UOXYo9vjBjw6uQrhn4M1yN5xeAp85iUp+V8+p46IvA4nSs/wMUK6PIiVQBpJAs/C1bJiXKTKEC0z
LpRN2wrFHXpCZh4+ijCdTDaLaZgYSqRvUQWfHQ1GshK6SOYLX63d5nNKbe2Xac7iha9TwqfDl2Yh
oNIv2O8UY3N4fTx4zDC7Q1ai5iKj605v9RZKyd55ts5CRFzvR4hmV3bxcrvdbUU0O4m5Zjdzk1LH
6GnExOpPhds1YXbNf0r6+H8FN0V64EggUdJANWrQgAdlWnxcTwYNYjm3PbUCoxFkCXjsSWgWAS2j
p7f1wMaPF+82EM3RD0l7U5NUBCqwz+jtCXGWEjT5mq/J+NVO98PMoD3O5c4+jPp3+wCKnPXTGJOG
GK+Y2JCnzctxrbJYXR+crGljxw3Jr0sOAvI3bhPqdXfmpo3nw4pCQ3z/xLcoWBHKv1iTDejRlN4q
FkMj+X8k/r5zTRwsBH4we+95rFCX+Ee+bhTXqjyDuFquGk396nezZPJP5yzVMSAEBSsR0MvekzOO
KLzphOwTRYy72RrJqciSeAfyzCs4zdom7CNSn8dAmUWbkU2Qqie45ZxQxXKUHWdtVu93N33CItAQ
x+s/D1dLeNy2Ymw67Y7wmEro9DuBQL5cMStxtFXfz9ZSu6ZVc5UnODP9ymLLeMYRVto/3jUyxeAs
IsKk6feVRznQU04R+6KmJSOh8JswNhYPaGD2ROfyehr3M+u2RwTnaf0keFlNxWgb98laBp602LzC
Io5zQuswAaeLRmdsEziiMzS7pStzVlMnjCNpQ5Q9pFPj7Uu3JfTetoO2SMBKH6SLJ1nz20j9NSAQ
cLLUMx1ZVVJUQ1SwaSDw94BMjKaqKtu6rWxVzMNsb3vdzfjhOnqa8tXUB0NT6emLLdWFr/avHtDn
260zUpDRj5+EATJrbUYJiRZV56JeELVW3Ek0E8pMkD6AmiQ9Qyo/5whCY5eqZCgm3TP53AZmcIu4
PZFujVY9CxDhL8LY41JdNx/DMh0Av2qecvYjJN2V5tGnzvNmoSyuWJnGCiTkNfmgxvv3L6NJPlkt
b0ibn5djtfOrOHqF1/jtz/ARqnAmmFzlWL2aCbZlhq+qLHhIcpwTP5oi4XUbcw4LkSJ8cdhuKFKH
oEySSZRyWS5jYCTDS5O4qW+pS3fl5cwDCBFXlRecH9k/EUHlKyu7BFX9KVymAPIEUfXzN3WUER3q
BsrF5gwa7ZlHPRovhraL9sa1I3p/SjnsRYs1Kxnc1J47/I949nbP5OEN4AMx0ab/O2xlEAhHA3Zo
4LnYMFPOROHL2wMvABNOCSNy3Yhu/krU9FMlwcdBHkQH0H7usRbRICQouseyXIppA4Tt3TB2DcxA
knhx7S3vMeKua9uUL6JshaJeZELYEhOTuN6fZTa1ygleEj8jysn2ehN8Wf6b8QaqHLC9FyYj4p5B
nvzJVMuG6rdYKxbR+Zl+GJcS1p9gxSc6nEkr9aUU5nPPQCCIqvoY1lMXPknUP14mezk+WgF9/3BO
lHbZVg32ir6eZ5Xvxx2PN9bv27fuosqvIKa7Kz+0NQqY0x956mwgJPe22BKXRVALy6d3aC6jBZNt
eoILwsyoa/tYFyN1jbhB+bIoQEpkAtG81QtAElntqc+RYd+J+iZ6NnGypGsfxOkZ95GtShqyqmxU
KybASb6pVT3Ta4AYsW706APbd7b6Su8hzfKLEzf7PQFeIxRPijYnvXAg1y6Nz969ArMJYRUgLzTi
5UtqEC5biLcsFk3gapDSd+7B6ExfkTN2Z8/4/1/AFQSrD03xEF+Bz+cP8TD83SahyVxOMAhXAb/6
xwDbqM/abJ31T+cbwmx4q0B9MMKdftkaVxu7hmQIkKCJ7K9gAZXBdMeAux/NES2letaBuKqyt56X
9DxZlE4SRcGX7a/xQTaIo2AbzXbuwcr/FYju8ZH0KTckbuDDg/DGx2yu42QPS8bIRO97B9g4JZyN
SDCrikUnJXkbRkxgUF0qytJ0ynzrR7JFd/AGqKP10/UNHi/fsjUY7FYcLtoE6ptNdpsdMalBEaAa
FiwMyl+D/TYtNVKUA6ugNQnxzTtrrk5EKevLi67JBpZUjuc8pZ7yF4t4eltCbZ9T/3lPlnQZMKPu
AdAujsFi91zMJzeDyPljflTFuINOdCBxYTu/j026uRBSuVXX1onTAVTZXbBK83OFE1Q1QZMkiEO8
fBtIBMu41oBbwE1z7m6j4LEssppXmeenpLNZLqloGY9N0mA4bqFaWwUQ5lepjSmMSjVwTm+91fAF
d8Z8EONsHYGtZppiyaK2wAbqSTPkisrWY0XKZ8+PdloogY0S2BYpMgpaFzelUtUrgmor3QPQXIVB
dWxJiQ7c2/bemn1/zCI0Mh9+2yaQZk+yc1yw8calDYYAn7kLmlAzsBzaKSTK6aVmcqf4r0VOJuYt
KiDNjafGwFsEmod7B/bRoe1qRdzSuhrus+XDX/MFJBxzo35z2TykqRRWdBNDoyYC/LuimK+Om6m5
VjaqyQ1cpHxpJ1/gf+g2QpfnKjBJKA8piAKDvPqddxho5fNKk6BScy+yM/fVYXZ0U/PNR1WpKwcX
hQ14ULVCjDpeJCOLFGBsDlRz0LwVNxEqCxErbnelg4hsUiAksyvF8E3sL8RLj9idbEYkZTInS8jd
V79bAekdgpBLB9XH1PwBZWwfAH6rOVpTxCTuwem+LRpKKBAu8zskbkk9vPwBIjh4GSFRnYCE+Yfl
F4gq3sUN29hc3LaML6Ds34e88BFMrj63e/dXVXpdPyQVYBoLpeMtHJ4ZGrob8HLzrNXBvWO0yyfe
c7iFRjFdIiIgualC6HfOl555LVNontX5EYKCHgnOel8PS8Q38Fc3lt6gdSdY+RqOtHSMAHcGPUl+
nZx4KEKeWpHTY1JUz/EFTndCTEcLt7d19otSVqknZ4ETLedjD+UwMZydSkARFqLci4ibPvWLMY1G
tei2+sNZHyJNdSnei8yfI+rU6orf+cSsfJhxx9MVrPmgCqU+dQIcvKW3Jrn8QfkWRHuQcm+eBDJ8
mkRPf3danoI+bRMGYEYdiusjC2d1gdRCP+W1HqXGkxchiM8H7zsGdVSKYiMw9KeAtuu6w+jebCUR
xeWNzGEsRrXxU5HOepzleU6Q2XptXFLLCHXyNs+ylQNTBS+iRo63uYBR63JiljnIRCN1qMB/A+x0
2qiz5vcA24DlESUDffggMyiRxeA3xHazQ/XYNUMrOoNcPtt19nLEci5mBXL4Dw0jJdw4+ygSItxM
leSlXQ3AU50RfruoeIYud4WtbD2s6XH42p8Czl1UuRitJ7Z1AMpcuQE8p4NtccwvP2tjNQ8Q7a+m
Ttcw5eWYOCUl/6UgTRgrX2qCU4R2wYVfnNMUN6ip7/F09SP/uf/kNkmQj6rpULdI0K83C9OJYoEh
5llz2R7CYEBOAVYJDncVqe0c1eNUvthvNFSHUUWkzwSQ2Q0gBcwfEdjkQ9lp85xqmZWS/BKLYKzt
Wukj4S+l3BTv2YnQCbfo/dT0JpLfuy2NWNxK5WQWVNavD6QxvlUAfI/yYdu9qy5Ml1jsK3eaNFm6
Nk7rL2W+KMARJ4AlJR84/TkTeAOC7ZRePM9iXGvjDg6UR30dHuH2NcyFA7QIFIkjsJJb5UR6t1y7
84HhMAVNlr0bE/uj6HLnu/EyCWG+suCsyvJQ3Bld2tK3tDeN/rHqzNFjnO3/s68k1/ieZteOm7PM
SV/I9lH1fRIWZ2ZmWd8aQOGOOUjnB1CTona/PwPxs6pY7V+SXhnn4mLhUt6QXVDXq8VKQC73o6jo
8YEPIrWpUnZcttkuP6tnxfNbhAGmtWh7URC4yr65Zinv0xQCTo5/wu5F6aeKZSLQuZt1FV8S4EEQ
Fynv6gHtkZcIiVALy27tdR9FODSdPGfqgahsVvbeanQkchvQHmWQsQMLBuzYuPCqLDE0F3aXCxra
nFHfH3FFE+Z9K/WEzp25FEHRZn+tOmlDdyRFatqM9CRjIfzqcSWefodqRIXhu7FwvGylAFbFd0Wo
pl46NSJHxmUjApHpRaXHuKU55ecaYSjS6RmTiv4LGIeqFH2eg1MYJiCSpZDN3YilQO2JvMWGg3NL
lpudpVjpMMRcxpBkp0rYcfx6m9l6HFGn4tZanWNIaBkiRttBLR1VFoxlLD9UMlQ8l64qiZyrBzd5
u8TzoDWHwr3EhCTpGFl9KB7pFPxxZ5Ouxw39WyT2BH14IdP5FIpHiCV17mvi/0+IJ1aCaF1SBNhS
AT9lV514aVlVGh7kHpJusUf40EPzhb+0NdAPQ8rVG45502AAe3WDVQEhVuAemNwRsYvSFA2RLtvf
wM6WuCnS00heD1ANO83LJ2hZFE37rQBdqIn4X2S3J4q1xs2mVRLiElthGzw3wuWnUE7+AtOiYjhx
qGnNyzAoSO7j4prJiHB+gciGdYoogOrWtD1W6v+B9IWgxSV2cW9i+70EAe3PBWoVylPXibj+vblm
2z8hrp774HA37zGkgsXZryUbnlwsyqmxmanKcUWtxEFZ2/WuUdZPkeXF/tiymzQ/U5Pov9v+Bge6
9dLTI/ngtEhC0sdKECw+1OI8RODbHgPMpXbXR3YS6hkqGCb2vHALNNsGKfmQ5pNJEECt4UIWcEJs
8uL3/w77FmrSzBWe5Z4ptibCxqkjsEFaiSq0X/9OnQeT7js7QcfWUImwfmLMGFEn0lXyIienkC3F
ws+UHDcVuS09xjGzF+6ZpdSNlYFjEKK3x18Hfi9Bo/O8ytSK6Gc0RLHPql/rivDqqS0L2kgXacWC
NKFs338Vi+/ULEueyPq5WK//UwdBguk8S1fMkBA1bCcvFh8FbJ2aL6pYN5RZCPwxVLpfDi/+wjBR
/2bTd7FoJkNnSy5A8LWknv+XAclHDJmAaP9+4ysSYkH5dck0lxOxdQ4OWY7QIHI0gr/IEB8xkMYN
vm3c2p1vnUfyLvPBaIyJIV8TAkQy4r8J+0PLNPxlRo842EYfFDn3FGwF0iRHZQXphGBRsOGg5Irg
NkdaQhftHXBYSyfcWnbT8uDUFgwz+k5X42DvIAhEkUEkjNSnemjkqcXl2t5qIDQ4oZTIizfmQiY7
UX5FnouXif+4/CJZu4FikAUeb/QCp5v5Zmi3xM+3/jhloAJo5IZRx97jep1Uzz3Oss54bPBluqrC
2cMCLxJ3NNnJBlhPaOdoFCdNbgnFOaHhN9mY1Bwyjt3JgjJweXtXsQ5oNUMRMhf70hT6WJ9XpDLQ
VrjIPaxmGU2n7OlqvlmTmtJn+MqURk9o696M+il+Zk7rgrx5mJnTghpj6g38yuflIVrecbxY3s5o
SQPGLqs2RzDq65NBzJJ/Fr+wgkh+p/ymFLl9cnm84toZAaW+aqF/RDQ8bcwDpUAsC/RzOA5dfZo4
pKS5wciogXKWmmAYKkfzbKkE5vZCr+8m8UFW9623he/Seg6bK+kZSWtdHuL4z3Y1WN0UTUBWKHN9
SGkipA2o+scJTJmGl1tbN/f0yLuADe/mtrKfyuKjAEKwGfEJUZz9dnTFo1xB6Lo5pOyAWpLjIP0x
77GBUu5i0zmsY8rwTY+1cmzsuwgcpj8cj5UvYy5+EDkkdP5PxcUVfivg7h1pzmog9JV355Z2l1/9
rvNH63d1FGDQqya4lHHKb92RNsv380RwPhqwCMqmlesd/F+zuvSNojU1eHfridseWi1+wnDylcFD
0Bg0X5GqJi6qS5yM2aPjiVOCtnTJ4R69XBmuP8l6lfhboycH/ZZ3j8xpSO44oGyb3RkQP7CaLHgZ
+jxX1GefLoJcL18guoIgOzxzQIcz4AZhPHr0q45uLgS4wJqEB2XxNz204AhTHjC6SJJgKHFGYqUj
13yJznNOKFXiPMbZiUj1FUk0NRUoET1Au//eCfUU4nC1RbQs4Ps7wiVQTHFqCv9ovS3w4TYiZhw9
a+D/pzVJjDMCuWi5Ah1GEmDWZIrmupIUeyTmp47H2UJLxNoDmXKfg9mdzWz3NiFA+IuBeZX6rlX2
HSv5K7frc0XBK2oGjBNi2HeqlTW+nr81BG+y/WJSgyMGyW/jUrlIHkYrwgS/GOeom5LEeTb0NYtd
Z73Hs5CV/JqNQvlGmgwmIlFT/+uMUTNTc0p1UHyctFVToipJyc1RjijIuGn7zWK47bj7bTnYH0jP
gl7zSd5OWZbPI/4TjS5yqfVnQbyEjA/QT2rKpi6/xxHHSiu9Zcdv+4U+zgH1SosXLVIxbU4jSl5f
4/kv3Pi80OlMDsZJAv8ZmCizsfefybdKw6xMfc6HrB0UnhdBecPglCcwNQPRkVSm4MYIPL2eCIkM
zJ91M0ou15kg4Uy4uTDIbdnQvryA2bY3zAFOsv9GiRrGJjfPXW+swAuHVTuS4+LPFkgykoq6iK1E
fqOfi6ZRN9vy9dYUBeoSPdqeXSOACBFG1V76ZlESTMdErJYv0ppSGM5akFuPdWnPNgGCqir3lFBr
zRTVVtDFMUxNyzQephHdVhiJDFZTW14PlgNxJXqh917gzeixy/k1J5SRaPMHSw/5F2MT/JYlR+v5
PI9UR07SDI+x9zu9pvrcwmoMFyQ7ilHWMHpzKT5t/FZ1gjVAI8GK5snDen5LpQsJ+N/huD0gCWWw
FCPAFM/s25D7TWP9PTBjXFzFa+qVAnx3Wed9l7N3CucIcVnPLSfdWzzMhkrZPsQJXIpru81+3Emn
aTVF0ze0B+Y1BmKUT8dCxF/QnJXyvvBTZesxeUDk2Dx3xkCwV+4rl/ZT+1ryiXkcuFX5oaqTOE08
Iv7siD4ya8K9+P0G/rVHYmqlZe1gf57T+i3xBsTrSn/AFEb66ZWB48t9v+tftyVPDcNtOBtfX7RR
m9nOZWjAtZz4sl44kDWb0+DPDFdJr4dcFTnGPG64qVJm+yTNaRMR92cHGhhZg0vSin8v2R+MzKB/
A8pTIvHOYH2LPtAwSGrmRoVxLlxe3xudg8FKtkQXW9BQMoDs5/8dzu0LfNZYgKAvdKs+A6YCZPqW
HiatxOOc39RFZOGQZqs+JZ0OSL7vzDAUxsZxW5LdwxDV7Yj4pf/aaS0cg3ffZgnX7JRTLYKcDFmu
0+0zIqzTKMQTsnqrVBiQTndviTkkMuwwZ9l/ZT8hJd/TIRazZNIhRBBsWiRI+HJpv1uTLFeusv9u
exiWLWEBR1g4av5FoE916cJbjfsU8zfGgzZveAW6RVLX/w2Olfd05mae9W8fo15JZvqBn+uBVksj
RxheFZxZQvGicxvwn3IBgX/tvgxQ8BtfCg/cuHThZ2w5akyZj9t6NiDWpEe6fyx/7B0Yn2U9S8mq
tkaMNEC7h3Y21iyhOFXpaMPt+kR6rocdidFxxa9ZnVjwfplV4RuOK+cfsF0DzIeGYND5kC0dRUl9
zz3RLUzlBXx09tp3xZntq13bpet/vgUv9GQduy3+KACQhrKsDvugaoHYLm7L1tRAbVPv1EHbLp2O
fP28+JHIuhd0VLWYMA771uUoiOWzFplFTcbHvzJNiLhv83996xLR5aJPyzfFgTu9GJSL7k6eVbiy
mxmZNnMIT7QOHPYSJADENsHJ74VUvoWUrFwkWkSwOUPyO2j1PkBrWfm3Mx+HlWsXUi2hq4gbJdwd
+7aT3m9WHAXEZtuiDuS0vklOUmFokwCYE7mQE21077gy6wIxADc+MoUCYtrWK44F4UeBbA0XWDxQ
Woc/VPDY6O8rw7cw8EF3GBLfRKX9NkmNlSExCgwU59ZzjCoJL24GY5smINGSfjvjzJjL07pY3gbA
a4VRxOIZ+/tkMZxptgPOCw6nZSItiT5BIbyY4UzDkLI46ceVY+XBLLiOdkBYxFNWIYVHb6hrJd+H
nUYHBRoLsXcR4w65d/py6YncDZ1f7l8X0AH1thWDUD/FiPwo738TWMFG7r/IFz9v43s75VpjfCHT
l3nS9wksB1Wz1RBmTNcD/DQR3AxLNsFRgjGGB3DSphQX5YZg1H1FAyQM24aGLddBFYjgtvV/u2dI
hGu86K5p3JCq//mC0XSRo3AbBrzXe+i2esru8Rxx0xqECnD8T9PdIuIw7DjCESIb/aXzHufvl8f4
igrdrUvthj2GsL+1jazUOOQDoIGn4srWGVgbFjOl6K0cBQkXpuYFRsDrA54S+db8KIm/xcZaxb3Q
Q8yZFbtIY0fa/QuT8CYbWL3j6OmhwsXS8L+bh07NRCMSTHgPGXU31c7agoQ5un5mXXfUPh1+S1cp
zEk+vnnmEbW1uuD+uNQWLp3LDIYzQArbWh08eRy00mh/OHa3KCU3F0PY4MULheVEGEN2WOtIwCaF
gvWa2AQdcUY+HW0qXz4cD2Pk7VXXdYbcxqNQ+DVyELFJ5s4QnVrlSp963bF3SZrd2oJDLBDSSpVi
ip8HoWwbcU7gfMBmvONjzK7tdpZcep4zp5yE+89bXT/BfOkDwR+ImHCaPMjqJ5d4aO7sUEyt/gD9
eLTonSUiYZxoEIajDlAbasSUOilwJpehWxWiMXTQYYiDham4re+LRyLytfQEn0NOFuFw6M4ydoVn
wGe1dj6ZpGEDj8y+i4aGjy8xujFLOk4dBgtZ5jy4S/4oqDMMZfnUAu5zhicGOYXeHzA0waGFhiI1
V9ww970oKYdyBsQp9GbIhcu/AYqUXV7XPB+0qMWsTCtwWGeLip/CYSYL4+ZCf0/C7K7UjSeVh9HH
l33hlOChNvkjI1+GM/4RCaZPtVd0vzVntiubZkBqu2vZhhTJ1vXVBCLS+FeNxD6qzH3gLG/4iIX4
2I48z8xPlcTXyfxYfvpMmPESevAzdiPcbqI/2IviK8UdynIYQakB/dyDdtlluX+WrzqM/vjTuO3/
mPDQHBhPCSgpEOlYA+DrvkrPv27dSXL7zhk5gHlw7bBkQ20dLT5ewjggtIVGv4jDHx+/ma1CtnyN
uCyKokEiJpJhbc42RwexuRQmDyyEjo9hIXTFgs8JOF4uUqLMy8lgItfxpjjqLTg0NUYC7czy+Tur
7YjrM0T4Xh44fnc6ca7B6BFlp0s9HIM2Mmwujz8aK9UJ2kEDDWulJzWJkVVaAfwFbnpmG7wHNu9w
crz14uw9bLZXO1UY0UKFWui4tQlqdLRAhsLXmsyrUlKlkDj+8EpcSBtXsC8yhOG7UO/Z548nw6Q/
1CI83LpDY53k/9dQItQednYQgr3Tl/2fC+GcfAizp4k3aHE2o+VGgE+QKm3RRgghAwHbzNvq9Ygv
v16+9OvwgKkZQHxzdPaZSW2h2bfF+F++PGXqkYt2E4UIlwjyoBJ6ASMBMz78gWv9f9Sq+CEHaeiq
c+6nrD1vYUgINp2MXxzbhD9ytep3hvhUS2zbSbdC5mYqzC58/ftwEGOBm9WuFMzciXqRXyc3xUvq
W11nsHTKvodc7uMFnltUiXiFwxakhCiRBeiIy6aLDl+M5AxBTXx9T6NJINH2U73bpkKdUm43qh6w
p+6MaCFcvb9te5Q0ycM5i9k/QKFDKA1er1uMlB6BLLAA/nu8v7vrZdu0WtvfRU2K3tlVfOOti8Qf
Mwo71MjPg4tVwf5jxV8iBJxTNzQvt/ZxB8f+Ec7qPWec6v13u9PgqZXgzlIpPwpTuOKTH7O16LSM
IJABKc3ptCsWlVJUU0E6Je1BM7ZIP+Jh/z1n7Xhy6igqaKUzlQGlmSh4W5IJf5OG1XJa6f5brn/7
McPQApi6RoeaNegviQWWxzUF6tbwjlfCHqrev3joEtgxd9RR7OCazKj28VM56fNRWcEnMjAr8a6m
qplTo8HmpVUoM/dHQ7Fe7SnNZFg/FXhJ6gdEamM3KwU9Cg7FCTtU0tc4HUdNz+6GvFd2pfdGtq05
9VQhtH+wiJURH/2x+vW3Sfzvh6QVaO8IQ4bacVKNAyqoGiluu7uf4HX4Y/JllOdF9/JU6KGe7bC3
S+uWa8DCzS9Z+c4hIf2fd/bYjw+88yx+W/0EqxZaxZuO7yfgrtBtoEIiDk8rHq9o/CjWtEr3RBwe
/bUOozsfcTj0kijwd40Ygs9lo4VIEYSDFPf2kyKfDN8H9oJoQW1SJnb8MedDBvvoAzCfqs6BnKGB
kxvKMCknDp8QlJuGpB9W6oEOxx7H9Rt21Yd1lZ5TlXlyV7Ey7Kmcs2QSfSefg1N+i0ehpuqcz7rD
SJWMxsngILYBCYQWG3tuGU3ZHutpNQuJg6gyEyfxHiFCHfhT30hywD+qMIVNT1ZkI5S1uSmadd5B
shDmExq932Fea9mjc4APBKKM1lG3S/b6abicJrtZUaRoHW+8qJR547hCOwxH4/eUUH13uGa4+9CW
eCe9RrTbzat/dMnfGTHePlLCOyK5S00slf8nQJ3Vy2SjeNzxIGS9/WktnLBu0YTp53JyHO4UBX42
xYrbEvv6gEjMVaY4MqS4rybbM6aB+mahjt0cSR1Vy5M6efDRDlPtkU4rPGTgqM7aB9HQHGL41pTN
NVFoG8oZaxP1oxEEqgZOa8y4bxt2LzPiePTKRedHnJNConhL6I6vw19YTVh7i02KrNXD0ZZaKWR4
IboYdkJbQ6Cp897mdF3tz1g6eHt+ZNDROjHXLZz4thMhMq73HzEWkdEI2hyDFK06RF8ggdsfdnRN
Rcxi23m/2BGJbOstuhNZnaarIRR8RSf5LFJhZ6WTG2Q4/rKtyuLo94/eX4qPtJWM25xxEeWe7CRk
jR9lrr34fiLGEHuMj4A4omMUBSMOQswscUJPRq9obXN8Ap2FPxu8LQCQLxpQsyDkVSriCVWSqqms
ecCtj4Aj6l0EwFU9z0ONkXSFLJURnm+hWC4MPncgvYWYSwUSJexwHxx8zsd0otJyRO2udBEM7y/m
b5Siht7LzsH0TSb7dIu3EnU4F2rrrZHBa+0XNhTpdkjMyBsML5PDvgr29tA94Qic9eGfvnmuJW8I
NYZ61mCD55kvbMcHeW4GaWX3j+gfDwcV1clEMHUMEnlK0C/ME5uAFm9lvDpykWGE+Kl8jyF4dEp3
0D27Ex+Wk2KAbgIDPn/iB52FYax7TaDSlX1SE79SF3zekWR/Lm2i4XEVV6h5xA48hGXg0BUTEaA1
A7zPVkXCSFJ2Y1Zz+wdryF6ILso9KsbLxyP1AYmQW9sr5/NJUjgacJO1c5yfRHsLU+ZM4ED+Dq4R
VyWtbZvZ7aQH6XYlNS0Kw7GlPe4Ig53HTmVGKTLbf9qCH7JtOdIEmF0RwrVL8dm101jZKHXq2P5W
XZezMBqtlqjpowiMwEE5k/DwXfa2c7eDvX+3rdnkgYRfl0lW9Kpb63weulRU9Htuj4jNg68mxxne
9/ZxQ/eVr8vjyw+ButtNW+moLriCCKd2dgo4HZHkwap138ft3azWvUl52coBmD3EIlla46LI8PSw
BrHn5jqhQQcdY4Z7zjuw5FAk1cmDFFSzI3DS0XqUl0VNdWbTfXkPAofGeTuCLiA5RW6r+MqspdxZ
4IDYxnTPuhwHkd3B3fOLgpcqlB62LLnmSBv7fKTEO2dzr5wAUdOlQu32H00MQpfnd02H5rXML9cz
QlROvFrkg4qFtXrnRpsFlHn+BCGZHlwpqQdP1yDKtem3nys4dSI2yVfzr9JMWguHpc3fSQ3eF7Ut
s4lD1vNbH3kwlZcEsRYE1spASo4G9jlBpZnKjSqbZJcJHa/+XWaHeriaio4MAXHoIZouRvMAFamG
RCWWF8xLcEn2yQuuISR2/dNoo4Tly4Ltzyw7GvPj/oO7mcRO3GggHHI8adeDqR40cbHAr6P0u4H3
tUWKscMw44tcYwnaWF8kqc28zPerzaTtzGTTpWN+IdR6UOKoKGYhYU/2mH6HX4p/1yOP4tGIVEkc
gAhF+He30Z/sp1W0AEua05wWbWG7vnttap1tR5mLoVHjg+EEMkCsqAAHlm8VXU/jMdoi/jhj83g+
yIZdeypy6Md5iiySGuA7baZC9R3vJjRqOHmZXsW0nrgb9D1XwfJzMq4mGFjuXkrcF+fLU7YByIcR
a6kSD/rqMEM/bHCi+hZWgxSNQM5yUQ6KDpadYgUa2c3asYXl4cFCgr4WC38b+HGxRnsQD6SnY7AG
F85T7XxnPp/uySnTkZzrx2fKnmZnBsxPCO7moSyH15nXtWdqCVtOGf8TGnLF+qXPHUTTbzBcSfni
Kk5BzSd+KTYNOueGE81JGAL6apxfSX29mjxCjwOZG38Ndd3jTe6HMyqp4kM3bma61sYtupvdNQm/
QgeKbygrgwYPYVWEvt7XQCuNJoFj0KmUr8ntw+VbE6wB6+kockZQnzTLexRcOe++Bd2EVLfOICSt
BMvDSz8tvOeZk3DxmCVrC1W98eNHwsX0jBue00upT3lfbRvGNG6/8yVmhGvbh8aW1Rag+DpyPhfB
HbWaRyOdrEWH5ausUrsjHr0iYRnlrGoF4gURgYs/YYetLACjxYloVuElV10l2MGnAFrvkB9P+0K2
CkFZ8ps3Y/GZRE931Zy2mTGpDVMhRLjJBVGlxnfyjheKtQt/irVjWrpYxxb4E4gd38pcNSQh+RCU
6x7/Fm8IemqNo+1EhTqh41i/1RlSekUXYpK4IvcZiCdjiY+XoVSK1il1yiJDlrW5411Ia11AeqoE
k2okVslNY4wFb6lkfrqhNkzF3SGqHAdp5sYCsB/mdiHN3VYUMjzTc9U19D1VTJmC4bF4o0PdOpkX
moymqKOt2bsXQ0MyKyMTnccxW80BfkgBLYpPl4zwQ3Z+dN+5L/MxIOIHEIympUG/69yyAgClknd7
jdlRcuhgLBJkRLycsAll/jXzLEin4uQIWFr2DtbcyIZkFEGINcAx4BA0kUBMlEJuWligTLzy+ftf
HhH6bqU7lFbXK0Qmjbn2oV4VQb9JhxCwkTmpz6iglRkXJFNtjmq8OxOGALP98rYreXzLcVZf1zz5
jKbsbX8g+sFlXUEqJzNyKvYLqFJ+dOqrgIqVt7nYKZ24sELSWSS2M9T4f6Uw7/9v4rnXMI+dfTlO
i2FyFBG52fD0Z03Uv5ABzp6u7ep2pp/7x4gClow9M1ScYF7d0EcEo4vqFtUvOtCejJguQgkvL367
FfzAajoLhfd/9/6rp2eFWttpVJpNRL9YJIpuW84iWciEQqc1hq8aXKksp9afJw/O6YgeGwISy/tx
ORIQfsSV065AheUnsL9Vj55EMlnpurgf6jzCkAbAFs5/rz7yab9NzQB0ER8lMGe7cAVtvDCvZ61Q
LYLiCLMN6wXhlr862QXif4XxPQqlGMhI4YM3O59owirrLbpRN5tMYl7ahZ0kqMNK3k48SwtIcGIj
nJhbQOcQn9DE6Ma5ExX9JCXdSZ7yOa0Ii8MNwu2l3rjx9wFX0q4RL+4xibKRUFvehnNvJsLb00aX
0nWQrDEX5LgU3zPPTQq0Dqg8WxElEQ+e+BtBR4K2QBwW0rw7Nv9SxY9GnODeDuFlTMhrwqw285di
2/6g9BxbJIExxhPYR/AKfh0GVmaHh+n594Koavmlr1tf5PcKRnxDiHSOWvSrmKMdFqbY8PNz/hAs
o7jcQ43Xa2fFlzMD1tBMUJCXVY1BREiHPjVrELHOyF9LINzTa/b7pyX0uZnlJZ0vtdTkaFOnRSww
Mi1EAyOkLGa/4nPvK9W8v3gbOHSb8P9XB/cpPSjKvAxE490zzYoYJtxr2wyWG9Rz7LbqFtowfZqk
9ubPuUcykqDJWeQ0kPCHiHSOmVqQ9R+gKVZt2yx6bBUEy8D0TUJY9TrckJLKAuOcnXRlhAf1f9/E
4zovMt8bgdDpHD7ywScKTQ8c9rOlG3L7q7n7P4RVOY9ckyGNnC5kooftXeoro2R7yVeLgCdFjEv2
lWe4lAOkNYHjwp/Ll8pF1ZDAkdmyJjfVG/y4ftOmpIgd312qDutr/r0r1xniZ9ohkSZlO5CzC3bU
O2ZXgxRICHgBqGpk2Gwqu7PCPReXwCvTCRbYUVxl1Bpmc71+x018Q5rj06Ceea5FxAIUOhrjueoB
E5w6XkaDfkwQX3ghbJ/Qckwv1BdvypY6kKIv8ybOO9ouBzwTgW6UKO9LxwdVeA0hiidx5FvjNCVA
lgI5Pjy5yDrRCRNtUqluCKfh06QksR+RwaoSfhvkRIZqOj+1lVY4GGmti5q61+FRfKIT7Pg3Bt7W
gjWWf7klkwHSHJVkC4XjOd8HNIrzwKlStu8bqrzqP39DZ+Q8wt9RIHjX3NXiBHRaxwmfN9CPqagp
6ytYprP+69rqS+VbzSUCLWhvkzYi4M0fuuhWi4R6kohbCp4Bt1B8li0RxBcHNg9B6x7fDb684yQ1
cY4O+glHho9urNj95GtejnyKYDeCpOYnXA7vHtcZM5SvOq+7e4Ark4E2bSYYdLox2JJJlXH/kO3v
+gX1xPFGt4/2OSlihXsIn6uTNqFoAXMijBppPw75crrIlv9ejNLo9/3phXcAg59rqu13iI50tk34
xfqX8PsV8AyPq6phiRYTHxWiRap51SNqOEqDFiLljb9HpB2SVQE53ad3AXunpIXvYws23bTNlACO
rq6Sf2zF5gT2LUoAM5uCvbV1MRpda7lOwnOhuOlSc3q4536hxVxUzHs6yBIhb5KzKdcLINuCQULt
N/Q6M79PM/NM2e3PIgCV+EacgUOpfZswUQlrqL6sDlPajtyHqrvVoR4YNgk1ClHuzgwsc+GiN5z4
iLSdNctxa7tgPIW/H1Wbsp0PNzIQuQa4c18gN7r5BNlp7ROq4un8Xz2RwcK7G10tSlfuk3bFfF1n
E5Rzf080CCqhaQhyh/CnTXOlfLxk6K8UP+66cYckvtWwS7HztNOrujgeJQHVEuBHAzdy2KyEoyFu
TiQODhqy/slz2me3Sfpgh+cNlscMEQPVSdb9ct+iCEvO+N/lmxIoUwPQxlIwWRvN3zRtv6mXxarr
TEoZiNzXdy02NEGqTHqQnoXu8u8jqDAyhvoXr/WP9tgpET04dVnwP9NoDjCHE0nZcFqsonAtuLnd
i0dpk8GGdReYVW0ZX36N5P8R4QLwyEa5VT8CGTNNtzP4at7GR6sCroE4N7B9wTTHG68DJR/SLsAu
TARQ/QG2TYC5AOtBPq+jmLuq52I2I29pkdRMRN9Vz1oaXwbQR6iC3UvSrBmg+V60mmiUB3eVSHAy
4Kly2pi8mR7qx8r+rE5SSCcg9c5CZ9tmru3nV0CeUIxb+9hBu8rAekplsaCkGvXaoNjrSYt02d6/
Q4O/wAZH36SecYQI8zTPJOFS7hDFvaYfEAGgVaM+irE6GDDOTojfCq5B62jA5d3lfTnF3u7b+R+O
mXsDg+zTXO8OcbA0Bb34uZ/KLN4GBXziaMsHMe8uyD2D7MAv6BMtDnvY9fwBxp2wt+hu/Vz7qUYl
gsCh3JlmHiiOzz32dFqDumgbzrmm6Bho4BsEd3EHpa8H5MPziArxHaxcX5DH2256D8tui5s40V7l
jgf0qMb14wFwXzNvstLmll0uQNiaF5z1C2sfxWSJUA/bNyXbxXoIa/elKu90n6GOv8qNG458mzNc
El06sG2ko3GWlPf/KOtY1DIx5NtrGVNMsL7MNZvXeI/l7T2TjSNVXxFmUm/0hEPiziqBSXuscc3z
CrlorK8vpwMYe1hlW3kW5Ua6Zc9zxgGxPACZQozoTVDjyqho7se/UdXc1MiEXWSnx6iWoTVzksf0
KYFecg1zR3zZB7anZcMR6sqMnaqHZwUWWm/+H4w/+resZ7DeAlwCJwjf/P4XZIL2PpUTx5yHwfxg
dxiqVZ9uFcPskhJ+ACltowLiAXsMU2rwlVO7r0j8dRX1ZF352rxwczfoOwMaG5ooSjFgpLmpEH5X
yz5eQoeC9KjaLwGlAaUvhOka6s/1wMZsOzNye7r72BatesmL44DGxdDI6NcDDgIZzQ+6RKzFy2nW
6cen06QYa3yULx/HTEbQeHDG1WEkzx+EDSIhspzoJ0SDHW+9jm31AdR3lWD2vutxoA2tZyUi3blO
HQi+Q7MTjJtiYSy9v+TkMkMNcUVhAEbbm61cmyZWzuRnpKu+KxprvmP5/n4Tfndg5F379akUfkQd
P3FwY+A2opy7lu1ddiFazEozcrTS0JBi07OZUi+t60TvQ8Mg2d4LViWlWznW80CY/sXrVeqkzK4z
cht542hBu87mgISw6br17PcTgkQkJ8afhK+1IgIBjsPE5alLpLBFCoYAS72BVX0nl5Sj9yXQUXEk
cCV5YS0HBK0NDb/BCdGics/hhHbmzRrlY1UwtmIpvdojKB8/F34qmTOHhkFu6UjJiaDjMONn5IOn
yINAZRqnzCICzz6vhGdsUCvMaMRzuB/x6/lNMN0Cxkfox+lk/z5LbqWzCzSUav/rY5Tc60/nbvn7
/w3HSssdnofGQo3zC/PGziyq0GVa4N2OhSyRn5M5OXuudF1hjsquRNXBMJLMhJhLt2LvQt4LgX2P
ZMcITtDMBGQof9LX81rbXMnp7dGGvMLyxcize0I8i18Jn0IO/YVkZoGmRPfxluEYn5g22SUiIqXo
ME2AmWYHfWV0nezIa4e5q61u0mNDNGUdATJjjq4JJj6wHtAfeOpECusH5GNg2nbTU4Kd3QwwXAjJ
JeY3pBqyv9+dk/pqVIR7GDV3gkv3YszfodfCWoT4uZRKxFGzbG/Y1aYOuiRU3xflIuqBh5/wUvVm
CJ502Ce1P4x+6MiAi0i/7oOxmEoXPxF9TXF0igYBYsP8rh/IiThw2MID8KcvmrqiXDN+RfNt1Y66
SVslMgSx+u+/EoWlt4Rv3N/weKeh8Mx9HJonDjmrq74Xxgh+f7GFhc/AzgEKML1o7sL0gdzWB6dc
xlIbhCe+kJQUfxipwbcIlEiSXYBjALknJXWLdDoC0DoMd3ePP8MEQilnLr0UP0IEibg4MB9umzvU
u8nSM7UFknNiNjVR8U1RNR22oHUEaysmftbGaiYmeWxSU8sX8vx/YBGa1B5Cu1Cizrsa145rB6co
C+ITyCNbGjjFe4MOuGwDTykwsme79C9IyXDKC3M+5kya4pWIipuFYh2zeHs12r/SsKhA6D0tbZI4
MLCgVw7lI9KlRQFWfH353zt361JJraalgTL9oPJ+CCK/sWrs8G9rljbe8oMSGwaCNWD+Cku104mP
WlSj1PYmtDnUUFwi5rdXnHJFJ/jAwfXlO3bDScrTaeVRvXL7bGqBHR1JJzOXKrX+J+vj/QipdUiH
XVrxZi77PjLTW+ttlbp2sAQWGmFAFTeOrZi1M8SU5jqItnEI3hSuBplt8kq5o1ds4vMCcEBQXY+D
SYlv8NcjRurk0MMxUEmARacbaQ5yypjY6c6rVNrxFcWyHIp9TCkQxOpSuWwDLrtjZnCxvEQhaVx/
kw4itD+ArfetbiHvA3Holle46Rlb0zzVxVBPaWl+d06Gx8tTTRov+85c8GKGnppoPiyQMXhJZIaG
lWHw1GXijHH3DT9ylD/UBoHWayF7jnZVmijpkTLYOO1M24H+HRbSDquS64yvo5+kwY/ocESrcjfP
inEFWspcaUyXQxypWmesRhBHJQ29kuybO/Q1eAlOgRE7jBeaSA0fnrB9alAWdfga1jLhXThJ59+0
A/u5TgusAzg5WRqcoi5mVP0/OpK4b4xiK9CsaHL9an/b1l4wkRtg2/sHPAwbhlAHFxe1CkgGdwz6
vVQ3wGi7pSJn63S4Fi58agll6Ae2C1kve6DyWViwdcIXVQpf49//fhyWo8BD286sBVvkCeA0WsGw
C8lJQlN7J9Zz1UGCfpw4eVrnzG+560liPMixSea9sQj9du+LOwEuKYs4ThFZ/VK4fg1ncQmreBmC
hGuJkFJVMoukcg0W0rsLeojsOq4VkiqPN8ES0kelWxfiQywiEC3jTPopj+6ZBzySupr84wGqt6oo
V7mvGZptYPK63lN5qlh1au90POIerf8fFnN5pd1T/+Loh3MV6utaw+WQO47GrklOef0DsIfocInD
JU3y2JrBIPoZOccpisnBe0D3r107YsBbZUXdtCoTMq+Nl32nZrTS0y/AuVbqm9iNT5QNfcgvj5uS
cZksVH0tpmq8tP8lUMk9mime9LLHKaoS5QOxToF1Z5vf2AK1+kvPGXIji0MlEqnYrDaRBUqsXYUp
trwH6Tbbszuu2RTa1FC+Nkwvt/uCgtUrIxsakMCPjatJdaQIuzpDEtH2VC3COZPUcLrGxonchq4Q
dHFu7JUe85wlL6W97bmI+Geaz1CrBmorAeBCkyAPkT0rQzecLmhuKbxIQe83KE9SGA4vQlPGLmBB
p29xyn35DCcD8fRkE8QGHu1J5O6WerskxqkUVRnMortgosqb4PIr4zHhf2GeOLKL3yMlrR0TBp4P
ILdqg1deVDzZyv3s/+Nf0WrKIZzLMNnkju+OHUqcTOXu65gcr5QhUISMycWeS1zA0CUWBIcxUEV/
WZOXyhOr2ldzO5Pzr+BsEbnhbddJu0lrVKkROJRR9IUSt2/trx32j/sA86oWj1oTt4jDx9UH4bK5
yPfJt48SiaKQc4qtxmq4Iql/tJHo3ZUZLoet1fsO348QtMyFhbNnqTeFmkSSof6mfqvExhzZIWP6
GJflqCoOmZHCizfHLnWuQaEabmUbsu+wvysWn0qX9Fwb/FzZuGfkzZGo+DGUGXx8LcahoTIbeepG
XTzQBwBjNJmkHFipI2zPIyxgboB4JBE6vHBvm8ne4YQAPnUeM5fe5qIsEmKkOOxO9NdNR3IoPaZo
P9u/cbiO7ST7D+GfLkUy1hty8qWIJA9AyTnhhHI9pREwh/1r50KQEONsBP1DtvOjSVI5D5jaWV1O
o211S9vkkpFK1En+l5LBxqGLck8Gp5V+sGcOxjcoNnK2axQ0saQRmhQSQolLZjJTnRejYGkub9Rt
ByL/G/oD+UKBIT4Iag5dp8PHS5Zb8A0/LQW8rnX89hi7tEKu4wqCoBqcgcxnv82zJPMbF9RbLh2j
NNmzSXfwXfcg6cEtG5ViZXk+LOdPCd3Mu63/yesgBuXY7xf9QSZEWlWJfVmazi2l6V6RagCi6E9Q
EaMr+PkYkX6z3kN8TlN1n8T3cWzuX96TIZYrh+KS0R1OPvD3nXrkTBELKJGzPuRcegTSq5bUxUUK
KW9typxq0utqQKlad8a1RFiR8a8oU9tUTHs7OJfBLTDYNoqLdw2/JwuYz1G9ybbgGgISO1Q3tkvL
CoHNvF3n9fH6c1L3l3a8NkCrDX7TzPKD48/7eZPZ8HFZoC2+M44qnJCGgbR8cw7SGzNXi1F2XJ4g
I7lu16p/QTrHhnfugRfM7NPVlqQ3K0hhTX5zwtfa17jzx9tv3jFpkxLJsE/3aL7t0tkAy1u+jS/h
a4cHiB7CR3o1/9EArKpSbvOWF8bVo+aywLdn/nOfUYOqks8gzTAg8tCQX9+/AMuBohacBEsa3bnf
Wf+UQocuaYe8qcB87pDEjjgTKmzn+uUt8Y+nkDW/XVJo5jXBYzX+N1I/Y8K4jtyfq6KQnHIZRcMe
jbFFym9c/qj0DtN6A5z63V1a4OzzXdq4gIcO0GNUuOUu1A2RW/LVi2cSJYAQG8VRxtIXuuJdqva/
Ki300HmmMFW0fip3Pe2kWoMqop2w3gkjzAP0ExhNshbUQLO2AVLQLnYcBjyk8cpngfUGLhwPWo5/
I/dcl5eIP0JxyU7e9T6r94H0J5yCmUjqly2mmnN/gvoO58kjIIdOX8nXxpqJ0/MDt/cfE9yhDvK/
YqCyR4WPBP5Q4EHKEyyAaubEMc3IyNUoF+2T3/qLC5LUh7GTjYGs5Tn8/Ydv6DQLfasbDd9F6//E
lcMwYlWFd5IZZPtCzy/cgDk2BtVoXGlXo6h55yTIm98X1ID3Zlzo5qV5qLWUwp5kvAazacv91I5V
+LyNEoF3/kppMfWyuIEAV9ZqyUQa73wpHk1zWFTn7Z0wnu1W0lmpa09omKxESCzixl3+GQukHmJG
U0OOmH87xNBfMzkYVYGowQpU4Mee2CBKvgkIE+oOfyMHdTwjp7Dht8XaYWafy519IwEiiz5mSyiy
zvHp6Gysaxumg4h7fyva6NmqH1/+berFpKYJ94Cp91NAUiomeHTsV9V58m0uyIwwX80v6Usrr3cz
1zajgkPdiVmrdLUI26XXkKIZJA3EQcRi9oANN3awxYj7LIJ/BUF+MlQVCpfR/klqHUtxx2O+we8E
ulYI4E1iDiYenKEV7OVxi9QEfmQHd44xBuE+sA/6E6WEOCEvb8sYmDyiO8d+6siJpc4hKW4iJ1sw
R5FglJhxvwbhjgsYVwZsBkcrl72u55kdnP0lw98YPQM7GIWFdKTVfe6Ius7NTVcZ9ImhwUAi9mRC
/kwwF7xXgSyBqRelQnh2Xj8vt3rem7zGM5zwemdjBa9pVgBNh/YPA75nzNCVUeLXufrZYWTA0y76
Od9eEMRVX1Z1bb0LwIpNMX3NapuMXFzsIK2ZZPrxIZeLVtTmF79PcmKMfMnICcH6piPDnmn3UZsT
+jIWaqpZqawiG1cMRhW6dYrF4S1mQadr75jMQSBAj7Z7+wEUL10OxlB2gN6bQBY+1Uey+FHh2+Dz
Oo5fZAwSGaip7QAUzSPhX8afhO4Q0ZzTrKYZedRJS8Wkv897RMhKzb8t7jhpOm3DkfUnbeH4o+cV
7Vc8OLiQF74q/vI6VG3RD9+bL70fZ5LiyWsnBRBLvvaYdyFYtq/VSRmqWffipx2M3jDl0wK4JPHp
1z4DPewD4IfQdPxb0piq9af/Bg+KCtwnwmmqhcEFVQOLFeS9Fs0OxiU8k0j71ah3eYnGm6dCBaXD
pSkwpC9Ub1c1gWZcXIx8dq1OsT+XSHtzFBkpCsEgq5Kns1HbJKwkiKrLUo8NRGfK3fWovG1iqakc
gYbjYlbbL6cDsQrlUFqry2g40IwYPqnWHuOOtHvlpNwRp+u8os9Ts3/HM4MqZOKqamz2sf4ZNl5R
ONgxvFxYJ6eOuTnW1Q8P6abb6bABOYsKBI27iIEbY+eeGJNWoy2hIfUH5a+ysqA8EsuNNQ7LhGRa
XybT8rguMlHRBUjek3xcrtOgH5VtM8uLICZmft9+due92AValD0pXTzMB03TMQdQKKqRsIqHIske
QX15q5+92KFbY9Sn1FxWViV5LPCfd8ScFN2cvGH9YkjCoyHUDYh9t5t6H7oGcsXptRWzIY0Fr7ji
0fq56U1L848NlCteX9OXRdWoD0WDqp/VITG9jlw8KKVkY4w9HrxWBeNlVjQ73q1ACZqBDZjt7HnF
VD+euJYl81wt6psBoyuyBbFPUcaM3Tj5/X73k1FHV7v8Uf5b9JuIjTo59UAkf1igDjqUCPDdZHvu
MFAsUB66fgmR5ZjOPlhiyYn5PxrICwMdQSJSSuAbEIqZsLIzPLGATQvuvobYJJQrK+UGNXCIM1WU
OtR4JINS2UNTAoWY0n5IItJ96F5eA7Gqfl/yhlA1FlMjTC2CXO0h85zOtj1TOJxhlkppeyxry6SC
JKUai9FicoGokmGYPaE1lMYAekk4mY9zr1LUSL9QnG2GA8v/Lwd2AXJZhLzdOVLfLIKLs4Mxb7+G
MVaHkp7PeuDb81Ksk4NDozyMES2ugW+MTk4+0F0gKOQwbuGEm6TQZiqNSaURKyrFPmZzoMCI2g6H
lIpuO2dJaUnpGyRv25fbfY9IJz146XHyji6Dlyc9y8HjFZI9eSZSkp4QaLYeDqg4wJKphevTSqKq
YbyBgbbybF6dN3nilV4h+9ThiwC4AjM/DzVF2645sPKIBt75bgrRck5AEyn1oMLHYdLD/AarEo8e
frtuvEPb+VEOnjGzs4WcBJ6CJHQQutLIqJe8tK+miz34wr1VBl5jXqtVGTsQ68oCJNMnwvcp9FTw
fWR7L1ZySINkhT6uE5zVPdpp05z8QXKFnMTII3Xc0K+pUC0nkbVSBjHGXAQ8bXF/0GDqWyWUQdBl
007wLDV21vR6BifEbzLXAnT7nK8vgjMEueJ6R6HjEteCXOJskWjgTmiGOHoj+KViQcfC9ogKM1J9
rPuFRVqXDGmqk4vA0XANh5Ee8y2yIeKqxp+2elP0XVdv0RiQkxOLtaBujsKthGPQa7wK1cgiaTlP
711R+aRNt0C8bLlxZDJ8ra/LKVMoOZwaqCZGsDNOgWbyDUiOnGCChcOc6pMS0MfYnCQuPlaht9TK
FmwfrjN8tf60iL9AEQB2IWVtvgAp/BxJdvdh2O7YeWSkUBeb0/s3M4DEUMS+zc86U/vrso9KMCtB
MinC0BhWk4X4ShDjjxTFwsQB2yfwqsd9MvKhgKIfsau84yyzGP208hyQgNaE+brlES6DR6asKE+p
jZ3lco0TpbbnPqS3m1imrqYxRE5ZaupkRoW0rH8YSOqib2UxZILCptpnG/tUOXp8HfpcdbfeCa/S
C17QzguXicNz6imrCuZ//2DPwKNgeRX4GqDAbGNwXZRcTWS9+C3+nyW4EtyQC1veP14tzwukl8kN
V8hB0seAK0VEx3bu9GChT/o8wh5l0EcQIK5pAR+0XsYinRqD5iwoyp8xybiev7HpXlSCRusrsiBw
RrpAd75iyqRHj8wAFLqUpwzxziiFyTIxzWgXoEtrf90RvjQwZHGpHdwjmRSiiQbtwEtKh5Uy0ATv
SiU6CRZFYouXVl8H2xp9HHufO1nyDOxfHP2+Pg2FtubWoYScO7f6dSz/VFp0WZuchLQRoI9gWb2Z
3oPaELa3bpow7+T4GT908z2VsuXr/5T1Y8POzfMKyfMIDpZ73nEW2cHXaPrqM7MRzjmHIuzFc2qU
OXeVn72bLtzS+vFpnZOnMbDk6R+vN3SXCorYG2XO7yZNUlnZsNA6RajkH8rvZPuhDgcqcxdyXyIo
6zThs69VpgiDFhrmUaFTEcmYKtmSW6e43jDOJrJsEmXJzln4JsYEVEZMQsVU7OFvKnZyN2nGolI/
ihZ5KcjALULHIFzencA3Adoh6w1c52rRhQw4tbOc2VvDekuR7D1wnnpUj+K4BD1DU1Bv0y6MzJ8L
OxZGHCKXXL05b/LNng54RVuGMV0utRB/z5qiijIqkyQjnXlFR13yE6eYZS5ZvjlKkjpQq8DQTmtX
Msbu3OH6s23s17jK0tFCnLIZkFeYLE7hXdmCHRgr7JP1wTi+P3FHJ0LyoJemFAqnMwqHMtVqzavm
ozwwiD+dz79EIwBtLfLFIHmcxpPmxPsxGnD+HxGN5wZiMmmKh9GJoNT0DqKYgIabciQKNSMczvwd
3ZskwKWkNbeBjPommcuZDZrDNetc4bItciRtBXN4ziiCL6YsrKBT65JuSQnOSchQVwjX6mTwHlJW
WJgk8d8w4c3DJD59GlE8ER0z5+0sRDyzdJtDI/+Jl95lz9Yj0g3SzRnXGuF7soMF/XieMuEG2SpJ
qlgGJ/u71HhKispJ34o8OmWBv3z2Z84TjLg/lbaC7hDX9XP1HFo5AYIrAS0BUKd8EyQ9b+n7Gp6U
7bzVO3h/l2u5MWDYv2RSfuD/X42ibavthql/w1XFUtraVWNSEXO1O0dbLY2gqgMWEJ7a3Q4anVCJ
2UptB1G+2NPuatXeczjXXkc9rLH6MkVk28ovP4ilC6+ikyr8DqyrQ00+J9oMFZ0tNR+6Rn84u/az
xVH8lbjTdVSETnhVqGupRMMxBGQHvaOKTjW+wu1cy3/nUkgAnnAowi9HV603umtlThipBoX9bvjG
TZLbp3+/vmusE6Pw896gBB36pRhMCRatEpNMqHSvb4qpBO7/MGz2Tdgpk1RzqOPQdASxg2QWR0IN
gB3LLqhwHKz6rD8oSJm1f7lPV61BpMpdVPnDExEyMNydCJcm2Vgabr0DdC1IP45zhh6JctG0L+oO
fVJyP6F/06OxLXBaSH3Vx7KXVol5gA7kCuyzSeMn+1JeDKWvSsWqssMFl22wi3gWPjiQ7r6mPyJY
ChY7S1FjuMVbDKZDGQ9i3s4Bmc5+wt2yVSfdfBUQtQ9F2F+yO7+muj1rXZ34AlcSZDKNSD7YOiNC
4rep1yQB5FypylYd2I7K68PB4Kh8nsajv4B8vNpLl9pkllnNUjDqwdCXKMWDFL9KQpfy0k5am+p9
rFbPPejZh7C8ToLphCFJJ8XTul2w8udDZ+Zteqc3RjzopeUNrT+gHJ9LqmEh4zkvxkMB6bnc6EbO
5k+SExUPA7bXmmQO17dUnQBV/2DVSd1gVnpaVR/GG+2QvCWXTat/umWsjs9y2KRtkpamBGfpaF1a
dhMAZjairBuE/0b7mYMxLIvuPRSKk5rP6WnEOCgd37jKgEtbBDFye88Bx0nSzM3zuKywez6PVy74
iQkZFKXslxHjLM15BT2ILskfUSGLvZTJdks/0C08+yHO10px4RGMtjDORJz3xX8sp9acIzYY0czn
RyNoR7OZvgwESirmV16sM9xkkKJFBg41otKQLeCUt9g67SXDXhfyQCQrt5fzPQ3PMKrRflkZTtjP
ZuGFqz4DLjc5ct569XZWGUPzG+d7zyZLn6QZ3uvjYHnLeEi9NPgzBHpus25KhKSaS6+evMwm6b5/
WCVAP+TF73AOWi3437yFuR2DHTP1uqcVyhKbOXLgVpfUV+rQPNycyzUV5eBIEsmvzRY0XWvYwPyR
XqPYf863ECafRk2ph/tSchwH1bwxkmDAAjU6lfMByzwTKx3fGmVEZ84Ysez926swiilsjcW2n5av
2F4S015I3FZ1vSUbcwdxelhOB09RqOQMU4u/VYGpCDo9kQwPdKzVFdNxLs7vWxo+OxkYfnrDGzPD
OQqaFwlV8X0pC98Vub6vg0MFph05ivzLx9ufGP7IOvW/pS1ZJYHHQpJqPho6bNLuQQICP6dlA9Ov
EzL2lyUXFN3DfmUcZ2plGSDlVY98Hy1r4pK/ZTTRy76sv41ffArpnRIdlxGFo1m1m07JSjy+6E4l
2S1yYGtyfp/PXOopsx8FvBVa7tNwevMgksnvu0ycAyB4ywZPFK40vmIDxx3cEJNxAZuvEGfXG1in
64lwpc+2hZ9kcnxLU6D2YTLILu46LAHpuH6I5gVF7USWG8svcVK+33GbsA9lfmoVLZki7sXJXh75
iRQasFAZfCGwejxUfyLmfIrObj2u3uKHXJfsmfnklLKd5Cr/H/3NZ6aCKZ+qWek09+j7Lktn+0Ml
6ilGOeYd/N7mvv8flLwfBt8dC+mKtc/G/w0IJmXATs238F+Sl/GuRHj4nDRoXS+WL9wMh6/3VZU7
ztCI4Sx0k0FPBKOjD+sL6qngXXjOqL7w0tXKqAFDTX+DygyxhrYWDUzvIx1nDtF2tq3MNyLZzR04
dJ/sd3Yt0UV27WS3kcG518KknYLjz7z22409pB9JWDEQnnPTKf20BGsHCzjIlpTU6hY6q95WWanz
vV0IRyIC+KQMHCML92ZMz/eTnDnQ2nuK7bZaUIw+9SHliThTVUr7b5+f4IReVRTFhds8yB0y0cf7
E2/D6KZGBnskk0tlInnMG9k6Af2LUkI3GUzNISupBzA8SbwZT+j+c8tC+2wA91NL157yLnj4fySM
YEc/Za+Oj7cDTnUJQUQOIofre5jNndpHCUiacAB6rKSok0Xi6i3gzO8VI3MQcnA24FshWat8b+3X
dFXSc9Ws89+gfBGWBQb7hIIx1HmTIQgocZ6g7wKvvWTbEGuNGkYQLG8seRAzeMZnLzQWa+QoAXCN
V6li+By9XSBk4yHyj2yFxqYt0vO6bCbwJnEJeTLgwfCwOaAuIGaEhj834HTuJhGSKesOxAPVuPf0
otImWQzxgB37v3mOSbd603oJirljUQ/PvTXxBIkHOFbRH88IADgxayOozBwH83aTykWiouKs7H4B
zKq7Cj/wCYB6Z9ADPAWbQOLPGBTo7ZSuaaFBpZ0Wr2Qmivleh9lhj9ae9w9ygOh2B47c7TSNRZTX
DcI6LXWYGlnmXriEHDV9jWdLGgkGa+iDHt/oXRgntKyxzBKoxequcZBtaSs4MDPSAP0VJY40AcH3
IQzoTvWOTigNqw9cncWIP4BPjmLJ/pZvCGwtMUBYiVLAYh/D1Elnf5oTMmXeJl56d61uQEJWeA/k
mUfEFiJSkO/RWoGPSsCcxMwbb/98VXKRIyD030Bejt6tMXbqb9QDAIh3IqY3HMzIsLHE1QBSpQ6x
XZDRDycM/D8OuVGYl5QI1w4YXXuSd29HdgFtUIRuxBnePYRXAFxY3FfrB1zJvFeDlNAO4uKCJNkG
7x8FM3996lffXYu7lx4aJxDr51dcR/ik5ptuZz5Bk586rsnt0rE11ZoYSU2No3M5V0sFjMS9qINP
zueV+HTAmIYIkhd9rTeRpaS/v/JEJwQzWVPmjKQ06wn0GjcLTr8n1kZUA3v75dv8qhto4VQFb1iJ
K7OFbf057XGUNvDR2dLypeKRC+A2Rp2JYXAIpovQT0FGMSkRfKLJ+q/rv99xJnYmDHiJUkiFWaiE
xB2ZxjGfiGpzi0Kv30wOfVlAAQJsBh+LWvIGMZj9b/SfPGfJqytba2n/9l9e0KfMk1tVtYXFB7xb
1elTpxV6TAagF7Yu5hphvmMoCWiW3B67eFa43aN8tfC02zL85WuogtVxI2XfqWkmXhuVYwzzgX5R
F9fLYOHS51Ov3Q+5y0qp9weF2Ii6J6ZouEy8lzwx94cot8e2/6b/+4sA37iGSp9YpPTuoV5y5/97
3gypEtCVmnT3qVi1FomrGlcITzmzmSHFScVtnpA1QCAxOF0mgOCXFlW2n+OBFEezp06z76+3Nj16
NcxsUPNjLQaoxTbb6Kdz2XWs/xci54cFGRheQxlxO2uuamlSDIunaJ1z2yjq1vzEV/eJhos9l7C9
nhdt1rqxYhqBBPclqiahqbI0+RWdHlDq05Hkl49ZONYxXVjyeYPAJceo5YzsIDPWGJhrwRXWJfOV
O3X7fptARfr2beXsgHYKXG8R/2taknY8q7nOZZkUPopF5oBJsoFDq4HUwivVwcIZH+TdJ67Hw5xA
DHVaVZr3jSHF/72k4iX4KqESfswWsyXdNT8P6NgJz83tCrmw+sAI20R8FgRpSCkwY6as7JlKuyvZ
EAjaUWIyZz7l6AWZiCrNKm4odJ6PD4S81Zrm2p2/0pqjLynSU4o2BfQPdbY6Pfug2kpXMLMGMoNH
PT2giFg2u7V8K8116Q6egkEuYKCeP877ON2aVqn+YrE6u7K5bgmiAtyX3PXMD4sti79rKs50I7T3
3JkPmArJr8Xs5TKSZDQ4EXUR4vONfwClkjH+76ipDrSbBcfT3Sy5QzAe05T0LOWFiI5qws6h+JMm
0w/vh0/OTqxCWlFCJhV/5jOBTbhqli9DLIhlvshg9JYyJNQHxl7zUoje2VmDet8k0lPcQkDhFhHS
DPIIwGmVnYy40ezS9zmreSJixk1DUGCFYLtLTfB1TMhOksl7mRacyDMKrtgmZfQBP7bqcNEDoGWR
gSaiKL9G2If0fMMMWr62v3njv3PEDWugEh40vy7OdEXZWDwdLwGTquDjINSE+gfsMM00VKoBY12B
Wj7bG3ebbcza/d3qPMkrfG3aUq8Y5lKHuwJjwsVA+SZ5q4Ea7Iy5C45PHeahO6ASAlIuOlaZD2S9
yvoDDY46gseRTL2N0Sof97K/siaURD4bP0dAaiHC3WvcX6JP9mgT5zMt8NXjK/bLvMFQI07twj6Y
p7iL9kDqgiY8oWfBGaVuqBXo+JmbyVBmlC8OU1KuhWExK1IPNRcux0ZlvwZBaulSBKY+HakD3X5d
7lmhGyhenU42XD574fGLXrdhGrR9WSbEjdBzrvuGGmBjUxCvclSl22uMOMflUWlCDy9/ZxXuA4KA
Wl2d9Qd1bhubyWACjL8T4xdOjMR6AHcpka6LGy/zl+m95VpGuq8nXL/qa/lxUl7yxA2lHonW2aDZ
/zTlqzvjkzRHOaWTGOul3UG9UAKf/o50Fn0VJ5DLq/Acx3DsGoYDeMN0RIBQ1iWBCVtMEwN9sxBI
A3OK+gHQ8SGBmFfwvp49RCSokxqECVbBwdTXzQkxiJF8gmX3lpUvz8vUxz4bXfbJM9zSTI9MvPPo
YCSQc6b8I+ysVXhAWsI9pW5KFxMHFWHiH5KewsJIt+33t8jbA8Ubx9PsIwtN/vkIaCsGAFW0V9SW
gP5v91veA6kpIh58ejP/lpvnsYpJefG2b++Qxvbe3JDmDUoaAxJZ+XfCUV+gedZUIkYSHWqQ4RYj
TJ17E0lVIiTW9bkdd8Fh8onUXiILEGHgeRlajkEkH535vi5Pyd/mUIGTYf6hFspJMVdb6ZEPkfP+
1tnyqnDLNGpgwx1m8+8i2TyG3d0xUocO3yW5rvtTRuzd1UQ7ZLTp7nEkF/9W2V6MpNgjyct/YRD/
SDkWOEFA7FpqJqg58kgrzMHinMjiO91LEv6664TAH93hiQjWlF2rZXuuOtq4kRRhLNN2kcIwUoAy
v/JsU+2MmfKID78gdfqNu8gosQmAK8naMfphUQR/Pg2n8nKIIcfYBMWh6W2FaWIe6w9W2O5f4dRm
L8Ys89dJCJqSr7bnrlSoDxwMm0YS7cwseJLrhgD01FD4bZ2YT+5O12nVWHl7XHGByevuR3jnn0wJ
JU5BbNuw+B1Znn0UwoZ0LuX0/gcNR6lO6Pqhnq1jg3fk0v4mkoijwt3nRPdrp2gFVPVRa7eK4rQF
LXPoo2FbJy0IfyMFrCFtSGChPavLni+qxc7okTkGPp/Aah/+L0GBrZZ1XhuUbgzfIY4Z1VDLeZOT
9cLfKGoHTumglD0WUmtBYnD4D/cumQAZCINOPgeog63X+eG6KkkJPyDnSF+7Ix9eOyJ/Ye1LGdjI
AMgeNRyVebyyhVIm4i4G3buXhFLLcVCvTHok31VCk1Mn5WnGPKUawe4hi7s6SxXH/Pv/7XBLuj+N
CWH7X1DhIrJJHJJlwqA/xfxY/Ro0v73OFqiwZmpN/20aTE72e9BXZx/zwNwcxHJnJZaqno/AtDCi
oD48nuytmPLVPYqW0/WFwwbOf4NCO6OgEQz0dlfy2O61dadLzduI9ZsghPI0zDG/SoDsqngE6fhd
61JYhth1ibHI6h2+QeZP+z1ChOZ60Q0szuMy9ClGnGp+7frycC/Qikejn42hyOXqTS+LB9GV5b/O
NA61WQshhavEJhfjf81nVm6WyTjE74zzo1ZtDvdE7ZKgu0jP800bOjVhFu0gGdRXhoclg5kPK3V5
Wtye4/ciHRvjagNfWOr2qzSUh25VINMhiH209kuKfqksIsMgxhYGPzpnR6m/+QvGTAdUr5eCPIRy
/Mq2VcprRiZWUm6hSeA7dnGWIokIXTTUEPUUFlYn4prlMdDJ6dlvL0rcqv5jh+K3842DouZ1rahh
mptdLRhW2m10JIT981w+c0VYICj9hmtohuouRvSs2MkRALGrDSViI+Zww6e+VkbeKEDzTl++Jtzl
29OLA8hYcbeNSrX9nRr0vMvd79GDHqHqFH4ACGfMYe9hoIr4n24SWMDKs5LQ8oe5yud1hBrD/QEY
RvawhLlysA36zfRR/LXyXX0fcSHgmAhFYcNBanF0GMI6F4Rf29wQspCxDA6FqOAFG6LUfJrA7QW7
OkxXOO+bn389+EpLZAViL+JNQ+miOtXNNXiS6OwbiNwVqUCDRh0waymS1ccdynnM4ujY5NpsnNGc
Gwqft14FrRvh2b/r/aNyaKNZ17TeprSGkc531DFw1xgc/knMxpOucSNsj82M0ddA5AR5UXNr8ygf
O/9RR5kh5ipNwsLjNZERPBMvlJ0xAME+BD4HfSfKuRIa+N3t+9PjjAEHiQ8EfkFd1JULxMrC5QFA
dw3p+HsneBAPT9TzwqFJfVQrX9edm2O8DNpsJquEyzrCj2PinTx4N1z0J9OyRigwcw4Tzd/+XXIS
YQlcrTy6tcgWE1rNIyDEAHKmZwkIrtX9dGzVbbYA6jidQ0D6QKZa0my79b/95Aq+3OsZ6Tj80Fvb
d4ozxZN2NUMVC1ZF2g4Ty8EpalHdHh4et2MHJ7QYTlGyp6/NCiK9YSolqbY0CI0G5eJwnbNFgF4F
P8dLQILLgrHx3l3WOwlmJ5FX7XtachEJqMD8Tn39yJkNKwQB1GWiLsRZU5Mppgfm7euQYesd/Adg
OMIMScciPlGRZhYou4xLX7AfxIPo3s5x66d+mIm5P3khoRxtdn8mb/JBB7BHKxLR7LHlzKDfL8IG
hHMjS8X/BplOUiAWHRlDxRYHNAhEb820raKhRjTfA+m3K5tJQ8fX3gXzOluM/iLCcKsS7Gxvz2Uj
pL2C1TGVdpJHCt/7zQE5lIv5MRQ7rm5YVXtapXlb/8eNmVMB9gG8y0SfQsx/AmJQGslmXAvrGexS
UZFH5jtmzISDValQ28negFLXGpB+Ftb4XlG8UQ2Ghyv8pYtjTlQgVLQKXJL6bdtf7YOMPrkZu3AU
4npyu66d63N8s5NjONU0Wl9tppFvAe8ykVMf8tyjC+P2D1iRFur6Xi6SM68eIU/4gHpOj9RCi3nv
UdqntEuYK+uq/z/3eUzSM/Evf9vvPIBDG6Akf/Kyb0OHtfWguCEJqDBVaAFjd3QSzNp6ztdn7Fiw
/eeoz+qiuVXKUyyKATDnCV4QBagyj35UzksL1RbYJNKrbxyzhXLM/bJAIeHOdPO9LsIg504/ytQe
igUByeq3J1dH7OfuVCSjk4s5/tCxtoB5kRjS6MEqSvVSSHTfWDgdSnWm1IRTESuBHRd1PFArpy59
iQqI4j0rYkkOea8r0hq2AKEqWq5VX4oH12kTLAqtJpU3L/5mLuTsN839FQdvGvu5XBbaEwpEXKEq
QDBBD9Fs5JEGCt+VbAH8dI1cZoH7ZeFn21IxLjn1xaVLe8qzMK6Hot8eDgqcGWpo03tr0kTR8Lpq
Q9YuiY6Yvam/4U50deEgG6ryBy2y2fEo6uuVOg5R+CJWLE2GUPU9VYIyxf/zSAjwXV5AurZKbk/i
F9WnvvmqQAUdKPlwbvORrzMEBl0SCyKzJL1I35npGrDH/9bZrFFYzrvNtEpPJwyLLvw5OlJXYmS2
PFP/vT34WiePxOPlxhPWiRzHEfJhpTM1lAlGPwE33koTg8fW8b5CL9VRbfP3kMruzyrF6oulj1xA
92Sne6WP/ZPviMAoVp7ARkFu5M32MYBS2gL+aRs1iF5GRb5NCLFD437Me4DeEr0ZSa8zzLnZ+/xz
KJffbIkvACNEKz4Zbthh8QyeLQdN8vDo8bveC0EZnrZ8vREIrk284zHq8ALnbtnuzNbCGa2pqBrx
O8F+dhk8+tEm9IXxwbqZ/5p3u0asd6zt4VnaSBK/7t4PvK3k5FmHFXkWIm2b5jH4gkkNYbWJuv2C
1ty9JF1PemKNjq/x7KLA0zxC+l55B+jSqgZF0hb4OsL0fi1qNLSgtVgWwvmXPECidlnTZzdokL/T
Ep2IUMEUQorIM6ZLYlvX55r1G8VcuhLRNX3sNKccR0hFppKTTXR05Y4WnnNyfKC4r7huZxVF7N0s
HehQBGQeGXGrVBaJ0cda4/wQftmQuXMpfeWEnObRuQroOW1ZpbyJntsva+4mC4PCzQvDHXnppKcI
wjh7mEoXDkjZbXPykOFTslJGW7d2OSfUH7fOpctj3DAAfHI4bK99bAO8CwOXOn0n83AkYqY16CDj
USnDChda66QNZrqZ8c/vnrnXTHA3joRCi+NNhLDvh7U1aCWI7XJ/cY2SCxDKOrF4oty5SvM8N6eY
yuRwxmK/55I3mKWJTjGRlA7fLi+LhjFtFVygWMS5ISh/V+Fy8ioDJCGvZBwgGLOidX7gNymtlpVY
RzxzTk7tYR13Ir42Sd+ERIjBdR+MqBmU5Nfjt8/3pjnmUi2rD3THQYnHyHTLvN/vV6Vo/zECCuug
TEuP/ajZgz58cax6nw78EC0H9LsmaKZFQ2Mbbul/E5K2UwvI+Mhm7O0B/1taEd6+pk0T1cDzPJBl
N2GBcXUcmmHFwryW3x+tFQk0e1jsZxWXCNWEXoQp1X/gQ5FRNsrWNPSyVscOXP4J8EkVSlM07dMR
V4BR+oYOnY3b3ldsZN9EN6hJ1RCYYmExDstf54eHtikf4JD30oA0Yp1f4zsno8ndV+JTHbt/Rjn9
tXeFfwqpgTv8bnuDDFPOK+xpxnVQdCaoZntCkkJYqsjgtIW6q00Slq8ZBiusR80qVmYVvccz4Wh+
nKzea6n46eTjIbLXjXVBF5jXFNtwqG/DvM5FPS04IGwVzKh1S4wmDW8HTfPZa9oipv+t/KayULJS
7oGK2EO9cJK9SfeUmVBAPK+3AKakD44hD0WfliWsREqYnWI6b2i+ETuhTJVdXQcw6KO8FKdpgAb/
XITe1uYWzos/OWt28Dj+8IWf4fQh429LmyUOYlMiUEmY3ymtHe0gkttipgoegIyIKQfFyx0HfeiI
R+OKs9Yt0mYSI0JH8+P3ksuDO/tKcVJb304bqlRPsv2Md+BZUfdKsVr1pjfhoXAtQpZnMwmVeGwx
ncmdeGUtzgggRa2fUmyNvdtr0IGVNFfVEyaPpBJ+h+jzOOcjVKV7jdWvT93MQwOHSX1XEqiESC00
jAy4PEEqBL2wi0hDLVQXMGWFOF9tLuB413pzulI6Z24UKfYKbK/HdYZ6MWo2D5+5fWus0ZXMa3EW
5m3DrBi4MPkDNLVs7vCTMKIx7zoaL1jjEzPZz0aD1ZFZ8/Nno58UFBaiAasrD/+3/yTSltNzzTbr
JN5eT/6h6ngRDIwyQRZamkH+5gkTWaacw/VXz5VeXRLlaRA0Z1nfO7LfgoPVf04yp5iydeWPgdzm
S6Jn3ZO5XTe1vFZgnZn8czYE/pT0zzQ/TW5xadD+PUiIZvLS7+aHDv+PZq5dgpFPjHT9CNyHAyHd
h8pKcSZUfwxh1XPIk9nuvlJ9JgdWdXmG8+U7Xsy5gpX6JF3RhDscq6QPy5cegfmcbuImi63q57Ap
sF9vGFcSlTheoE9xH3i1oZYzz/kmwZS8XE02vwlbhoS4IOQvv9GiMB1vZo8b8Y2g4sTBnpDo334K
+Wgo06IybTTqEhyCX9IUBqqJcF3zInk4IhO+9VrJX7FTsATL7YBjx+baOVMh/zDPLPGELT95VAd4
IX35oAFL8W8Zd9fFinOw64zaVAk/+eKJzpEO/30KVBUIG7DeV+mx2dBCYArP6vVi8GGm6oguMqG4
PUBjNdpa85XINfRWOAGMyNFYkp5LjdQe8RjeHFHMBY+OaWqVssOceBdY0fCYFnfTTeiGELaLklgO
qPeimpnySOjwx6t18ZPiWNYbCB0vn0YrdfKSr/BAHZvjr9inZ+PA2tVXs2KztDtzhuw3V8/tCTUY
kqFw+cnLvnm3d5XD/PGOitJy0mFn0QaZl7FVL+PjtPh9qm0D+BL6+Ax9fWwbaVgsFl/FWQwexzoy
6rmPuKJfsHni6Pmb2deq/KH58o2ZWqgA45llMqo1xlc2BBHM4gwk9m1PM/ke3vK2AzYGNTDxGL9y
ymrqROdznf9IvKMcXfOBpbs0B846e32yu1Ia3OUZYrp7YUXjepmh0kHKUFBHH3m0aiAnlOiTPX3j
0hZMrrVEOXQMWRmw8fpKOw8Dr8b1F3zPLkuanjfQfSKR0d3RfICPAHAiCah8HUClBTy7mY0c8FV5
ex3eyTtOHjQW6Hf4Wna1Qudyjy3eBzbpB5dK9iiYZXfdk9UZBILeRe85nd2wzoWCBZZ88RPgKQHi
uZl1jg1GpvLZdX53WM2pGpTUEiXkg/XiK/AVT7tKRZafxhmbNrYZW+Tzb0b6UHxNLONdxg6cDZRu
KH/59A/tsMjsT+4HVYXRzK8XSaMejNTA0KKT+U26UYHt5nBjcIHGa+Zqvv+YLc7xswx7ZuVH0J9n
fsw6kabCkTY0M10aZNeIcOd1u4JdmhN6dv2CQgBOW+n7CJwqKjGgzTHqA9lpF8ACxipqLKaFn7AO
rHBNmq0KdeMn8iHa8PbhDbI78/EGJ1WWmozoKNLpf9CMSJNtlW95X90RxqBWwk3bN8BGDGmdWjpZ
EK4AG/OIpEUcSjQzUdLxLNG/dIDajXSeBlOu9HGKFrN8+sr+wQ48il9zfzhaIkEdUiSrYYC+tBle
ZVWoLQIwh3+Jdqcmkru5TKRmYsuynY431u8Cb/cb9nvyxSwNyaCslj2bkJapqAMlVtDbo3qZWgoV
kOJKQ2Af4y49lOC/nAakT2LlcwKTkxMfNAx7v2/5Didw/dNeqBXl8kjAVd6KrEmJ+XLsaTUqYuYz
RjTzbCzknIzsMLCzZ7RtvaFjSSRjl6tHG83nFXTgoGTVfuu++YnFGI3DrRqenEW3DkKD9nmz01te
Ssm8k5sANpYxMQUdf2al262wZgjD5Fs3Zdhb1ARtVAdvDNbo1CBnM7NC6N/gbb7SSyX5HC3Cg2eR
hvHhK5VqWfgDTGV11W0ZyZuhKiYXI0rD473JqC+Ovh5Rg7r2FbMbzBnikH7bjID8cYXCTyQ8gSFF
TazlpzwDjpd7lqw+5GZHNJm4kWB7kAM28JrsFpRrnwHqaujA5CRFDynWctB9+i4U/7GbmQnSU2ku
QhrTu+ez87EQQxUazcfq9EGKXuKurr3LBaV8Tzl4BUVzy9vbGfncXm9WyPf7Dhf7BVsaObizpFk5
o6NP9+QVWLfGTclfFZ0pkaXxf2yYgslZurOe9gdMS83lBRuuBuvTGOyVIsL/P8nZq4BaXHZg0tlT
dWrOgT13uMCNi0nu5lOLOKgzXTBkX3jKoBTerGJ+R9HVqYKwGCYFzfsZ9WjJwtscH3gPeY82GQbT
J3jc69A+JVa9TSfTD0Dql8KH86BClulVX9agtTd62ywjDafOO/I+B6a3qoAtwVsTDIukeK4TKVOV
LT8mflNfKhnbIHxkVJbipnKtjn+9lAj+d9Jr+iPDJumWnv5l6qpiWQ0xwodccxR1+kN2ixvhqB/t
xwqEkix0mMw+NeNa4fGKe/qYu3e1bKjNySgmSMfK7vJXRrs0MIruRmShq1ZO3poqYmNqoEtOmJ3V
2n2YRtZFZva3wY9JOXUf0ciHwfm18Y5nO09SEXIta8y5GAZ9FEi1+puEgkjcthZJwF9/fsekgplf
DTuRsPuAK2Jcawko2h7mMTUi0RtIXy+I/zwQAeKFKlBE0bupEJY1PApmsMV3q92bD07xLxKgGNJH
hc4ulv4pUezDjBHVDzLGBbiwQuOVI4YCS4B59nmAHhPO6/+Oug7BJx9mO6XVxzj4/BsHFPZxf1V0
f/VhoOmR12z/aWql7hrVxNCiZGIprpM3ZiyUFWZ4JgPvSdnrXAaVq0DVJpAsHdc3N0eV3qhA0vGh
XArPftPmND+a4ZgVafwZXOyFzRrz/0wC4CF8okCIYpdRGRVAtBgjYll8DQRPcYYRWWltyMml0XyY
NRnmMzFOBDaOhW9eHaCexOYQOotkEm1AMlPBsi9xnzd204k/I0fnCdFTqCcoAGpVi6rhi0NiqGJz
t9bHIUmRRwsD70TZaSGFWDnzTOM1tDJDn60lRwR+MbFeOZruENB7RPKKtNZ0wW8KNXGY4F8oaNKk
j5AvW5aqjfhkAMUUfjiKPA2MQFSO9AHdLeFy0mpfXT5lsClRcWZ7U1w/s3n8Tjc/PHQVIEu4SJSI
y2MeULYd/Q7sMUm2OCevxBGbOx5aGwh5qu0P8KLIOLMIOEAWZgTQbb/2/VMidOqit8WJGXyWYoq8
cUxLfnpzp6n1Y2WWyTdgj+0atgjsYj5Qt89+8chsad/db0mHY1cvdMO6Lrl9Te75oSm0c1KTHRWw
umfEAMEl/LXd6icdjTQP40s03wzPSs/EpPJsv7YbuHaox8bXh2n5uthWTHg2cKNIBEdH5rKcerrJ
bhG6jIKnw/LwF/cdndap0bd+dk9K2wSwuuegf17Vtgn1qghKDkMIhhw/V13NHMLr4GlmAbLWnK6K
1GA7dRHfDkMNxjw+UzRSdVSeaVa6C8fSQ3Hks5m3KvYcSEiNhj0WrVTM1GM3MOdEKdPGDMTGB9ZM
R2tJ82oONA4BQhvmimdvLraWAKXhEJs5NB7VcLqnmcrfPmK6wee5c93SpogkFENph8lKePLAb/uh
zVVtYNhkHD9b1fj7p8wu9TYr9a4pW9i5EQUEhrqvVZRLq8eNw5O6hRJDMkgh8/tgpAoK7tTFv03k
AmgjOT5dSKKy890oFd7Pt506MhcOJ+5iJJMXWTX1COPGr08xd1oc+U6G/ubsCA68B/aPzk7fsj15
CwwPfIzd/xPZhOA7FtPv7tLve92f50SU5Lxnys6d8jXfgJ2TOj0cUJBpIDEwdDcbX2axa6by4+ip
k1rXAzpgIP+mcL6zzvbK05h1S2h0ax3fbsOFsDMOMSJoZY4oyh69EWtGYUmiWZ9piXaomNMY5Z78
JalA9cbS4BsI3fMm/hSN4PzgGNfBFHr/Aho/qRrjvXStcy8fbElCuQP2lcljMhUx+FCq2tiRRnDv
k87CN6fK9fK6Nh8pwSM+pChf+bzzFrH1zqTI5wYcmNIWm4v441CJNoW1H3Por9wibhER4JxKucel
rrW+AYtI8OjB3++5ETFv/uiM23k+LLRr+NrA3bom1l46LkqQaXoiCL3GwcQzpWBCThNG0/V3+hvj
iPNYw6BlAo2Ay34YUbvZwwWlzXMxhEWhNsTK7gvpjOp7JKzw0UlEF5/57yPPtvCJDreOkBbU58T1
KVC+PMB4Sjm0d7vY7hwXdCNkocl3Sy3E0DA7+GJgRaqlgv0PWCLnRF+CYiGAD2VGaBCfXYiGnRc5
sDFJ928uKm+nPIV4wNWu2uPU8SWTzJi0paWPLRbHDzXZZUjCcTFFbnpbCW+PiL4NFseqbR/7impZ
qIU2dSFNFgMgxBeWoWggtyUyINr6irlpBiy6khxyMWowi0ZrksvUzF7eNlWsBH5ejodRvKfjlmxo
RG7oHxdE4P5W28lSSevT1avrvVBaVmld6ztkk2C+EQfNTKaDwuzRlggS7R61vNamz70qYXztE83w
Korf/6E6YWYpnLywKCBhGJIEAj5V4uYQlcJsJQiWq4aPO1+xz7PJ6jSkAH1GoMOjdWSZUjLHdF5m
JBgOlfi1uVdXVapSGIsHc/gF5nJTlO6ETxV+HVzZeQ/gHmdo3wJ7cPq7ufO4Y0G9yRSdxx5jNGgP
Sl2baF0dUtioyCVASvjuKJCeOW6MoOxahLr5CWCwks/eGwfCQUTGiESyqGfTX7eBmXr4TmtCQJAz
0CXm+xy7zR9g2xHBHyw/EfqTc2vhVPqIpeHtpEtODVF3EYO4YJMptvMWfHKHmlUIThxBbHDeYTwV
7UMh58rPWi8yGCDP1iyY+njx24rbo1vKruQJlIl0i1oBsfKGHs9MTp+16pM5mPHi8MqZi1s08SFu
nf68Ot8i0RhU1ds3IZ6jiXEBBZfcGWfKOeWo5EzcgjsLQQ7vV6+XkyVIXahvQY722OAqrtmwnyrT
8Z+XVSATIG3PfAga2A7AU7CW+IvdDql1U5+WJeec1k+2S8jaMdslSH8vSofSnvJQNLP2HWCBSZ2L
+yv2+DXbaRl7yRILeXbyXm083Esh25m4QMLrBQtg733jCgCOHllOz1jClFPabN6JTQPpQdIu71Sp
ZpQfN97awp5LSyPKK1anND2u2+pINgJXgjoHiIVYMvJchoje/OqQ7B6Ff4Ofp9Ne3fD80+a3RDPE
cocV04Ax+JJu66kVKmmMYEfwKUJ0t6+2zUIDA7YUzpWJk8EL3dHgahNZeSlqW47mdQoBgL8zfq86
/JXL6NrHFhQIjvGXi5/Sbm/6dlcvVw/zkkc4qOewRSpjgPKtUyP+XEjYP1qxA0Fhhn0wYseUSDkv
fqczf9GGRHUsHZnxYP97uAJzkdvp5fQjtKpnYEBwlO6G5frv5IRRUTN6o0hRPsyz9ipEgVyzwWkF
5kM7qKaov2iZprg/BRQFxrZ0byQCQCsJqqQnL01Rzt+9Th7g4ioQRWeoTogcGPSFbAevRFNlpJd2
Pj6ua04tPETN42ISKls1tODY84oNYWfn+6Jt5b0/jIq3OMKxF16HdX0vKI+Gj29G6gJA9cFyCJ6Q
B1BOBO80NULR1KZmyDfqcZYl/FfJfxzgMPLimZblU0Xk38jhGjJyG6e6n9cr2ILd18sQf3IBdWog
/nQgJgZd9uOBGYbJfV+moskq8mYpsMuhL49HNSxa2dWOazQnTH3FgVCk4o5z6F7yiBN+QwwM1QX6
n0BU869uIFBW+MsqRIX2jZV7P2vpFsQMyUj9iaGCDLTvtZasurh2+65vYDUFd9pSzt08grmeuvL9
xKIXxT+uxyk2v8UTuP0kIrnVv5Xtou65fCL8pC1m9LJC66VJQeBKspFrMuQYOOooOiRzKB39JQ2k
7k/CTwZVCwFr3YzMb6yZZljW32h94DOYnO476HW+76jqmCciMSN9ubchsqgg5H9vISvlTZlV0FpR
AClau/pYrIAfXXqSiqLrtqmpzWFLmxF/InftSisLOIvRjvi/ZqBBLdcvHkV+FaEbGOSb2sO+LDYT
lgwOccyYP1uXAR7P1dxhevvbkgBGxC8AstIDUMuKalapplu2yn5baBun9kMHkuB5V8BrBpF4oIdq
TD2rYHG/TCvKw7x6HC9mBzRNcrGMx8MtiGOLPLs9WVWpLCXFCcaUCleMFcfL8MQno5CEBBbYV0qb
hRJ2PFBlBD+h4b3XGcZWNUNeKE7nDt7H2IidiB2M7BvWSRLdsAISMJeqVBuDRe26n7g1bdZBjO/x
ppsyT+yXWd4msrEhDiGHZ3hdYzY/COz58mUcPVi9KEr42HNJ6VxXJ+iZilqFd/JEllabw2H2sGyb
luPmJ5kdxmOLMZfNvOzg26K2pnaaousFBP3coO2KbHMkJkUsDUXwxPaAgxVNhsslHOKLibgQdR2N
PxajvjR4E3udopkpCWLXcy8FNfMlvjh6vjI5k5AjGjwyyu5vhkIQUurftsBEj2Cdab87v7NbJ6X2
5pHx+HzY5TcZEM4GvX11lwSNabFDCaLwYDJSLIpE2qOPgmi33dwmkGwI++xuq45zmGOXawQarD4X
GEBNOjetdHIyD9hLg+biSMRQUy77gm2wino0JOcJao7boZlFmDNzJriPr9izhsnQyyss6MW9wGY5
k7r88zL05kG4cGh4MYimamG2yVFUQsM+u/XzGyl5vmdHMe13oREjNCg2mr2LRMQ8MgKOZ0cj927y
9wOA8mqtqaCWzdaobuoTpY4yH95IldcbMo50XWqCqE0gjYk8ghLlZnZ0//45o2Ls7wIZKFa6KEH1
CHne+BFVaSmh0oepIHh5LhBS1NukK5kNZN/Trwkp08ovxkUDVqrFQtG+6+B3H1o15m3MZ/q7lgGX
jBEmzCds9iZjyls89AY/zeXKvBW009ysAvaT6ysKO6PFxt/aVY2B4kwbuVCS3kuTmxxikGuRRkPg
4JUWwN1PwXzk6mZbjQuetrgCl8cgH6pxX9yqwSq2H+tPdF1/VBoiSTCYT9F9AShXhiYNH/BVbhVV
UiFjrvbApqk1FcbYFqvQeP4tHhwhxxd4ccDauxl3DniZNgTdUO8XuMJdpKGW6lPGxQv8Hb27FOUe
APBhoc/q6KrYJzyFu12wN2CYUGz2uu0dAuT025dRkseNDkFKtB+P9JG/07LfsM1AEP6x9XFGRS3c
nYGfqPB7b7MHBvaW323CHi7z3xMpkLEtunZR/RPXR5EMBW8DM3+dsacNqs7nFO6EV+uP0kfhaUBD
wNA/kDHlzyKWKszbL/qxy6S1QWYEfaOqymptD1JEdxt6tafTglhcrX8PfeB6VTt5RJc1N2Q8tZDz
TEeroCXxFlFkbgO6C4kgS3PE1fe0N+9D0p/fiVlQTAbo2+JZx2xf3pstsuelsWj/FK0PtQzfG46i
QMM73FPlyOhCGaq75OVBVeqUsRbZwhvX6lm2g5sRhmsKUa9+cvGkU0wyFNEAV0oB15L51LNDkj3n
05UUtDwNmpguA6s7YlxaK+2Ac7rWHR9p5f+/oQLJdGRcwrt2xAQdwB13bWeniA0z+OpFCBv/paYT
USIOSEMotxYzALyUINmDrrFtWHQqrQJeT7AhPUDtDYuInRwsPrnDVkBvwb2L0pjAkOee6jiDYtZw
bLWmW7EvNTP0cE7RJ94o+8wBtA0pCYdm7UF5ESoUyHopVVBrkbQbhMUvKwoKW8q7JrSs+Jn6jUOs
9GA5lJC9lJqfdGZkFQYDCuxgIPSTSniXc0ILfM5YSqgZ8GVsXnArYgJ5Co6cOxJa3hRhy3l18PAW
D8wZ/4gjcDDREFq0yKJEh1jV1KVrKt7JIB5MaK2odH7Tw6+/qGSutZ1zaLfsn4V/pcEYQ4IIB4HV
hC3ZnITHjISsrlgdwSo3LSYgcb08n+O9wyVg2N113sRi36/MMFeejQXdoWBCHBuDG41vYWDnZXwh
JG1pp4wQ9kVAyR1t4Y6Pw9fVvyq+mBs1KC4MrP+PcFB40Ol7kC0zyJtSfNDCJr5z4oXHwfZNR3cE
AjbfEvfM9QlVT4tChyNAmhwCE/L+TE/8y0DxtTcN47tntPPT1U533rJGcNDiRc5FWjN7In3s7XO+
1RsZGt2fLoBQ3UWdERdCATz56ikXLLTWLQgYX/Ss3c/7yNlhVcw9mND21FS573U6uD83yH2eBKoo
WP8VRr8jpFGIvlyifGVfwdYBFQ1Fn//wFI/8c9VweOQBrMzawZ3wD/j4WcSmnqWbU25k2M95B8Ot
2yzMXDjGujnG4mg6A80qwsB5aD805m+VFBT+jzY8rIhhfQbeNAHfwe7mZC8neqMd93v2ncg5BJ69
V6idkGYR3aXocpmZYsCUvth8P5x0KwCfFTNOhZjqlmBF60QqdEAQMmLbQuYUWXInnBof0OVrUVxV
rsvKx/nUd/YrAxDfj+liv22oCpvltbGQHbWhEdap0Worn0g06IkpG6I7S6uftqVvd5ooK7vcPl+N
/knrROrt7jwstN/F6/43YcFDPPe7wbky9DZJQEekg2JMfV90gQOFzhCzuzyAbjbRHMr90NsBkL/H
dhfLZc/JR051GZlLrk1oqF0XO+DEOFy8R3N/0wCmtF9FtHEiFOD5rDH6hqxoNrXUnz34oxyyR2Hm
LopMEmU09Zlj5oLApnHXzkBgBWgqf9lXRUj1WChZVU4r/OdgqLVMka3gEOjKElMn/LJHaCcsFVg+
NTJHmeWuBDzNRQXqlL+/fEC9KTOMpszIOoDY4aGqK/2JUKggcJblv0pQC51cVI1QthJPz+ohgfGG
G0Y+JPTgU6mYrhjwf71d6c2zwA2RFYYapQSpLMs5TmWhdzXRaTPnpfokj4evkmR+Nt7Mrd4veHQZ
pvoU6i7zDDhJ3ECAR3X23GdecMYp9KajEbqjy7tBJROXMkpJnLKzeWGZF6MiFAAsNx2JGVgBAqok
h/DpyJNCBXIUHdgFl/vkMQNnA3z381gOaLcLooT1bRs3RCLoVYAZ/h+/m5b9daapN3nvh6rqOgSK
lsfcb377yH8lBmUAHihjy2KI2kOGIehttXXnkjkAbOH6q9TtrA0Dlsb6WFKK5418WKLfDVyu6AT4
9XYPBDtYCubQZfB7FN6+ccXtuLHTGN0g7hWT1+EQSKWz5bPe6PvDQcdwVPMUPUlk1RrM0zQYi1k8
MytvDFD2gDDQ5bNAxe7rYCB4NOT6ruYXD6N03BfegtJqiVzckQMNAIgNFrp5Su0qQljRsFiOG6P1
QyRrSSSclfTg5qO91Y9zs85ZpCE9AuXQVheZb3JowE1YZonrSjp9jCV6ZTiaUzxSraY/fJrzLney
99wrLa2NGYPG/BVsxscp0NYf8eIblPDH7r5tqWAJR+KdCcs7f/1WnST552FqjNglkZLgk+vW4hnF
xrBhiXLacAZgx5GJQQCoSkXvjQtprwwZqZGVTM+jG2PF6Di9fLVtf9Ry4I1UjuJxRjR0+nJYytXi
tN17MhToqidJg0WiGHnBUFqS793YZtGMu1KA15E0hlKic9BW05g7qpZKCj+YEu5sjVW5ei/LM9ab
o3UMb+FAJ9IBKyk9qsQnHLwPmwSL7hEIZK3TGrCdDgnONJojWhk53N+t6Elby98Oo70GfiGnLfum
B8fMKK3McgxKeuzN/LP/wzDUdneiDU5jGCzzLwTqWmXp917Uaog87913ubB5sn20klRZ56YNAFvC
tiJ9DMOH/2oTJ7rLQqHCTlQiRPVA1bWFaFUgSsPQn4sYEB5fgKgBy8dxFLa327de6O0uFDulBSX0
q8geemm9VQh25na/RkCBiG/pnSoaJlFvRhd4hsBP7NFraUQRwXOjjzPIgeXTisRvgm9bz2ezTfod
z9gD/OvCEfbEdnw0ckDx/IGRMDnvclDsjnDVTGD8+b0EevKxlh3V8EFg5OFLxrB2D1ac3t4fzsJA
v4te3rYII33PdPwv3Qbv62NoOt4KT7tsujggVlrl0KWQo3XdTBllrCZTbMMOEqrzILkkmpQr2i6f
EbKj3rFToDzMGDNmjKa/MZK82+LF77thFNdnEObkMBTFKqzfQtDWFIGFtlEEl8n1kgiolU1VGXPf
FBkz5dEQf+UC32MZgRwShItWmOltURbmMjw7sJ0KVo3KNPlkyzNBGJgcX4UIYmzL3Iv4sqBF3PJb
Gkw26t2KVxltutWqK+xsMIYpoUmNi7LshrYu3ry/Jm/4gTv0OkX858y77OmTOJ9Sy4g6Tu6EVZZG
PMsjBFKSb2PPiUCKqHkXJjqRfH2BuFxHYlIxJXKYdbLb4ME56qW1KWBFLxfeMUJ9jnJL1oPiDdca
C1zl1JNmolX+U2UvrqfRUKn8HrtBQNY1geBnteUrv0hkTi2QMFYWfu0MPlGjf9s7Yr/hufPI/hjV
2vmGYcJyZnKKQfWIqJrttVzUOIVsrvNDN+2frmuPSP41SL2h5XbgS3ao5Ie7q5v8kEfcnBydZI50
iwfCT4tv6EgMeKRrCkNRDzVggpVslyRsICB55MCF40+6bqX1iL49UOsF1Qx6POi5mNOIZrzoJFwF
NsKt8FQDugnOsFHjYP3gtgeUnz5zOntdFc673q0nUGX15RAU9mPVvbVUpxKi7OgxYhv+hxaW7u4Q
s01niL3lpuQqPaIMOAVHQ+N143evd0kU7Lk0h4lc9zJYQP+6VQGtGmP0mg0MT8Ur5MjJirYczOuZ
9B0rdZceos86BehP+kivjWHz29Ot1nAoNcy0seB+w6JYcnv4XTSrZILRIxG5yiM4W4uvHXsIqitw
09jqG/Y+PccOLwolc+UmCpmAsJgS8JiKWPxHH86J1ixzvudbc2BTnsyPsIwCpuNoiPZmDsY90H66
wvV5EN38KxchttfATauUztfiOEFUgba2oXG4MupGKCDC4aF1XDUABgIFm21//hQDyJmL7Dj37NBw
+uaG4dGCrTXmpsah7Sdap7lo/xagyCzT6JMNtxjv95uYfw4qN8p2KbMTGOy1Ln5pl3dNsqyJED4Y
sogBPfeFvkGoonhf78/S9F5ZvkxL5wokSIzvJQu1ZDemcRO9KCmffIn3PX5/l5uHg5iarPpvrbKJ
jexuWoxpzcIEnDOzakfsaAooElNJUZL8tpJTD6lprqHTPhvvyu2/5p9FrgM4a0aoPSHRV7H4U2gz
Ti0jkb8n73Zll691iG7oHoKz/8R45BpgdXsgEn3gbaOy43MXiEp3cXKHxLyiwAduozr4C7Set3TD
G+NiH8z1D0LMMaa4dFkm9RlNnKGdEHUH/MB2gNVdlB3D5Fe0DacWLyxDA8ehpgLyQdq+NauAjPZx
FxiR4GqcgxnVszMUc0PHojZ6saibCZRS8jUBkW7fJfPCG+/PwIkI/JWNtD66cnou2JWjIBE8j+9h
nns1QdSPZBC+3oJW7MrHfvaHbknbpY+bdOd8rG/3BBKFFa633v9ZOdz8c8IZ3E990D+Hl7Z67dbp
G9iBxLyHPMR3WGLIWDFnsB19nhOf604wme2yXOnrTCXV1rVIT0pb+ZRktXGXDlMPpQObW3Vup8ud
G1E7Q0duQYxy1+oBaXSNdTatQesKsfe5ZZwp7QhHyXisKN20xoTA4NQWP/j2RWgcsdLwSiVW8CKd
0zyUXtxVaVAL8IV+TFes4u1Ghk20BzaHsXYJP034jwlkUGjw8S2d3q/ejLoxEuvaWfAVem1Qas1G
6zmzvRMKqRRkVzV8v0tmFp5YuEI+AePjHmU66vGIvHcsELX5eknEE5Le6AiCful87dUQoh5uCQ6D
75ViX6HTkxDtGCuYYwrKGhppYr0EWYYr7uSt3YltxvdmGsDu8ePgz9qtbva9ouCv2tIBVsisBgy/
wVPf+gHBPUbr9JfjESiVvXvc7e1YC7+giJdhg6MxNYZg6PM2rrXBdpRJHFXEUl0WP+Hyqm5hCalQ
cFAyaXpIghUck1cI+/j8n8c/+n1ijDk5WVsTOCBdpa961QJLYlgtR8zjYSBl04uKzE9XezC47A4k
1rWQp0R7Rohd9MLggZETm04NsN9mf92VqYGGdGwF8GpDyLbUwz/lwEv9BnCWzVX6Kg4t9muNZsCX
unDj8z8ZtW6bA5NCRNmyCFvyE1ITe/NxXQCpVNeBGx2I8vpXmuMhBUKv+PCxECfnl3PqPai6kSEP
23OK7sVXE3PNI0jjmj0IAtk0aIYh70eHEutZyiEzhk3L8/kM0zCEbdA4bjr4fWrt9JWwSHCNZCZQ
KCcoJeEgMmUpTIPYHhSXEef1ZqPM+FP1mMM9s6s6RVin1NrkrI1xsdSM0yWVf6N8ARBvE71qh44L
e2FmdLwcHHg1zNNwk11AQVZWD7bNSHzcZBKJZZresG4bRip9LyE52bOsJnnNFnPvr+xGSDTVsqbC
HnhAIytsVYle++9CeNjPjHlwdnCk3EqePi7q1JMC3ki4Y3Ne+V5pdU0G23cuto8z1RaBEr0Qihqd
uwTrGeUqegpU8eYSoYm6QA0rwWOjnDMJuyHQrNv4gnHZVoZeaxXCBPyAwpRb+1x6So7A/E39D5SC
0fAfh0d5dytC/DMazwpJ7tgnOL6L/YCAFdNfxiu7QKJw27LUZDeKtCqxjCTx6bTEuwIhwVEFKDfI
KeHTZhDDsCfNq88xBZg6PfwPx5muo0mNJy6860HUnbn03EqEDIoYqWGUQYzEeLvDyz18SDWwt7Hz
ihojY+4DklcXcFRNH5ublcEVqnDcXap1YBeCkvAyEVwxbkqMFF30XkN5Fqkfm8GZzzmM/NiTkBl3
wecT8g8bYmvrRr6gynfX0/2SvRpLvg0IDDJ3pT+4x9Er1vpmTh3gNVEBxHjSIu+sOsc1pICRY99D
qsbBrkpVr08qtQXcr7IOsd/D/7lXyrGUvvYJa+WyQ5oHP4vhfXCbJwShs2De1ZT6WjCyuDhgiEjL
+q5jKW7AzjnLCqSY/z1oRCjsYK1GHrxHurydO/dy0GPTrfGlirsj4DRPv1BSu6eu/izLwLYEq86d
sD/hHS5r2SMruBTHW4x7rjnY+z55wqN7xNQQy1hEn/llWr4GQolaP+NyQDvVlt7ReAi717ijLxEC
Y3Kuh7dSpuUExYNln6EMKXyZzxIIrrSVYE2W2Wlp+Qpy20HIbAlrceduysXcSyeHFH3xKLvs5lHT
ppzsd+y1uwQjABZbtWcoIXit25NOPH4NW3kTDbBiZGkshfrM2rO3K4Z7O2KeWx+s7kHqM/HT250n
GFOX0EN9tX1UXy04kzZpE27JbX4CG7nB8KN0bKXSbMCfa08XZ926v/VEx2so0hisxYsz5KKH1Qh0
RICZkgxtTDkvRH947/Os0zFT5pNZbPifc0t0bm3Mtl3+70xmLFiE2eycY1NsJNGjKOOn/NQ9OYy4
zOnvnwLeqObYIULWheasKbCTP2rRfJ91MWKr1rxYZ6XPmpCliRfMD9U+so8ObG+6jopD8aia9myE
+Ohz5qS5YtLuYVUD7NBJKBt94lS7HoxnV3xou79OJX/2Rk0NH7Gha8+Roo9SY8na1Lf5rSvNi+7r
Im0Pw5h+tR6uOcZTC+CgO5QcAZ4MbN08hWwp8lVChaFSQlXGe1ulT1x18Hm5L4ud2WmPWu/MUqkz
Qx+hIiEN1h5lQC2iwuji6Wwh8iSLwanhRhnqfzTe2rdxMvGezAF7Rwxf0//ABDzGm+/si+cXHJ4g
ltc6+UjVJw2Ob+qmP2N3srFHUtpHUo37BixoPveDw0zRNPrxMZkf6tj1FqqWA/ipWiQ7IP7ihTgj
bV3KGVGw0EmTWK+kTVZoLBvzxtcyzTAPysYt0Oc/x8+4VmCIitrTuWTtZT2wAJYZGU7x38vpwnLG
XunPleZui0OJ80bdtarRsZKQ11aD0I6thewNjQUMSOCcTlj6uwKdVLDWp4MNzGvLvquodAWVPyF6
+CEty5aokFkhvfurNyAx9MirjJmfyqgV67k7HU0S5/en1RwMokUteg83nGc3MPy3gy9j7VzjTQ4b
dXsOwuqHcanVrRYAGB5ggo2UU04MYiLMSt3a3NfZAATwJ5ptCdv5Arjs5kDPeHtZaMjr72XV9Dkz
zV/Qgql0dw6M96gHOY/zKiFOU6sNaLbMBWs0P7yfPagYV95R2Eqf0SRVsw64hivQSgha2ZXLWTMP
5FzjHfctEkNzepxkQb++H3NOLX6QUTN/RKCxu5X0Lgmo+PlqYYE0trTL/FaYIZZ5f6rq+D6Dhr06
v2eMynfh7uSrcOwVdnb2apmy/oZbMojGNwPypQfBP+mDBB0+mpQ2ug9y7gMaMZnkC0zpjYG3kaxJ
KdzJv6c3l3Pi3RmiguuH8zi+mfCfPS1e7dLIlhAEIZSnv+kKAanL6OpufHPXaZrOYN1ws/ud8ka/
6lKtNtmh1AbsLdy+6mSkg5+zRwcgZ6+YHni+0P3nN/wI13UFPm/llMyc++GvcIb20M5WkYBQ/6bI
KUNW5PP76FV5DGXH876nY4g0EKCEBZSUSuu70QbJEmufx2ruYH1S8L4XX7MRHbW8T6+Cbelgr/6v
+l33ieF8TYZ9JDzhjHSdD7A7ojqQ9WgIDW12IZNrJzKPd57uePCAUjriA88l6tV29UvsdVUCaNhI
kOOdddFQryHwGaPDmiQgAlhBBO6KEwKgL1/k1+hMBE0RBWSUmMXmxRt0fHZXnke3u5yrPJtQmeXJ
Dcon3vU81Im18ZMGdoWgabSTar8iXuyyE3TxFnN4U4Q2AChOn1HOd+fTBVqkdAstAvsFXYfP8YOL
ZqtI5O1Tg6QdpEjFs58q8roZ20BtUVY8WlwaaUhb+JuIc8qhQCAkS4UU17HykJ7YdvD8v5ooUe1i
rdDaA0v12v4A3ccJNq3AjGtAdzRoaUWVxUJInYV21sl3gC9RwmKOxJRdpRpYYsmu6nhK3MNc7rJY
HGsiFNS+74k4eO8LJQ2+/cDGp2ofD92fH/MFq+alxsroJQ1WCNZab6czy7XqzE5LRz0qWMK1HMO0
5u5G6WgoE/UmSjdvcZpYcNldHWA9sy7qUal6iFOeucxr8ZZxtXh9H9wzs9I0Sf737p+jum9Pns0G
g/Bh6rs4s61Ny17Ovd1f4mpxwJPPaoOjeKvBttpRRASCkUW4EL5HsXwYY3E1+N04DlzZZDikyO2r
ZKxJiTkjLlCZLIGpKtxhUC7jj9R9DFjhRcEHGlJtkCXV/S1yjOmTQG5o580W3eS6/LLxU3ti2EPR
o+iKpDls35npPiErr3K6zVpMl8MFtT9i7ldGBgFjjBvQHeteakoUxj4HYh4vtZpE/YTGKBN9t3bp
s1lKjKCnA1m87KQn9B1+7Y5dUJ1WppMBTBB9FZ9C6LZg1bF8RndNQl8nRVztr1vwxNHAoSrMGo6d
FQQeCYADUdgFb4UaAjZBF57cMASjG0HrQtoEKbFoAa0lbapWTcGQgqJKURW6D5lZOWRFDML8/2K9
Ihk+0oY9h594+Xmqk+967ikbqsBLM7S5ADlfTMpWBaDbobsVHjLUvx6+PHeChkxSbgwtvuZFR3d/
0G+J6yE6wTT1UyBA/2XObmpU8U91Gqns5B5GzPjQNZL+q9J9Z9XWk7txz9eiaFXd3BpWdKBoxDyB
MWLStSW6pvUx14ElaZjg9WMOdQPf6pe+Z2OA1MLLPpdvXT8CqZaQY4jLG0z/C4QN46KhQHH5dyj9
LucuhXf8/VV9dy1aZ7pwZcu7Hviafk9rYmQFDTc25B7s/1GEcUjbCXhhcxp1I/nWyj3Py5XOuujb
+3LX8OFGB6ioZavCukhSs62evXqKfZO9Kah7A4KIQAX+uO+bV6n47zPKQSAQG8ps3OPeh4A1gm2b
kt8OurkIGBqIwAh5fQkpcLbsdj/cwLCK6sTvParZLsiqOcY2StJkwoVJ9KxMCprPr4miDNwgOkiP
C+ciy6rjWmCF6kZIpCaQhBkeW4ZZ+aJTuCXh8qyAA1RERGqJs7jmQnqdxXEj7LkaSaeBbIue5IXn
LQP5MWVU6eFdnERUyTnNNSEjFNDyP6NTQXbW0j4DNvy23dnw7Qi9eAX+8INKEZOFsy4EJ8QAbLEI
5VIVExKI1tL6komue8k1+04ij2zS7wRnUHXJ/yzvdurajz8Tc55Uo2Y3vKPzrOOJYOQC/6t1f2iR
L8MB4jDnqIayOxIj8paj4slMjNJcdh0vU9qLAGPBh7ii27qE0HEIZDYJbsMKaqHPjGDVLsl0DAfn
Raf70dzH2u+G2XaQnOAIEjC5PEopO8HusBr1cgdjSmYTaf9ZBHtE+l07vByyQZAuyikxAeDFIL8b
Rs9osmzGFvT38QA6cIGQ7YiUV46e3RaTnAJ7u7F53Le6mP+ynoU9o4icaAFH5vnZ8ysW6REXosDj
HxNKfZ6+MKbkGPK2fiSQrqODrazPncKSXBmtAE1ywvxwNnqzvUGH+ZjNQTQiJrd+r64HnVr/cFgq
PUcnZ5KcjE68eTqKa5XJJfEWFUj6X0JDEo7xOL12wYXNkCHyWVVLv5xyBObe2KnX5JRsTyztf3Cm
nAralW4wOVd0E5l+12CBeC41Z8pY0joEQDkDPt1Y6+to6Htwg2kVQN57OF1G6noyRfMUxaHp5JCE
PgQh7X/TelziVyM+TKUxiJV5gpqSJ741fXoCeBNI/AbeYd1bU61l0X97lKqA1uhiL6VAnRydNI0i
04LMjQChdYDJGwbF/dcGtwFwrFQue9P9pBrPFuFE99haLnH6XaPAvulDMt6KQUlC329lxgSFrq7F
a3PmrSSpGQKFXj06ixs+5MsMGA1MOMfQ6UmQbI3NKYoGUZx88OhaLbywHed5u98DRPNmFPEQrcFE
aGgiYfqqvmQIxsXYJuNxVrUJ1SaAazhqooNtYHcAHC4jkYd68cs5T+2IL/PdMjAK+OeschDq+eDU
0u7tn7WQ4WNW6HPxIqDBNVOZ7eFDjgpimpcFeUnRwm7NxAoO9mKpQmRNcG07lzzBRF8G3olMmRGg
wcu9gmSswct9v7+5mlFI83A2cthrHoVZFOA5eNwBwB6Ij6lj2VsjYJUE+dPu2sXDQ7nJaqnDg9RG
j45MKe93inb9/j4IA6gd/5og23NIH5K4w2qyzaPUMCx7w05zixUJmKTaiDDdgjRLNrIhlk+CQPrV
Xtyh9lMnEZJrS8Vwe97lnxARHQ3Y4olowcD4/NhfWMgrExjJ3jdoC+nDjPtI1xRGACZq/q5kvTKV
QihBI/ObKpBTG8LrHA0Zi/gyQoavJhAD4r4IsI9x4qIBLzWc9fmSMNdddkE6Ac7iBsFy1z9fQwVd
Cwp88OMjC07krsDn3uT9qe4IpnliXbZYBRxHrhmRvmSs2WbyRheYBufmfcd0OyQKubU+BRkdkNW8
20UiZiGCx51KEOTL/SdnwXuXESR88JXzMkvkduVftlAUAJiXVTsvxSrzyoft4YGlrLwqY8705Yh3
aXfDXS5gb3dfiH0uEeOeZIUT9nghyMH0woDBuHMmv8v/EpE7hbl2pQmQYQ91lD5GVRPNP/EJLAuL
cSJKS2pYyeJrcys2O23kkSu+FHmnoKpgcGwjiao+meH/55Xux5qauGCjQfqqSrjgkD91ReaJhreH
DQyy6Tg8+tdUX976dlas1eEgBD2bizlodHuyvy1f7N0ibvxUb+UkCnlypt96ixsBrLxO9msp64GZ
z7bG6Ei52k+VZD7ZO/EnAv+kQZA12mWAeKEIgPqQAke4H5tCVq7F9iQx4RVGx7ABikESIHov71yR
OXEDVKhvVWPIpsYPwk7Zrz7x7fQCwFevG+nAeToS3dYqPKrSqSXBE0QgHpEpL6cdLIPVtbVgEeBQ
hb4L3AIBN9/ulFfycW+Md80EH41B2HwOL33QWr1VuPdE8PPqxrDJBOqK+4qXk0GzUgYlKXZJWunb
UnoCGcKlqZe62pHDyZZBs0evDveVJWDscucam3mrhT3/JsljwF3sl724yGXA8SuA7damDa+2FHLQ
P7JaJYip19eFrv1WGI2XwVlhMirAN3PxGzJYnjMqm/LnCfeH11X2KorvA+aWmxsFh7pwGt3smIsS
6VvzyCyLeW++OsXghA6KI8+8U881YNIUal2tr98dUO4hULmEWLUGOTW8prwGXgBWX7noeQKcxupG
6jOGt8ggUxRhznnmj1KZvA0Jt013jvaKwW2Spl6zw22yvBL/bKHFzscrCrVVQW4mTiQqOvOV8o6l
zoR+jrbFf6VqBLZPUopVxYhiSTocD14iPLXDBZryzZkySg+7WUHx5316CFyiaVsT4YiNAaMizO7D
J89aJtqhPdl7LNQa5C9WgA0053IMmYGZBP89/JJBLplmle1S90yOoZ/cbeIUNjCHbcRepD3tNNa+
AY2/18R3jkOj3kVwvb7HtG2rxG/608u/VrUuRzblqNtJEbm6ex38YQdBtFiVdxxRmd4VKIl5sghH
YFZDm1oGwnoevkw7WPGuOEyTpFaQkEeBKZHh3LzjOHYhnaYAwnomiDUEytx0DAgcH5ztOBMSfBn3
jPLPkJIlGG89qaHIsjIQJC/idjDpkNay+wHs7vmXHPnnZ7O3mXOFjpaEI7u20eFZjDepYnN18UK1
fvGWW3bpSUyyYyDwkGbjA7Ra0rTTn2uPM8amcJVW+e/pUmmwJ6AWhLjYE52MHndWNeHPeauJJgsD
qb0USt5lEB9DN+icAEAT9PbI90T//rJcr7L70fHfNbzd7K+6TX7ZdWUhKBn3KnCIOks4jbZD7d/N
/ODVRi8EGbwynV+E9BRcvU7z6eTK5miP2bmLljfMtufvxCO0s8rBne8Q4JTumcSv2gNT9z9BhkBv
fe5ZpyoVOqGZXVEali5obBJk9oZS2j4T3VtJ3clCj3DjIFgBhFvUNxAdl+fP3u6k2SUicHsaS41P
OFEts8Kx5xF49qBUHA4aJ7Gixkgblt1KwWdFpZqjuoe67Og47u7MvrM1Qp9HJjNJk/a5troQEdIP
4vaQxtisSL14B2j+a3V7w4KEUhxJbmn//xr5dEgthue5Xx6/qJxlK2Man07IBt9Q9UEFAV6huQ7X
nDrd3RoqGT3et2vd8CR/upfG2LeP9A6p7lR/VnnS30akoihGEBXBLFzqUTAjQALp4zjdPXmQm8HS
nDMex0O5IaTEO5ranW+Q7lhkgOiY4PL0/F6CVuohu4L3Z87iS8fE5H8rOGrj17D+cc6LKaIsqkB6
InmQ4SZVgs6MrORtrcg3DbHZyo0OtfP6Vi5wiIcJ4BvF+jZNNhcHxMtXk1eFlQ3z5ZTdQay4BCqC
OXrwA208Zbh342ZplFxbSuryJUdn0b/+66xf7up2sOVTmEI26oh+GK40WRhJvcTSClL8Xp2aqQ+Q
MJjoST0pIdgNybqTUYT+Tu2Yox1YdDE+CW0FfNxHZ27bnY+pqJRWhMyvkhMVMlGssqW9kGCKyiew
uSbuQuyJUhKM1kcMiM77/rysk5HFj7DsK2JsuEYJPU0NyEmUZmi3fc4kwhkeQvxZtHJIKHl0KXVl
7CfMqc3SMrUruMCGNo5QtYN0/CjdR8KkR/ql/I7EsFUZy2j71YK9fqkfSoDjlTssEatbdCnJvF+k
N6Sjo/fGoFGYkqFxfVQMShP7VFf3msUSPuNGY6F1KiWvblgRVoMdEUaZNuFMJFczvXfuz+WbHH38
pcvs4nu+2Rc7RGzIvi+1cJaSBgewsLMYWnJewzNpHT2BZDnlS6xww7/SNUpzk70e2hgAj+Qjmw1t
JHp8nQPtw/fI5biiWpBHoKF+Wn7fjtPUbiPFE18/95SSAubqymhQaxq5OmkvOMsoRfR6pZhDQSf5
NLp099JjmZdVF8r5KXG/3L+iBacoX5znZLyp/+vrLW//ALEnuxSl+GOHnr8+/ybwoLoVZ6JIULKp
068l3VFS4qbmrBwwrUCH6vVAg32hjPzO4YMQDd0by5psAudsCsZrEnW2iKuK7A9dGLwpzQSV4iqS
IMcKVvlbZS2vpmsixQg7DDSlrF2qZ13SlqJEbeugljDZTpL4siyY6Z1E4Ou8kzBASXCayjG8HSgE
TGAFLfzEgMwx3v7Qi9Q7L77RODnTmc2f1H3ALAUkCrdNKX91W+Nl8shhVJxmCuZ7nYFo1ewXEmzo
B8mZ51/RMIqxHAUu8Ubok0BvAgCgOl6ywq6VvrGEGhoms9OBw/6a2KFh27rUoTqBzGb1UrypbwVz
Vlb+HYSQmLeDhf9nhQpBsVDVPI9ygdD4V9h8kZ3ax+/jD3kmpsKJ+TwkbuZ1VXEmdVqp4xEml059
YrF5o9OxUCMnBnY/uoRwjf1w0l2vIq+3JiHnpxdfOuSH5pqq9ATZPpUkOfo301+ZLoVL9qiGh608
9e4HSXbF9Oc5fdmyVseL4ZPoPENl6ZkkdXxf4hcF1sArgrYXx1V8O5Fxe5FVJFe7OwnSqrYaBF3d
+cNgYE06EWkmFmAyWLa5DxyHldZkETprG2dhmploIsxc41t1aaFWBgrn4upOKXpYIK0cXzc0GHrc
rprwRTLhr/F7rGd/c0Sl1tgfPKy0zBjVAiLpWK+N3rYgRNoL8ec8zeysxnEnq03UMtPH1hTcnwbN
ldHDnz2+awYjRWn2zOmCV8ckwOMPMdlMq8CxaQNyl1qDa82i37fhwTbp4NwuBLWWwoRIygsNEvkD
IGkRnuNIzo2n/rTQB83/Y3XtGTEQYpbE9ynBnXN/+6btEuOBca5HBHz+R767Jloqh75tfootl9fJ
WUDqZHl8hM0mzwL1tcAAlNSHzhhdHpYGvKT6FjN9BIC6GfEmOwo3NFDFemeNwiR04R+XQG/uV17o
XYcZhv6/Gx3hE91zwOXsEce0m5iMzO/EptDYulWJ+9WWjH1vO5Lu5oyTPsWGdP/MrfLRZQa2vENr
7+hslBGZOe/esf3jwkW1w8paV7yueEhYscAL7iyOqZsYZN6/f6mzYEloLHYAkMZUC1ljjBa/aMoo
9F6jurRYcXiv2ANJoZcW79ScJA/1mYCNsRmRiIUJ+JkUe4VzaY7jkQ2FVJk5BJ8H+hxWYXthCUv8
4r97BsZSdn/RDOWG82yhTGxnrHjkAqLBE38ALZzCICmXQXEy/Y0YE4fD7BJLm712BtwdlnepmDMG
xa/YNowEFHnAlXsNGa65Iey3+7WoaUa0ZZVt1TIAcd4VSm3OcuhuDLpkQVge7/4Kwgo0Fur9Lq4n
DxIz/v9EK4Ruxfwdb/K57o+TiIoIpmWXTowLP2ottbIiSG3D9iDpdebG6CGM4y0IEnmzkGY+lVai
rVSbQ8B5XAXT09VzTQe0LFh6iwe0FLTYdO8izdIH1pxicq5Apcr1tNiFQR7RPor/O/i6PTEAzTaZ
KdNTiQ0zE27ILtAVAdSvRAjCFSQxRIJyZKiMtg0KLrtqhWvrbDseO7r9Lo257cXSxGykAPd0QJKu
0pwhS2KjJUnbeEzCMZ30rHbEtH7sBlFa6b11lhydkU7P+q9YowL1bb5mOW067Dy1r65gq0iSA8NQ
a45LIDOSqnKWukR/TQT3Gt26mYJPpYMNgqak2zQmYWas2FenmM7148tL0hlwscUkf9IHjqewLIep
FDlJSy4OnYCuQivKwRtJ0O5jxAG34I93+YdtAW+IMxRA+EXIxzgkQe3jLg35O+shiwky2EQ05h3w
/47aVu3TIY7CeRiTRE09POK5dxGGVFRjz86W2NVuCydwjGpWiqRMa25FJ2aGIgDbwH9MJaVuCBdT
oxFUfhDoVrjl+zV/GwfLnoVF7UoBw6SQH/wJP7Auek4s3CV0qrl+VgndDSvFtxjvHK+II0Pmm8oD
B/lB3MfFwNrQMFpV5erqFHMyO4Tfna8DKs/DZjy629OqzHaoiFOoSr0kY6W+casZjzgoN009m8K8
vm6+6Sz5Zr2bkFpXBMqRbWvnoYJ8Csi0xk9RU/WH910tFtN4+VU7DIXpZkxrwRJCVdN+w+44/erB
BcFRVZTVYjRilx/2FObw9OGMN4YHEdE6FjCE1mpV2z57v3W3VGm4Imc8tdtF0oRU+R7oModV/2di
mdCH/pa6vNi5Amg5R9vrxVDWegqDp5VS09XPSVtGP/c5duhqWH9E+hHGiZq5JEmNRe34BCU06jj+
Kni2YE4sgnkZfMWQNKQsqFfopVItIRMte8Lf40bbqpZJuNAap0BLZaPegCwJXGPdkdDWsFaCOn1R
d0TCc7x/5h6bR7u5sWRuMNePrybSckp+lr5KNY3D2uCaAQmAp1EKhFl/7UXAfk9EzwIwCLOJSfO3
cJec0unYiMediOKbXx94sx04cZ+eqdhBf0TRCNj+iZadoOV/FnQdzvFjbmk1r1gWh/rSoodVggIX
W9wheIUHnrwnyDWoizsxAwwvbC/xwj276sAJkqqxudQS1at0HzKSuqdx2KaFIIJ4thiDY5HnXsd3
+F5TVrtij9PIU2lMPLZrbZ/hDw6ajdWfduip915zYnfpF48P7ZshaymjjgAhpy2eoXJ7UCE95Wal
f83Pdqj2zQDQR1QBq+hBYA8BCyFLE1bjzzXEJAoT8vOio2cEKnKF20JfxgvBlXLaDOqCWBDg8UiD
CXQmhvNirHLlm4otbcjto0Lo9jbmovVtrxLM2789ATsFLSQXrmypBlbssWt+xjHe0nRvCzLog0Bn
J2y6A9ThoSA6W1JisdichnoWUGQGj2At3vxHrRNXm5H4ZKii8moMf7ePu8egzKCf3dCjkxVm9a5T
bxCOuotF5W3t0KruYpE4aplj++LT0dYnkp/NEQH0XdXPuI87mYaQ+koK97nDTU+zBoWaNl3XxTG6
92uLeRQzF4+SCE2Yq1ZtKhcid5Jd/cMB6KW2+bNQc8Im9Xd2H+oS2n8f0hXfaGNx8x8w4+HS/tLf
AyipgZH0fz4ZGgMJ6M9dntoG7VqZDArqcIG1RR0rz5gjdqiIH42LMjOxNbOCr0PxlV/L5EdUq+up
PmX2EEe9ydoJLq7zjTT/P3AU/7w8Ng4dISCNXWh1JFE7+FEfp7aVv/gW1cvvnq+/wUPQTHLIr8va
j+h4Fe0/2iU2gQyWK78i9eiVR4FHDj0bmDiDEUgQC27HAH6InUDE2kMP8w9ctr1MTDLUSiYnSD2B
M30aogsfwH10A1I+9olNBUCMrvxA5N01OrXNe7/z/qEmDv8rTpP2ZCXw9kgCV0LDLJau0okr0inI
Ur9BKJqqS+x6+0ndo0c0t/KIasisOdYT+lVozuN4Bu5nWAdjtztMeah2nbSrZCoN5PAjhOBWLj2X
RUhPEYXJnP/DujvKjfkJUIC1BF9+gvXVY9mq7mYAFo/g2MUxoHexItYX7z5LsoGQ0pCup9dYBUUD
9WL1n4fogtOFs6OZbZyC27YuEE4fmTeBXQyRHeLmIffKfqWRYe8CxL2FwJ8ZMadEmn0whvuYMeno
LW4MO8F6PCBy9guE/PGDNYN5kWI9o0hACvrxXHc7TtXY7GN/wZP25tzMrvWGtoIzDnZyYHLHA4yK
F4URoaS+UcvVXKkCfZQMYsTQbU0PqqK/YYFGsbrQhhKQQFBBu0ZO8EdLP0sBS8tHkQ7CClluBkee
/raOzX9jDzMBdWtR6pza3NubWe9I04gOkIfpf6AmFTYQN+gAEk6FNMT6Z9Y6X4MQFQtR5aJuEusz
ROu213nuVjUYUgojFxQZuO+ie3eqjbXHbIczFbDys+NCAONDGhSgBBwVwxPcAk/bbIDe+hEeB637
Q0T5cmnIYi3wHlU0SERz9mNLcv0OEyhIPnsJ/SoV51BU3LfhB38z8qQjeiAsqIAAePkKWZOMcVda
vjpu1vez84aHgSmU8wZYURjS+T+PFqOQDD3PS6r8K0nmyeigNzJWn1dXYc5QJ75TlIN4J5yC1Et6
P0Kzp0nx4JIfr1QEpuncCQtFNfT9vhB0Xs+EwfI4dHOAr0eQ9dl34Ci3kXiuy1npIhX6yCqNpZRj
P2POaY2e4/IfPsfimvs/lhj6TOtQao2juGr6k3AGxEldzukFso/FjhHX5XM7j+bP/ph5Pjat4++E
XRVQ3avo64ljGaHJCVElJ74XoajnLx5FG5JEGyk1ANJOkSncXLrIOS2wL0VI1QYnctCKfS+2ZkYX
piO2GDjLJiK0JMPJ28gqOUot+6ryAL0TaAvlIQQZ047P7wUPVGNTApVS6N5m38sXlbog8DwMqg7a
JsvzhhLaO/Nqxfl75LszKNp0uwrTFaJD5CIhOQ+hIQkFbQsMbVuSFmPqdJOAg4rz40tqC+eC+cDW
eJvYgidunH8JgbvEZOFlum+2A9vOFWopmVloZVa1J14/tg+lODPfLOW1t47G2+8lRCH/17HjW1wp
S4m8c4e4SGF/HZzWzfZDDS7WwzBepGSXPwXg7tIW2QlpK91ngdziWoD8Zd5iEBdrCKLBmZuv1ZW5
gRfWB/AwMiQ2UBCwSa2Y040oIy06OKq6qc2sZYVMsxJDHGY6h+Kx4zCD6xRnSBHmE9jKD7sjekxb
sj/WvgIXjyJMJ6tQsD4+4BTOaMG/UwrGgu49LZUDgH5po4RYGbhLZ2G3BA56DfJ9tFIGIt5KQYjh
K6Pt85FcTl7H+VKgpPUAyXxXNGRPUUT55eicoQPOz9vtMxye7kzQe/WVnTMlljhoSk+uXhyx+Ptb
a7tqFdQ1QGg27J2ciTNXIaetQem6kJrBhFBkPjxXuG93wAn6n8kDEengCX/TbzKsjC4zUCbEAO8R
MVePxbdMyXPCn/c3CBgjwVc6eyB0NaGdos2QGIGoU6tThfFIvGq6JdoLL7gtgJshzdUcN2upRUnQ
sELrV9Y0mOisgqXrgkazDOcPF/z2eIlSd3rFi8lV3yL0KNbf/guTL+JKzvEdUANxL3eMI2fwFKmD
it93QO1LoKR/URlVxBq6VFEg6Irvubw95yVBLN/DsQ8E4Q1cDCqQt87M1aw29LzL3yFyewPCLGaR
v+Ji6rBu9IIrQ+3vTYftxEmd7WkqKs+3v89VWRLNo1Slfyh/x3VPabxl7g4d+QGWfKG9npqSjBxH
GYald+dzBXOtFmmLTbztJQ8SQ+orTMU7leWbzqApnKwBBxbPX8+fpgbTHTOrsaDjtiUQZX1Z3aeq
tKDLAixiwSRPZZp8HltPP2XVXB+wvI/kdJgeDWUEwCcvXy/xQrrJIFvaI4AmNOUNiQHPHEMpHav5
FzWk78vFIcPfC2F0wxM5ranfaWyvKM2GekzQpGXNSL+gR6js992kqgor55yLxDcTl0RXhrTsu3BT
rC9H2JLlezBOG6EoaAO/skGWkMQ5o+UfTWvpO5+1RDLKuTuQHfHXo9Z5y07POVOTpwy9DtFy+X6g
NDiN8TZv8sMj3/7qfpoCp9UZAexuoC4XukB5S7M0j5pkb70dzMnugdnoMJgQV/gDN/iB0R3Y4njW
33XQ7T1oUamqHOnht9hbve4/ns3bsK4B3tCmZk4K7I9jzIp2aMGL+3xGBN/4Vx3hNkInAPlbLODz
cYud+tJseWtg4dENg+gkY/K5rPgEePO4RVq/6WyYcfc9vZmQaTi38u3bGaWghvENSw8ntx5tPjo/
rJ9Vm1/UtG9CBZy70QcQySmEz936PFuD2Lf1y3MJ4i/aP/ftQrX2QrR35ei5lcP73S6ghd0fiW7O
YHSFxxeO7iA0K/teFk6iwcejTYPXRHywD/dGs0P1AczFUkk4Oi3J8sjz9LwsOMfGpod7cFrk+Xkj
88q5mEytiL4XesWngRU3XOfO0Rp+drezJGst1Uz7mhWxaUAkr+KBUdkulWoWlRVmDZ5/wew4Gl1Y
G6XMRB+shKb3vbf6rUpRHzQBj1gh74SSZPdSHPpb3ZFyuyvJ7v2X40P+ebygjyykH57rV95B/A9J
TVARggHKufNaHI4rbHx7XJsgh5qhxb41Zl0RoTmcQ5MZ2z1N6qFhxaRKBWIIDtqje0/GqQY375XQ
Tz8IMQqzJLBOaoyG5avpE5hMTQ2Hg3wMDGf8yY9lnfGMWo1mkxnwQ6DtQrCqyo3D7ljxEoKxptIP
NPFsboTIEcIuzsLcehh40hqmAWDZWumHhi55TuISLaqzNGfSxe2/X4ckzT74H0hLNcdG7d8PMLUP
DhwTmKL/66SVbydJqYeQGC2AbQ2mi+iB70k/pBFPqF4nDoASXsSvIvt3SFg8+d67xNioL3P/sIft
GcOLODnGal5W/DWpW2RdRVbqOylWRx7Oi4fnHct1CvRwcGgHGiDEzP8mk90/nN/zH31n9Aw94mwS
lgAK+zMFQHhnkgJRfyd7lxJG+UwDEuCHOnwg/BDLMpGffKt8uMZ5MOXLAA8c23bW5cKA2dLLupqe
BBdh1A7fbCQ0Ga29T3IquWd9d2nCjDpygTGypyAlE/6BEN/xbKFcmFnUBTWlG+IekRPMG9C/9wNH
NJ5qxKj0VfhTvmITylWVw1Zata6FkEBCqTB6T4dgemxj7cYCRg5SHAEyfmknSVe0SF1OjZKuV8B9
+5NB1CIndbWQmcDkmvNlKk1NMAZhNvFr+JRHygD35DjzYoEh9IBcsqTxZcts1n51pH7NpU0N+AOD
rz9Gg1VTqMxpXvCzqYXqwkjLatPJXoCx46mb4MvS1CX8I5exPOtEW3HZMZa3PP/HaEQ5JKtWEYCz
DSr2Ev7BvDEqFteSlW3gJad71TnHhYTsK39sukJNJ6aObn1sDC4NsLrHKxhXGx2GnlhuBW5fBaJn
Btna49inbLzdjr1CS3EHUGjQZvvcJfSZWQKdQtKe7Ll4g5JKWiqHSiDlDUV5OTGkTeL0GOJoWYmV
ZkVuLTTZEbKLPvYexMiYurdxTf6FEMA/vkgcqLNoawDPw5T2D3HUh0N//mXeSkKwXfHFGEOCxl9H
xolZXjjY8sa9M0PCvlGYOnAy4ulmW6ZOx9R+RhJoAg1tmcBcMSRiYxFJ3a+sYaqXqtQ8NuD0tgU6
5R8Zp/NJVPd7rvLg9m8UrNPBoQowUp0sjnQ5PDc7xB0GEIXNbFqy2kQYMqRfxC1QvV6H7wpFUKN1
S5FY40wTEcGb/ne8iLjI2t5cLHxSuCJYBXUPIcYUk6FRQJaiQBLbemimSLJYuc5IUTqMSrpR57ni
ouJBQ6pAR1ZfemaX6weM+dX/icEahKXYSL2EiueVQ9eURyS+PTt1Rtlmo5QGMdwtH9tt4pigvccw
GH1N6QPLxwt54lJJsu3qbcpxZ/kyXYjDuSwCKkGIvHcqTtMBlTuXMeLEb72umIxnlYkhWtcauqkP
KSCixVbQnzDndXVAUarnL5pic6GNmYsk3M5xNSg3i2/xfsr/O7ynXo5RUxuXDrQJ3jr2iKDaYzyV
VOkcQ58eg4Fm4PMTA13gIW4qmvJhbR2IvxgauEaYcj0VUCfMMGSSyIVM7VffEbfYAaKvc07h3L30
vJvLWvaP1fuYneArRCsvOFUhvW6pEmpPqummSfPTxjuO+Cve3hc4QRoFiilRu5bYmGBHNShZ9Xx+
NCAIdL7yK3cGXyS5L7E+RmMRZ4JbWZZG+gDHYMhCAevy5EsAAtxT3xpAT4LWg5bF4166VqhIJoEN
YLCBUlEuKoJueM4RaCkUi35WJa9zi9CqNxY/kF2Md/Sx8M4lWnKQVLQ3L+3eCWMfCeD0EiwxZpD7
NTrz/72MAH3nr7hqJGSo5fDjpH38UOcZqg6IZXXFoXN1tTikxbcNhC6u0rPtHv4ydjl7bbsql1qE
Acxh7MQs0tNgITFPXaLfxinY/1yBywQENVkwwsrHXxo3sIY7fAvxLvh3ocb2oc1pDJKCD895+bxJ
B6CP/96L90tIkp2RtDukoPV6fj1FjIJGPqgtVX5p1XuuHlo0VGPiaBLK2NwA7fXQssTBVQ7vDK0L
wN2KGT0USu8Vez3a9CZU/dQ9sy2q7iyWfK808prnCXzpEw4ED1+7qneQETKxbNUMPFA5GkRc0Ln0
3P7IOonEglJiYszi+HnOAKTrHUIbcT9hLmGZOuNDMbZ6Iwlzz2RdjyQ519js/ObaEWsLvXqSN4Gg
clYAZYLngge/uaofBgOhn9hd3kqPNbHtcyUktQzCa/si4FDxKXKMwMlOcqZbdxUPWZ0+onD+n1eH
CJdp5I0kp/miph/NqDhptm2TogmlJvQCd8+FK6YxC3zvASUzDMlruIZxZO/dprB5whr/UbBLJZW6
GZWPl/M+nSLzl4WrKq54aqRcJSSZeWSEpQSUv+HOAPhmg7QPSIMuxQ/MzJ7L73ShSwgh05Tj4iGW
7yiJnqZAF8OGkC8Bf8Ww8+bpOrkFKkK9b9Dz0hqpsPHCgyRlh46FfyCObZSqbqw60kfe0BpWA0QJ
rt2WFmdqaHMfCTWCKWM1EEmHvphdI08LSxHJk2m86fT7GOM0HHBboindY9Y5RFmwsbBEXIX1H6xK
xYe+zU2YOBTrCQ0/rwALILjpsq5fyHVuRxelTfaD/yCJbHmMJvOMxe73FqezeGgsBhuarFN/qOe7
QwBMBARHCE4fg/Fo8ZHoQw/qVfbUICrbtmA35SXkd01SCtlouPs2fpaIfwtlrQdncZaW/SToEzZ1
Y+YXlV5GOJR6pibqU1DkL4vxCl/mVN9nyNpjpFJ8a/icOj3kEUJXkmX+eMkYrZhng7ew9sXv3F2J
5rxvCIgjUCAFBNDVL8Eoqpoj/S/ldhoCknz6Ah9aZD7OgfjLakGbfRntW1wvOMkxcuhXyP+BKjNZ
WyLVLl/q2z582psH2uwvXol/8QT7QW3IavoGking7lGVkOdRVf6CWDPmnKm1/fY/M7u68DhvJ1Er
NpjC2qzCmhpzxQLXa8uYwxkrCEZfDTutYv0Uh8DiIyU/kT/W3ECDS1TMHSuuXGuHMNjvOCZkrh+3
DvD52L+0qkVaBB9Jmug0TDyGGOWNzyYp2P580mtiC52MmMNQCb/FCUvbzG6Mu2w4UNzWptXCq3yt
er4jhU6eZBJVlDX07bwrZ3DDU4+xt8kArLfmWddK5dUWbf72nxZdLD1yUG+AV+eIJ8g+jmEAAD0n
4b0otihm6S5C6GBofnHEeCxifnk+BBMQ7h2igDoiPa96NDYx4blqd1DWoM1Fr1JZaTkqoa75VS2L
ad8cDt/kofqDCnnxZmyV7IJ8Ywmj9EG1LEee66tMolKqrBw6sMTASrvlCCzBbVRQGlMGFBbEMaU1
FBT38aUpp2Z2w1BUPqznOyJM+m0rpa6r/u8SizcUIvhO3X/F6qlHJhcD4evd0kbnSpipT4pGt7BG
KAflQkOjVlthC4BwfcaimP1JNwZDD/NJHGVs0TD/TzCmV+6idicabJy5rK7Tk93+Q+h+RVp7LOpN
8AHSo+U7MdM/rxC4BKtCg7NFZ/JPdLJZy3M5JTGDXzrbcPZqIeWkxX243FO6EMrKBmR2Ek7Rdo51
fjVhVKeHsPW0zg2EISG1IVyALAHBdT/oefAedKQPOiY13tV9W8T+0PgK+rBcrenVnvgB4f/j/eSh
AyimL4V6UECNhtWCxOZhAy24dA5wzaBD0C4BRD3+jZSwUr/dJqj99rcEbx1HHMpCJFqgGlWp/VTq
pvUJ74J9a23Nj2c9PtTA/bEfUQOb2AbuxeFVCGST7CB46FbSNsYZSVlDzCesHDUUuV9oRrjShgrH
0cyELla61wgWHh+bskR+kAqivzPJGZ0sJ69DcASj0vJkQxJz6XWfsnZrFWPIGsNZPaxJS0ND3xNa
L+GCiU5R8AnJ1xL5H2WhUffbGOx6CD8ah5ZGIT+K5YHyUd4IFS/c5anNTVTt5tLNvjp+swv7y1yw
pJZnnsTkaOK/iUek+reUNlL9Je7pbhJA/8nsqlz8cEwDGsRQob18XogqvL2qvXMaACS0HhGvQt7Y
3fMfEbc6IlG9QuntZXGQMWSLaw6wToTP5bzZNKiBGeCOeasLu+eZhP4rPnKhRRp+/mDBz76gYegI
xGJmfGMfPq9AiPdscVt3eu3/D7whkoiy7i9VExqZnJ8Fs/S1+VYMAaDkgeJUg0DegLNhicZt0FE/
WIffqs79BobGg/7HuNNZTIGDenRJKtWNQ3aJ17EWqRkCso/WhvPSI7LzNExmDzwQQ6A/yY+owIcn
hOnptoyh0xaMY2qJ6o97w0VrmxnU4T/vnS/feBpLXaITr7MvkRjjGwK/wum1m1ltJnNe7B2xOjv8
aka4QWG3wvU7VEKovkzwJAu97qsGPYqGq2/cKaYf5s+t3Qv3b6R5fEQ8hzsyNTrdJxi04OMzkYu0
W1kSn1jhcVHFrc6y7Ux1fMinOMz72kmXmCvE8Jqt1Xbq/PD0GqlZ3smVaOK+Q615V9EsAIqC+Iz/
XEEUAT6TpmAX0odpQEKcINi6zhMzIPcdJjw9TacnvCdI06F7KoEgN+mSd0ovqd+t8KkYTV5MV9uP
ddtpMOAgPImn9bmKCSt7+MkKAD+QmHKrAKBIMLnrHHhUeJehaHQzlBovZGGdD2PPU3R05avSZzDc
gsCgfHMHHoiW847A5yaVoNgLQLvQlVhc+FyrqSm/+32Hqxkw2YR63hGrVWQ2rqMx3zlupWEm/zK5
7KwxquySCVlMPPN6OrRczUeGQOxFwdh0we+/B+8NikZDctg/PqbQuR/jdr0pjqtIV7JOaNC0/HEK
nokIlxVSflVUEJKyUpSPFJbCxWjVmITdrm0JC5tD5XFkM6p1qIxm9WDRX1y9Ss1ux8YeWm7m/4pt
RmvG/BxKCRwu/G5lMcCU2hHDy3oLEVcyB/CK6oemEaru/ajW+2GPB/sGH7+CzOWBmUlCbKTZZy3I
H6qCgI9ckku3udFFceGjoLYGgvvgapbjavJULHLJONpZAvg/ivJ+FU0YouVX+7CF9BGExYdyqO33
J2vFkQbB4Tx9vsVkAk2toUO1GJjSeY25qOXH3lwBi2lRMap4u3MdyIhgIPLi1HNuXF8Oypv3s6j7
r9PuiO2rdcikF4pFgRgp+CjNpZ9+pmZNm+PG6ZmuPOLhc6SgtDmnavVZ1NhEHCDXdnhSRQhXeCL7
n3K28ExZ6265IrwnBlvCWI28WUcF7dmzT0uEZZ2gTjAUuMg2xWGUIbXP3VaCsf6gf0FGy6woUBJE
1+sBHR2XGXJJPlvX0ZkF0/XCC/LMgnrpDQb0qHXW0if3/RP3XhQZIdfIm5wtO7FLdueq5Kpp3R9D
c6sMxSrSKPFaQY6e4BKzM1SONI880ptcgMnJUCwiDAFguX9AsKli2XuhUQ4bNrUF8rHsMINbLpIv
4iDdD6hylGibrGPqbq/HxwHKq/MuzXPhpu6DtTRJaKpGqHFeGT0T7QYba3eQeAVlZSSLfIkWELzz
K+utkYCulxlGZoNXM45WGXh42DXz6oaI+6eTvh3xLv0dIWEKcytmZzcEJc+SPvNnVutBLU5PKSBt
8fXprpWBd9yt3nX7ZJPzslpl6ITkdwDdKySNvmx7nsQ496xVvIZi4dGBOya6eJBSi++/bbOgzc/u
q4IYplau0TLTvN3adHDoK4hxxEnNglPVmAEgWdN2glBa7nbvbEAKV6sP9FmyRsFjNeY3wUEqgt4s
5odlKxF6RqbXpiKV7KbR+5JjpTyTRKeF6qfPDAMFMXo15KwfLRI4oqdnZb+61gJXOirmqnDl44D9
UGN6XquUzjqRP3REQquOyAIdIPSWCAeD1nFKhJZ0SJ5P5wV0vdEcUDmyVRptngQyzDigaBC9qOu+
xciCTc3mnJbQexdYtEHWkGJjO2/FcIUn5ZPjnqPmNJJ5TpBIpBD/6ErpFYmL8AXexbA1NHYBrCpK
6hL4cu2Fi7fNPSl7L7jY78OdPf2Ma8o1qAOzN1LTDnqbwf35SL6cl473ixR3gL/loMqXpn0vUM0F
/fduIeauQk3MlXGMl4/LPAd6fGvyc021ulYvkfOiLnyPSWjShC5EfzJCDsaH0jaJoG0MIipuIvRl
UxdmlFffpmubJ+W8owSzM/6fowjWPXOuXAsbCJEJshN5EzDiPhFk+YAfzfWiVuaz4jGvPBhpY93D
Xb7w/ET5ifM/mYpmIKgoli55mIUDzHZ8Qe3e3rDrZJszuc3cVxOly22Q4g6LxQMVQqQW4Op00PKG
C1JhhGFFbTLMvu8DZhNOcLM68fXkxsfs0Ffn2T1UhnD26+zpPnZ9UGZ1VsAItgzNpfoTsSzyevVA
2iMVxUju0uIS3fl/pEJKy/IdrebHGgBLPJ2ZGboBr1/lpE3oyPKVIUyXqpda1K6gdr6g73qUM1P5
7MfgLjRZdurt+lvMd0pccI/5rshGTaIJEMix08tFuPNdqyW9H7ZzaIH2x47WykWexErBXjAwCwjq
neYHZMsdbbv/K8AN5GLQRAMxYy0c6cXxi5iyb3uudQiXYLlrjwkfcHovA2qPPsIM0eXlA6jYsrR6
75IXsda+bBNJRNn/9X9H52O6Rorln2gll4xpDIj6zUzdBwLxEDg/2H1cET2PH06Iy0XYaWGsm7Pn
oGIoRL9TQZ4HwcEqNUNr9Pm6Zy/Kzyl/zLYsKCNuIK3J4UKCZbKYwIbZpUjTKTNkdzjuGvy2sP3t
36swSlUEyu56KhMI/suaWtUHj9oSMWZ0IOWV7RVaIUiINLOn6p3VPB0409PzTvkfE52l4Pqnzs5N
bM8W62X8NdhTCjpnKQ7ymo/gBZh/Gqo1Ed+CMdMxFx9ErimJHlwKOyPgSY9m+tSaNS04ljFh6vbV
s5/5ppo7+u2moRHRzjxfNyl7tYmKbf37PNhlwH5+iLYOSwUox3PbHhr+tcFUnHPTe1GoE/GqhSDe
9yhiiliMlrYf0TgkNrzvtMsx8wYWb5lwIewbHrbbA3HLPTb8cstdML8ggkmFhAgSKe4yEWqOtStQ
Se4GaULFzS8qRM675WSJk/9LqiGTkr62FbFBR66Mn8okCNRLeVEiszfwx2N7k0AnxGREOgb5x6q7
cHJ3x5zms+WO+jsUf1wPPCZZVnXXbKAes6lPhr32AgRC7y+l/2GBgsF7z9pBHyQkk9YDtpAVFd7Q
klu60Y1WpwMsJ9ptQPdGTt2YggYzcRx2DFvbxmti4nYrAVYMKJGhaRJ6QQca0oFZw8Mch9mnjnUa
9I/mvE8P2DM3nPaCm56LlvzWwR2yTsj6l9ChIlpD93c/FTjbYyGVgCP4JM8Ckf6JXaXTjPxWD+Et
Dh3sK7HIK3npUctrFjUbFG3zC5om/l2AiWIOEIa6szmd5icacMI01W415U6c9fLoK+Y17N7uEJnE
DfhZOQCK4n9QkVZ8fcijFARS9oA78n1NbJTAvrTyNKPPmipdl0VqtivtwfkRGavBcJEDpDHw8HXm
B/rYeebPV7OIs1vfcwMrPRF1UaOj5LnJqyQukGWrmNG2U7VCeWMuxTvgdsEW45s2TLsdCexfZ+Hk
CnX/z3/WPOx+FgeOmKEfx1R6Rd1UDFSLl+pZVDl30LsNBj2qahVPicVt8ZAg6/BS70P1pf7LQbqX
hqM5/UFVTwpxNms7bPANiEgtYnrpGI9LufzKERYz7/AK13wvLaKzeIv40P8+lzPZzeoCuIp+Gqa7
iOxKHQiUL8HYg6/z9+D6JEw7x0VpAEHgbi7H7L75hhUr2CU0kI/VlQ37cjxJoq6tRAcXFYTNa3nT
yzu06Po38QyPg7TCt0zYknYj/3lZLtfRfrLPtLuAVxqqdcCOBS/kJ8EbCvb6qeYTWEx/MLby/4Xd
Ekx44leqLUIuqtEvHK4vIYlRc/+U40Hj4aMx0oCkUkNLzQ+QYn9p1pbcJ01LdyOh1zkItB7/e2mA
Qc5HV92KzxE5fnhemsmnlxG3zhQcNCBI4F/m2XPQ/ZhrmETbE6PVs4odu7SFQU6rrSDMKOkmxnEm
zeQHOgPoZOVYIwxA5UCv3fQeTvwuFCS1h2gpGZSbRKGE0ce2OtRYW1ta8UfkZCQplm90Q07ly06h
ic/xAxz3Kno5a0l7Fl6beXlmm31QR57GFhG9sSy95tF6BseIhDizc4VUtV05qBaT33WZeyGFYydf
dpCoJrtq9vKriqkGRQNS30KoNxA+Wc6TCC/K9iabxX5wqrHNVgdqoT43rY46Rqhurtbv4NJUG3Gc
KmeoiTXLYGLRnGOWvamOZVCNnFy9ERyv0SQpsyUMLlwqlOeFR+A3Of9P3zd5NUrn9baJ66kZe/I7
j434l5+m36V3sC9f7+Rggj4fP49R2WWBNwDva+1pDg/9V0LLfQg1eT2eL5241XeohYIiQKRAXXYf
5re4z+cJX0NN3siX15zSw0zpS8o4RqlTBNqNR68mmU594iTam47Rx9cEJXlcFAbqtHSE594EDPTw
dCDGptzJYdj/TKzlb6shigNusrrhVDHL8UvuRh82QlpHDgG8Qg/6lH/dwlHZoqHb0WQmJq66nTqP
awbLSG9jWBpt6qHMirinZMuJnkav+j1oRYJGf304vfFqaIbJJPtNC6/61AYQ2oXmzYayCu/mzOu2
4uKuhf/zBMcJHXuawxvXo5o9xCE9FuB81W1i83f6XB+euz4aeurC0P0JYpo6zyj4Qt8P4II4zmef
Q/1Gt565ZQvmBM5jGvEgeVWgIwEx75rxb4QRRNtcsNHIFsAuYG2iQbTsEaf6EPNfD34RcEx1/CRl
Sh/uBV1XwGQzPJsI3rFM7aTfq5iJotYKOo4ZIyC2O2av6ldPSyqVJZCMQmCLVYhsJ7W3vseGT5Ck
oIjk2pD9MIbycg1t53ZI+wiKwGiTFzVDciQkPQgacsbYnAQprILnbOCng2oN/igJZOjolc5s0xrZ
qbb6roS+OL8JUpN9k+zNcYx3K8SID0SP8F/vuPkyM5yhlUz89G3C2StixngTrfkrpfAlTKoNPv+Q
eiHUicHoIB3tiegF5MgNm2OpH8eJAEhL6gFHkVArbWddNs6DWUE2Sb3q7A74QLv1GoMzcdMIGiv2
9syortYExJiy4tWamKjvXxBShSJT1TH7VkvjdFCn6p6FN+ur78S2wxaOFjhYxmE21JlDkfqMgYsi
YZq6DVQ99Y8faBE/LlG6T82p+kkRLgjMSvQMAGmRuXkUfzaeLMyvq8VvgaEoaoLbFNnxE6VXRV1f
n5QuoPULXojWUXmOEeLzqF80uqbFBy1lyQ5N+3on5FajX/WWiSxyO+iqyr8F9S85LCurulEqU8uc
ctuWYcIbEE5pDnwWNexzbOcRPwWjRF0V3P3gHjphtdPAOMsk0tC0JTgvwSU5K3TJqsMr+boM/j6t
5Nenvqi+kv/xFJ6SC6VeqiziSEYLix9FCJ8SB4jecguUxzT94pwsgMGol6yFcA3FZyCfxJ02iq7G
UlwWzsnYNuzgTywQLSdKvZ9zkWVrl6jF9ugDOD2OsnT6XcnLt79UKOopHpqLHvlsYalUNbuxCqmO
+QVNozalu5Hxseyio/JoMTalGlQUzjdPKKwGkx1QJANiq/1awPM/sPgM5c9M7a7yCHI8Ubo8KB1K
py5A7PwpxokZIaYDHlVCEyZP+IagbcHCkseCMwwC8c1pxG8XCWJljKpw/zkqj/dk5ynPfNxDI7oV
IEip46cbbMogyK88pc6IgB+emiBKQjAcOXHTROmLM7JE4AOLY+2PyXaDtoqci99gRPqys7dMnGB9
53GjO1M+Jn0mplXp6+2aIMtOEqEiDzit5MLbmkcAZv0ke30CGaeWZsorQCRGpp6ugxkKs1HsGsBS
oM0p4u2JVaerPPRYC1HdhV7JLmlMghxW8lZFnncb4nKLDDIMw/QuXEob1ERO9fJCm117sGUUkz/6
z6Lm81X1wkwByUnHrDyWNvFnXWhOPMzg0bBfgh0cTMikbAExI6lUbLPT5IC9sljKWcqZIh4vHDZb
qM6aHjszYAUjsjf8wp9C8pjkrnGuIu8cRFOEpJuXSRrjbjsPp9Rs77fkwlTnZI/obd0AAKzFaahg
u2R5iwsRB0hgaRaeA46btM6jg1iM6m16R5Kg6zTrrZhh2tP1SE8Wi3C1eLhX3dvYyO+K/3whWfAg
ZT7gE7AW1FDm14d6LPese2oqA+Kty4BVbiyHUdgkL+GHtQEW66rQsDhotprFu13jnZWXjHNRcU6O
u/j8EDVE2gQdwQ5fSA7mltNTnvKz1YaeBilcoZnFK2O5VioYaIp/TpBrpe5Jq00ONnaRyudITI0n
o0AVOzOdPjP9uQCnbDV6qjVW8OODic94c1czfmWXzZ/dQA1n3OYGtvs//0hYnDRPcJ1fnKJ7GB7k
jFUDlg32WZONCRAF+AYcwHXBzvWMBg9PDKdz4n88I4ogFex8T2O+KLQEMZGBeldTPhqkbF+3KUaE
EGhoMa8LoZtNx47p4T3RykzVf+6FkS1P4ux5eOpn0/IpltxrNjdb3CCb7Imp4bu7qEuGzg/H30dV
2ZWZdJgq+nFPhLR5ZkdI3x/DtanfNWtyNLdsm7YlWNIGn+rL+Z3Dg0wuEl+CjVYcfTBNM1u26Val
HLV+Zpy2mpvE86l7u2j8TN50WHeRLp0+U7PBoIi0eWXI5GQwqvn97gjRYeO4vGcM3Kik3u5Lf5Z8
XhNmBQy/b3Wb8Qj/iRsr579oR/Ol5/78NL56EGa3DzVqW8Zqw9+LWBRX+4x0cmt2IRuD06smAcii
NkKEzVjTJXy2AE+fssnu7Qc2t+VrsMviD71YQOcMI7VFrfjJnCYpUCzvjtrO0GpMhaFs5wg91l7u
30aqArWvhIQagFll9q8Fv9kit3PSlrWGpUZVhUVvhBWMWY2VhHWCNhvitEkKbHyfqO4fxIUk455D
4f2w+9d5PO9H1cR3dcw2iAiBo36m494H9a6OHHGV+94Y/WK+QFUtqGGmabO77uLJvplq0GQPvHsl
1MazTi6jMniKSIw7W55NJLKfF9fgMCFQ6HH5iBO7qjD6KQixkpsDjrdBeR4SIFWB/3kbG59KEPgk
mgmnVHPZQ/Cb/jO0WhJVDE7ILdUZLne6gpW7qsQB0eIi3jrzI6ml/CEm67CHvMQ+JKpwPDjt2se7
Bz+JNGut2Dh4I2C9F5qqLMjudAAxfx+GtLztDMD1KW4jIr7L6bwrmERskv9AOkgWlxhla8++69OF
CFW6VddLfUy1qK+8PpVlMxEnE07o/1nF3s9yubIaiLDQP6JRxMMmlk3nWg+ltmyn9foAx5msflOM
9YLkPyETkjhM3LZK0h8tG5C9RBwRdnAn+iglPg16dOUktC5RoDws2AVnperRQAiRKMdPaYF6Fc9c
DLadAhtHzgUTO6VHTTG1+IGCxyb1NX/YA89IVf+zPTGPBPvFyV6Zsie3f+ANJHmCDizHK7OcDOxd
QZLJncLurqY//YxtaOI6/j4mLfuLs9nc6O04fIPyfHDN04TzCAuA0Rp+c9EwVqK/ClD3MPqV0b/v
B7T60jfzG0f+FaCYN/+lkFPZ3UJAubDmGvlqD9ogA/OuVZurDDHw/RhLjO+kI7CPMWkbaBIw1/hT
8ffpN2M/oR4Ot12UeJKd/bAVNFXmJ22ai5VcR24gqhtlVa/UMW4b0NxR1QzPE7kV5QjM4K0z2W5A
2sCj7rJFm2FleVA8vZ+BMBVurh9VqzmxKNbnjfYHjkZSk0EhqE89R2faQyR6ARalKqj1VLxuyKm/
wBeYKAeSvaAu+OzsE6A0RQy89ptdkhU6D9kRntnbiQvCWoJ/iGwGbNGoIV+kCNYTcNOrFopENUYK
QT3ET0Cmgs2peabZZiuJ55EoV2QM0jdGihlflkIEsKR9XoCdXyozf2TnnFCMqFK+7r91Nkmka7Eo
4DUpFKg+MFnk8/wZUhw756R8KDrMySQ+7ZK0bI6dJWjFK8+3A+MslzDPncpNl8iz3qC8LsbBR6Z8
qnUgxxKVpiiq5vRV7LRRtSp8jKMtsaRPY0wEBWBZ7T9vn/TIsb4m0auWL6AP2EDjzpMq9PgYXdKw
O6E3WWMb9aeS6laV5Os/MJiEK8C+QAgn9mluYO3Tu8GPwO9gvNMgxatAXkwCrwAT/Uj/hWqBKcFX
QqERdqUEJw5ZHkUg6SalNpU1USgIVe0yhi9qzBxuTlbgRMYdMiLZbBwKwG2i+5d+77VtHz1rU2YU
g9Kj2umf+Azo5TbptdycnQJRT7aZN2zG58z4Qh7ktR6jD0Tnc7BFyBiKDytSngqemKnlSi1gkrRo
gpE/mXDSV6s7Gf9d+9IKQtXOy71nOX1I5Qpusp5n1w62cnYcz29ZS07HNOKE59ABrKVsAroEUb0d
PuqYitbNjVy2lz2Xs6avmAfjPpgkAIDhe0dYp8tuRyOppRydZ6BaEB8/PKU47b7x/CdoPFDuaycO
V46Wfx9ibEkG1zz6AxwrA+H91g0JFcalFCQ/vNrB8qeEYKj+KsZvVPb0WzRbh5IIR05054yAATif
Pb2x0GQ1UdqSvtBqy1mqH38qJk3p80pf9r9XB/Pk71zhv7J3nPK3+jQFUYH0/qu1wsGlv32etD2B
3nVGILLjLoCEdEDXQ9cj3r5kVeU5mZVg8Zm1MkQcqni82iQhpbkPOYybV40nLwL/HirV6is5RRq0
UVDA+X+PWW5l5g5ImN5H6ty71izTu8Wf4EDjkdxbpmB8VEqkOxqdHWM8eYVdwHPfsDPAj808lP6H
5fNU6RpwwkThE3bH8ZE99S7pKXKOOXXZe6KbBMsJXs5D6QGoG2/TC96tKelAQtEvh5tXK3T6BtF1
CUnT8vqrQZnm9N0IN8XkD9gX6v6/XhZFgoWFGeqRbMfslfNkCl5ftT7tvXTg3pLv3kZMSkBrvHd/
tD3yyVMXrswjkJc71ibtI2H+yj0xtzPHKjxc5jLC6BqxU0O1jw7NP5QqS4IrlRcqjVeVOgzMJK3c
PkCo2vrhrIG9+BrU1bdhpBI6Nn2I1lM5g4gPj8fqkhCGXGmZCoxZNpqvrVzv8MxyZi5mpZVOvbfo
Wm1SZVHc9/6+t5wsmPLVeuzpMdZNktYxGzVVBTxtvkTgGhuW+mr/UmQEF+hskcM00x34oCIDMKaq
hbtDur4M/nvd5uZessAmNiRMlKs/A4MmAAGP9KfygqWrmWx2BN8jSQik5jnBPcrjZKKJ+cUhhjpO
zR7xP2YPITOkaeqN1diobEuAIQJaoOaq/T4BiOx+RyzMDAe9JTCwOTwfqAVB2vELMGb0V8N3W5w5
z9rxqK3fOC8bVWyZbw9+XRRtrmLsHoCjRiD/OWhBIJC1h2ske32osdKRMdY+zNy5yfAq8WrkGv7N
x344W5ZjdszwsiF/kvoy9iaYpCAoBLDanBNZ/DMTglafPLfdgd8rxS/ujRVF4v9VlpoHPRwzVBMc
dW3MehWnJO0LVXBt7m0ricJpJMYSrYtxfI6Od+DrCKF3Co9tk8zixyydlQiuHCGnuOjFVkqa4aeu
f0nEkTwpdxs2CWgXM3evxQpxzJPfhVLbAk7m96PQBZ6gbC3Jv7SO3mSRXyiifKA3lpMZoCoBvT9z
kVaWShOLVYQ/fyBWvRD/yS/42WBW5Mq41q+A1dVDTNHyzDeDW0dTSLXIhazXHR9W+4oFjn8N9Opc
seOWcItIE72i6GqAPdApZCCeJfD/lYgaRWqURZ8U2+f6n1QLrML+5qRsha2hqUehtHnPGVOZdc0V
aXflM1ROMJnJ1/lSgTf83fDjHNNEyB5T4sQvn1JRqDnMO0AwV4Z6Yl6rob1nO0kPmO71fQQTZbJ4
7wL4gjOpacVRmUs09dgxCR1WrFGhHOdcAWUWUxSLuRLNLjC/fTaTIKKaJav79FiBlpl8nt3Tgy0Q
ndk+ZubL4oDEakUyKjmPho0631zMx8t4ng20qfcDgEc8kwkx8Ai8+m5/8JJkCYER2PySN4y4JohY
R1IdOsda9yFNvXKA6j3ckTngKsCwsLTJ0m4AmJRohf3w/nfwYDYb1/wCqRD1hl6OQI5ddHCVOGGD
nteroGSvhtbcmYsWfqBcfeRXMKOqkn78ePkFfcF7VfxdGZsSx8FiJpnOk7Dl3emHjWOccwuy5yy2
vs3bysandqaqM0HuZ6OTWylw/9fGquQLlc5uJA+g52y8uR4QklxcOyBFx7bfFASq8qzJVwFkbYRf
uKHyTZqizrBsUYacRhFWkUJfMmZnnN6BwA4tOpOlBgf6BvkAefNrs1E/S+P5MlmXo8YxyeQ9ih3J
qXjblzk+J2u7bi+ah6PxAOHZnWdw5MmO4aWZEOjyetci1eh4S+Na3PKFur+6URGBnR0jad2cyivv
jHXUJLUPdiTPlA0mk6wcxRSEf3BkwPuaaiWq3cy1CnKQNFmHvW6cAlUqIT0LEMdiBTxPhwALrjEu
KGoTMgP3cJVhEOP0wX8PZE5XhSsTRSqa+HNcHSC5iYx1wX2wQSkxIytcJHpPGECq5J7mjfzOad6V
i2wUunKAuY0UhAYhCrza1IjGfnuhELuWMYR3DSaVnZOQwkTnPtxcbGmtYNzamcm2mh8t+Pa/3Yqi
YaCkiFTb/R0YxIHT4BdRvuxMMLbLOWZVLfxJ4TUoSjczwqeO4R6miatlfXpWFU02Wj69T2K0A/sB
yGN6gmd8tjAhkmFbWljtzxtZiQlsUjSHOVVPgInMEgCCIMl+SHmnboW0PdZztcAhn1wlv48XD+KW
6x27Dc0dWbsRnEp1EakCZR4cBOXHoVY6duvTLoQYwZ0itq/oy8aFN7X2+BrAWTfoeZfQZyJ42BNV
cxmxMH1WcIMnSnKpUj1579l6+5iJDc/xew1SfnI6L+x+6zxmFw/fCFKgCsym5nTIhbfX6XUo1Cm+
3oksq+k1mFn5/Scy9RReoAOZKW4uu7X/isKN9vQDsgAzXMmARhi9Tdg6thb5+mbBqEo5soK7F54v
EPPgs9WaVElGRLne/tdRw7WG19HMtn+pZCRLWJ6OSpQS5Jeypa4/Re91Fdvzu3yEt8kb50MM9r0d
LvJwkmI3AivGUHBh67h4rQdZpltmp2DXU/PJbsF+zft/d/0JRd1evxL41o1x/rSlNxCM+0a0tP51
bh7smiZAddbYl95Dpj33ooOXESjxymZnVZ9j4awo3mqk5C0sdKgheykoxf0jvQ9gkWL+z5tFPqMJ
naPgu8sva3D7ccNQvMl7FtnZxLUBISs8Q2XbKWSgt9fVPS4x74O1VfNdhykYvdW52x6fcCDODhWH
s9hEToi6AvB7kmTex3oYMrUUuB5Z/WLQZwmYf/7HGAlggGcRbDLxmrdKoJoFMIXCfAP/Rc41lx3n
jRXX3eLpJsHHcUbmT9dwcSN4DvUlTgUyjiKPhsYulXFiiFJeF5FwXIDKy0lXKsrq05CvHVM4T008
/uexNjv+wk2n/SsxBZoSS8V0x6PUYwK2nh9w8QIQBKps0DF+VURCDCQgYPiW2/5w/Szk0l5UtIwD
Jb4LYmtWilRNB/Z4vXhKUKCiceYMzMY5OEjU4wrE3RiXqsF1W0ccmFCa74E7lRic0nlYSRE02pjX
niab5ptKmo/xIJ4NeeK1g+9isgnG0qw+mG3kUEbrsRIC1O7DenaL6TCNiS0+Rv9sxRebg7lIyLqh
ZuFEXWMKjS0APcu9B2o9yDwDhVwyoJnwHdZ1+KJht4Bn/UXlp1GVXvKLc7t7U2QUlZBNO5y9ayp6
Fkwgs6g87WNgDFx5LpCHEmx6Oo8bzbxPXn5go2cmRpF/N9OnEPNMdM6dri2qaLaUris/Mpw5t8Yi
XO9FVlbmgkmrEDsRZcXoJFhvc8fvWSkFr7qlg19bh4vTQtsmPlLSfJ33UDoy8Nil4mixfPElS/5A
hz6RFfbU0ZsQNSltP5hPfmsnRTpCS9JhQ2XMbRCPUBaLck4spRAvL4HCNUvyANk3VIg3b4IVazpU
iljsgoK34LSPp7Ask+zuFrctOvAv+wIDO1lEKIpXwD2zrFwnzjuR4AVf8a0kDImiPPsTJzO5fowg
bHAvKiQqHh2a2CMqtldwKkJVNuEOZSnkM25/VxacSqClzyPRnYl/OQngLjVyRY4Aql4LijHHViZX
z94sU0Uq0dsXJNsU82KBf+hsTlooPiS/Hy0CFGb3EfF0D8l++BkzMgQVexcs8BeBWc3GdG2Up9Ko
Smafo+LChjHc5S4NgggGfwqzPh0d33fg+Vb/6AT6wLN6nQKAsRkC+WuVbuTwwzoJ3Ax0ykhYD8zC
1YVwdJ39EFYR3Vlw58vlzp2X/ecue7K260TAK+lXSsPKXADR3Prr1J0lg6mxjO3IdgC+NALu8yOH
3qAk6bmNabIT+y7znydeyKR37ab1zZBbfI0f8/eMPsk3fjW0+Cyg7Jc4wgDfOpJjBy37qlqZI898
FWVViOtOmDFKLxk9gs/yenJ+CMoAn1gLGTh2xhAL74MJZNllnj1w5aj81GS2yXESRKakPFdY8MZl
2XPpyLhxqBtGu1wHGQf1KpaSgOZymG/CB0+RWAZcjiOktMBeb/vDFJ4UcwBjL9GzqG2CCGfmFQnQ
jGHRCUDENCyypjP6csDfw/FdsJVO0KWCFIIz+VFN1PFAEZVmpHz9TpC/erePoUTJBuFxsOy6tzSu
aqW3L8Jb8Nx2OeYkqFVCreMIqZLv7A11P2aFjkzJfq7FhLkwX+J/yYXRlmEFiptC07FhAocZStTc
SPuvrwtRaX4JPjzGeChvRG2vaooZ70E2RQpQWYtZcOfFmtFQhQN7JOWNIFJ8yOkqQCwwEcdClqy8
FBDvT46FCVI5lA7sZrcai6llNITPcFSXM0Y9rAo1joDVYRb4WXCTx1mW9qBKT5t84b3pPWM83Fcr
6VdBEiZw0rNiRcecuZDqgywJERvDFY4qnfkQsZ89qgJDccXLBvg8CeHBJ4yogq7YakVcFc6t22WK
wajrBCl91i1YC1d72YurV/EqunbIsT1NcK0zqJTqYDLTLKXca5QTRe/y2CSAae6FWPZpxvMbyZDh
WQZ0ndIrIB4+emj/+tTheajGt+co+iN8rybHZuPbi/1roXl9uBscVgHkA0xo0BmzTrFk8JEidfTt
3SczaADlc02xgV07bBguOP6RjhqKrWxjtFpd7Cuw959H8Piv8CrHk9rWerdjf9qyPF9YnRdPvxf/
mw7lsW82UCO8PGCKoipmt5jU77TvODqVYclE2UEnRZMmU+6MwdhEEjQWd8cnURJYYbRS++dlytML
RKJ8T77J8JX1T4cK8akgpw4WSqORJBHf/m7K/t/DVG21Y3JhQDdP2d+jjHtRlp/T5aqogMNMqTg1
B00wg4sVGONwtOxVyamoQoMUTSfHaGQ94R2fkjDJ+85+KeIr/2/j8Z7z9vsZ2VSDOZusLGTCI697
FPcBU43jAEzKTz0sHXq1V/cj2qDDAtbcV4hLyrDLvzSHcihufJcBUnISrCeFsZISuLoittVUHCNX
f8E1d5tbqVb6KegS7lGZsVKPe0Zyc8YqShcVXmLVIc1Y/s/IY4eJ3RBdIEYi4SsWcIld6k30016F
nhVOQ62mSIs+Y25jhV07PotabqkhMwtQ/8QYtsmjMIit3K4kf6NTBas2zNzWGKYj90YnhruEQdft
yxBYhsuE2gkmozbphaT4K4/AhfpRuWJnA4/DpUEdf3ld9PolC/n0RUJ4rDDOFc4US90NPFyhKZ37
VIZAoAciyT1SFUBHh4BVDqj/CI8NU1G3+a4TvxBzeTNCWH7qGjId1qm0QkHE2iIe2p2oFA47iL9k
nhM9D7zisMgH9IpjsDooB0TwBrujJxhf4up9eFSjeA+7nc26I+MdUMYF16HPmOSCpT/K8kqoo66z
we4VHWgtlOcaV7Z0gvlWwt3sNWmN3GNvtwoKvM10ojSnSX7XPvStMgkz1rvgnqzr55h/sKMKNsY1
+Iu9YMA/F89d2tjrRQ4LAWZZDN9LSzMRr2J54JIrXWarkXhE+VFCRexUKMZAig98rKHr/Ym2kM9B
KqkX3s195i/iEDkYJXw63nyl393WjfSfhisJub9xhD3GzQqI9HYixObgnce3WkWrjWOmOjZIC815
FUVkv3MyKXdLBvtgeKVPeOKN5LNET/FWPvcf0wTe9OzlsYFDe2id28T62MjKXZW2OnqRQhAbdos3
eQ03mH2OFnHp7T8n0EuSqu9LnTkcpmpdiobVd59eLeH0Vu2vpxpOivZIP1Ag8hixIty3GPdoIDz9
LPqMyHbl2XsLQgOBcf/7taUlMD0bEsr4GD64/9P9d5R5ZG0N/ILiusvuVwMVjaFK55PNSUwFjpHM
9f4NfEvhYH48ZtfayGJsbngsYZ3xufsrhVQ2p5qK9VvOrELQXWVIR7V4+jkrPNoWDz7VLDQyVukc
GQPkBK3XcH1thqwQBkVs3BGXYY3mWxy+FvuY2C+PP5tiBsyMdhQ+skt37/VSIRWAaQ/QtwrFXzxx
FUmUcuXa5Hw7+v4JFJfCDtBpSaaNf+T/7GQ46d1+u8Tc3SyZVeZRe5dC9zxroxXMzDXZoUS7o9SU
J5xodgAApBdY4eS5ANOHwnT+bS6VwX9i0jR5bIA1Xfmi+p+ZYRTPoCJtPTKG5XrV4Ls+PY46UDYT
+o9obO7mVVJr4bmlRl3f41XZ943jMSWnt6D47QkUjA6RgNm3z9WyTEbvpS4btgZxwwO/5fai/klS
syI3OVncqO++n4H6ri5a3yekhfc/W6POX64Uw+gQWVRPRfSfKUyymF9NDdv2EHdRxVtuvV7x2Bwp
5Fyhh8e+bhSuEY1AGlHePNOyZgpvTqJke0sMppy2DlLkUecmeCWW35379QRrECv0zqtKPvT7/wi2
Oi5ySSaTyq6zD2P488h6kya8FJr1M8/GiaBDZw+3/1BsnsGPmePjNkqyUxGgYTzcy48HfVEfM88z
FzmyViu7vyaFP/rOpDjOWYHrztH33CRnHoYEtI4GIbuINbt+ppz01YJrbJWOx6D4jEfdw1f2euQE
a5dqAwC7P1UKFjr1aka8e4mdtu6Udns57vNAcF4SaUM9xUzprsk5w88VvU3+Z9IFDyRYze8ly753
7M2hx5b00oSlTO9nHVDDsRx8ldOUuiZpyjeM21tucsc/d61m0u8cY0GxSJbsCQTBNjlmrSEZuNOA
IFkY/hjo+zLCM/e/29DuCsWwMVGiLNoahfB7btw48CUmWp5zwcc0yW50HyuyvTPueuCzyLBCSuJ6
D6WRHmzqAFv7kyR0NaGrNZ7gpuLI7G32WFPNfZG409bMUOuMeT0t6V9LGzEF09Lk9nYS5iHFX3eu
udYrhyVyfruayeYKhEKPcB6QZNjtnOvTzJR7QO38LuysysvCl4KSgGenPLu2BiE6p1htkscdinZo
LcRMllIDIRVvzxcP+J2HMjdlf6tU2MGOWcPFmCvh3LXsH12zC6K0UDGULUkIF176J+h9oAoT+N0k
v7dKpMC+ClX8n6uy55JWAvUljAdMiLgDf2+Q8sBKzsikRxU03vF/D0F5KDcZoYraH6rzlpe2Nzjp
Xj0OOvTwA61GJF+kxEM4xBUM+C1bpE+BoL6Tx6CIjIwkWnrZ2LLqqZ3V7Fq6w2jVvwGJfdn6MxOa
RZAe3hen404TR5sRGCHL9s2QGFzIvnNTyVU2XazWRSZYvg+a8wGAYmU55V8BnNwXYqC/xM+9PFz6
3l90kiJp2KeXjLyVzTKltn53R6lApJJUNEnJw58DVByWa4jEwockeFnbR8afEv8s1RlJjdVQ8Yrs
eqKmM/lM46TmphRuYROkCJELx1r7z1OAwLo4BqtAkRxlZAo5xdvXBbEsr95K7vxkjS79/7moT4TO
d8nCIQonqZzTomsDfdHuRWfgjiUKtrVNyOeqNqnDuvYQe8oGlZv34Y5rBv5Yl/w5yCCQqQDtuxeZ
ruWiEMvNJ6DkJc367Ng4ox4x3Ez8jHfRKQjxn3sfyaBoJNMZrwgBhobZUy17BVspwvFzv0dV00Wv
z5/V32arhN/XDTvAGEjziBqpk3TFXV+e5YR9aunUUnyuAvlIWpTahsZZdG93XkiJ7yPKx6FNXyTE
53wUqJ45l1OlpMkM4t1lbGyc/yvP0VcyGwBppCGPvNveEBQTcLlefV4FM87C8U9zWIOvobwYzMdE
zjTYdokH7LrqwY6O5SxLTyZ36DYwax/pw0zis3eheTT28iv6IZzX5gB/SM6JCu2xyRriMZorGLGA
OXGMnpuMUxY9MxTnNVBBL73J18YDsTJNPvMIX5Np+MqGLnt8cjteQYGA7LSEnqD6OJbaIkmCA6vo
hpyDgPScZCPP5jsP2TqGYqWDolNbNwWmepkfGZ2EnVYkyjFeFf62d//QEhn8nUobRhVXb6dCoWQc
wnV8InEY/GSv/mlsIMmMEiK+LdgPpkClrpMUUBthnmgOGvdpkRjXBFeovK5+tupjpfD61Rj61Y36
kk8qcmVGehaB1wfHE4rPRGSqVY0AepisryptdsaImj7s0fmQ0iSmdz6FKLs2+RVUlYKjW/mv4JJA
NUN5kN5kTDcGMlR3MTt0+GAWL5kl46ucb7c3577jV/Xwbe2Kop0CAL0qHHca12SeCAAnu1ruMnsO
YXkk8JbLlBkhG2HvOgnimHufVPFUoffk5yIqDS+Bi2QgIQFObDg8jhCa3R4mA3iw1vvUvXXpMwrv
bU1P1hhKu6osbzj5YxHrKhifDo33SY9UlnfhFBQm9zvE5t3+i8OzYAbwQyakrmYUdZloHALq6+oZ
1GvK3kCN5lGMJpxtCz4owAyZaX7Ykwsbuxloku/ezcf6OQwX4baqbUcbaKSzlCsOI5clDvvc3PoH
m20gdV9r7yEgYaY1cXRbhlL02hotXoX6KC9iU6n9rf3GgBqVLzvFNa3EvEb0J31NCv8iFRjeKaz2
srRhPmC1QmKaU8FaoI6yqdSDy6KNBJawj1nCIidIzQaemZFossjKBDBz//lcS3DPhdwl45Coise0
/EAVXDtaZBCJxhkHbqrBQzjQkN+yEwWfHc+FNtpnc4tqdL8TqLUk3YkIiK0TZ9xCai+FgyQP+6Tf
c4zbQ2FCOxmpMk8bX8fCseHLXqEv6KjJcmcKFRnn5T3O72db3zvXdWrU+GspJIdgc27zJk1u/cl4
nTAFWUMtx3W60LRw/2sZxNt5KZmqGTcfp3gYFlcFuV2iXlNhEIjfO3XcOhh5oNpurhR30Q65gvWv
wqxlsX0ieDW8qoCbEWsPpkL5FaW/Pu8QM0jKLE5gRi6qLXXOroJf7XI8VTi+x0l+iPgjliqKuLC9
coi+l66wjrWjCR6urbTUgVk/GkoZOzeZ+u3cVf4Q8DrnCbu+8axMLTRh3lTjJJCciacyetEYEiAq
u5pfUDbGMzN8lJvNg0/dX/KRWm5eGX/axdnPrxPzlYJthujZKXrPzE/TKjmz0nKEp/6/5CvP9KVm
dN8ILka8ovIryZGWEvJU7Fi6CLFha+HRh23DmPVbEdBPdoikdBGsBzJrDzs455biZL1X2gohpJkl
DwSAxoqNSmt1fGb5M7LgC46TsRLrkNnG4uIipBM4XTwsJZJVex1mj+iRfXqUO5oox26itp24W7CJ
7iLN/91ajz94+ZSfXxUsXxz9huf1l9SeYmfLtcYsSy+9WcI/YjzrPxvLxLz9UDP7mWoREsp6/KRw
i5v86r0HusX6cYPixCd1ib3631dJ2krc4Cx3/pIF8kO+9/VgO8GRORXxwTRimpumfuSIaz/AQ9fV
m1BnHouKyqQiQBoBBl4Ch226P9RfDcTJQGPAf9QeNy/JJoOWdPv0OSnb4JqQbv+QcVhRtqrVGAWg
zQeyE1rS2J93kkdgdqxTkkp/L5oK/ziYfN81g7cVHYjlnw6FhyBqHGKR5zzqCBTEt0cHA3GFykiO
XJ2odDO7DNeDMx/rZ1psbsVxIoACAWj2QKFRurOrL7kGU0o6ruphhlKLaWws4k7Skam+eiQ7Guvd
pkdOEg6K9IOLorim47IPGOEvf7A1Cx8UBRf8gNEq6vLTorNFwQLYohUWsF335dVRJTblu0Asg+G/
Lu8/C6/7T6D6P63awNq+14RodiNgZefc9NFtbRpkhG/A2AiaFsvk510FeIYbbsFjRYfdidkPlD52
/hOhvPGzwG9v0vmzTbd8FMCfw0m84A5nccXazljfLCfdQBcEyi6qsWNUiKUcCcRVYHV4c7yaXHjL
vXjMGPzPjkO57FEBaxNKU0r3wHshrYNkkxmvepqPj2cNgmugZeDji+f1n/ZEKuUscm5XqUBzP94Q
xEr4vcZPzGwBs12f5bWyOnNNtUJ0AYq20oxcFtxa185gUUzDbpt6I73qLZrsc6jY0Fg+3iOU9nsw
CEUW0bD9/G0EkonzGSmSwM0SoyD5ofwrj77RKaObIwtXE0v1MOD3G10PfzMq4Jv16BG6pInfT0i8
67A6y7NKn/LR/I3ZDMjdrmZcuZL7lLf2uR/DUwZar3y1ZyUOtQXruMBRW10JdA+Sg3tVCIZBAWbz
smHbWsADDsUxppVc5zW5qCKLTqySVKZKdGPCZ173zdlVLgDoAiWhlPk0WCBgRb4sXoKUoTCzfQiY
DGe/bPb+CnTevQGA7u5dJU9jHPylgaGEtZEdP6Q8sEaFhEK/hOokjfi97eJxs2hNDff8qooh9/vj
pe9szQJO7wg0obimdkP8jeadcUulG4slCU5NReKCy0g2l0GdanOHgWXadsr9qyz2cd8Q8zI+WBTe
XeC+Fa3iNyrcPwYDdhww5iH9J9a17G7utVYom8m2KNbsGcDh/WqFBpAVutpE0WP28FxaJuksLX8k
tMBiJphRL2LKQZOovRyN9MsGhq0RHZHHXD9l39A3Wky7GjvuNep3ukZrnJBwrCfnndDxnLAGtW2A
h9jVx19hGHqmHVCk7KYtrXNBzpnxliuMTPYqTnsTfF2WpHsPVdZNdqXgVKbuFTBER5U0G3tkGaTH
/qHaAk0VIS4boSqq8j3YBzXMWEsExwuHSJVK6aGqXIkTgIBYjzMngPeh1/CQcn8Veht58atp7zf0
gf0nthldLiWTRAkHCLtON6u1o3IOsdA6abQT2eMbNq+GeTilAWcJVFhv2btiiLnbQF0SVvl5nkUM
DZJgvQGuDdI3DvWa+8gsO/GspkfiC+JvRaCvzTcx2leuNaGM4pJITK26ofq2qhIqtV/Bn9iJj77q
0ILdXMqGh8X6MF3uI2Q5gbr/XNb+syMeuE6FdOVwA49Dkmj/XVC9wbPYmHYuD/OK27kQVHPiz/jq
f3HJJ3F7vrpOmVXvdpPhoY2w7EmHqcQha1TCoI/d9ynou+2W7GE2AXKGAkkHyi5AzH7jBQKp68IS
ges+TpP6lBzVvR24AyquQ7fgPGTXyEtaBaP0zKpe7Y2NyWiq96w/fGsZLPil9kuNtoE6V4Mr8y01
13s0qlqIDGaGC9VKBGJJ92JyvszkbiEFui6fo8ilz6LWWDu27LLpxFXMYr+S2Q4Qu3fiLZuNJqA7
2hmuHDZnEdSkadNwV56QDELX5TBEJQTvpmHWM0IqwSQxVjIssSKDfMP9RINijfSxytK32Hj4UnF0
dvDimEcczIGgjqrjdSYQ6sZJiLoGG+HcY995erjEUhW4kp5p1nx9pR2I/tE32PGw43DbMISL078X
R88TNQWgBrpeaWZ4u2SOSiswYgZjJkcpU7DzwmfBO5y8qxW+BG4GGY27jhR4APAy5Yqqo+RHqybp
rvOroPEbYNxQyHSJ5JuyN7aRvHkwh/c9eud1f06foz7n6+tPWw6Cqn71P018VoubQZ1JzcCKgY+a
Ema+IX1WkPOQtaQ/GonTfSLe0NtKhIuvIgldEcQMeACEys/06w3ihAPSN4OAHOdltuq4oTmKCFwp
q0s68BZmVrBRVCf2p9dninL/Me1kVgxLgGlxEXO7YPHMD3h5LrcJ4ect7Kps08n2kHCsVrqrNV+S
F9zgSk12gWwoIyLM50D+5NC2V2dVR/1UefDOPWfAScddcI5FX3uv1xjvMkgH7rvczwPM8PlzyXDY
RyV1dRPjnwWzRbvrcs/rKE8hVnRucUe4I2xgzNKl60Z9s2AZJF6s5mEqF+WURgcpuF9s77ZE/Bwn
aFEWhGkFRBr/TieyZbAB7L71toq9gvbkOxKK4nk5HCAJg5CBT2V8fqK1hqr2Euhbx8cpj4sz6ax7
4fxkoMa2r/DN7O3CeUp+8MAjhpHzay8EpiH2O6/vz0eJdVcDB1PIPQ4KQdIkleYPSKZGSdnao3cg
nKEpNVSM+SkW9WO/qzupFPgcJsOqzWNElOuo6cP3OkvDPtZx2/NZY/PwE2OAzso/ubgaGagYDnm5
uBj3G3vLpv1CZ0IeSb55ke5Jm/uvh6rlG/UxeNJ0fNcy3NKHFa4ONfzgRbGfbS9QnM1lP7iuNdwk
yJaFMepe+2a9E7W3tPrbZ9oCYHGgvXGYzbYpFhLH2mpJh+rbXxWaVHg8E4aZ4fyD57GxiqfMUTDm
A5427Fd5OxxFsUroEeoyzkqijIn16dVHs4h0Js12bFbJxPRZ8wh0glJiXs/x0oMBoPI0tamINLbs
7tLDq5iNmIDcd1Z4s4LivjxJ+RA/vDpizMmVXO8RFbtpmNSGyoaywJs2WdI5gEW0sXQ59N297l5B
HCcDokDufmxsV5dQF/WItZoBNfG0d1rIWQMQajid3P+6Xm74S16pgXS+msCG2XrDtAQvI/BToR4H
bQnic0pej0Ey7d+tcQ0mtDY308Avkp8SZw/a7o2/kpmaX97Xda9h6DUoi+O7upyGIpGP/gHFTWDl
LPEyhlWe0KgYoQ7CqizBBEqtn0E2EMiOtIHxcbHRHgmS7G7kRfBlA3sRriHYV4IauIw9OCI+dZx3
tcPqzyuoaSckPVkvwGsMiCfllfsN1ZpkzcypB0oWjT7ydbZKRaiWX6NDHpb6Fk/YLMrXvTHz/2ib
RcxKXAdq2WCoEdX5MCkFoYI3ebjesotR6StDXtoc1YvEtAFjyl/9v3X+8oehbvElacMVMCQgIbG3
RWEM09JPrfj5Ly1PkculL/fsZfkjYTSePJ+D+HbK1qorGMBGGBSZwEJzzwxmIYzXCcr/x7I9ree8
jDmQ2W2/kTQwT+dtbBF3/Irr0SNOm+KUB1dp0cVE3CFxqMEAPQjKRVlTYLi6qCMQW9p/keUD3yLC
PDQkmJ2w4tYFkV1GqUQYChqCPakET7fHPlYFA2n9cLlFoBjQ+GeuSgs28wxFa3IXWaGMHV/XlKvh
7+Pg/o5PvQpD5gWB/id/DU5klQGW7FJFHsdEJtn6IQAxozeBcSWEW60dZh0eWhOZJzcYG9eWdM/x
W3OBzQ7fMFetE0lDV3f6EaGz8Drcv1grJZJrrb9bZ8pC0xeD2ydjDNSFHJfWCPZpI9JUXyBiooGg
S5AVq4UeE+666H0uMf11VWW3faWTtIbEvuDtyHZczwwmvptwtINmLtb+Gv3s9FqfYeek4uDFS1NB
999GYHPWpZF/aSBtOukD+Y9F0ROwXus0CaWC2qw7DKSfq4dRATClOjbCq3TLvu8iMMF8bNQkqhkG
sTLaONVj8DzMbPVVwwXWirQrBfZDShf+tO78oui8aM323f6z+Oqt2urP/zI6DG6dh856QtPYjtJN
3FLI8jgHkgSJnoACZE1WZn0kMcPUFgqoLYdIgIKzIgIvloYxqb9rHvTVa5GpcvS/G1TWJLCOp52z
y4FZPA2owTXgFkdsjEiz6AUfDE0cf9SUc//IeBNKXAxcgM49nbeAsXCD8OwXVtE7K2UsquOeltEI
V+8JK+O18xgnFZrvZmd3v3u79oDzUIeAMw8B7AWkUzWen6D3jw4HoxsfGmY4IY6LQyl4DGqpXIqP
gT5RtGeyZ68MViZEON+HoKfUQxRwbOC8YGGUf1uUvljd7VStOFzWrl8CK8BRYT29vv8gce/rmxG5
Gw+xlVvx6I3Z2qyuzg1hcNHxHnkzfPPtf6bFWceP1O534QJQqOxNEsTuaR73hoKqAcfMC96/oT38
3iBHScOjutLVkBP5y2oNc/6F7Pqz3KIG3Tm7lof5ymHtCNMf9OmPGk5K2MZTKag6gD1rkAILGf+5
Qzu74jCq6SMA1u7pQVSQWMrj4KHFEvg7Knt7EdIRVKa7t11srnp2D0B6CuevY6qaPkr3l6CBE+BY
a1NjpqPkIcRKIcojj1hNczoOUZG1Ha00zYpaxjCsp4ED6yR/68obCbIBR4REz+vSeqWnJooyuwTe
1ryqn18Iyt9L83U0vOk2OcYVMvH5YKqgi4oezxQ0HV7JLVKLygiKjqU5EkihCuHjs1CDSIoSRTxw
1mYCBMLAjyk/N9MunOPctiYHQX7f82qAWHXD24aP/+9FMGMS46QyS2JL7oSCqiaxXRIThQ0OOwdx
FGF0wfZe4VKOyMMIYueZer7AxVBRPS7psbDFqAY2T+fm4dkKbKXos8eA5fEdd3jRis3iawwxjkcm
bVZ1LRagwiu59iYTh5XhFSkCCI0nz60Rv/V77sstAI0Dk9oUH2nCSZI80XZqNQzxJEELBSLGMSPW
2JUvFY18IqW8F/5r3591xiUEEklvoZoS2IMLNM8wSTX3WDyFCmqySreXJqzFul08l39iBHw2etKv
NOrvwGGeWRtbZo51e48BiQ2SBSrOh7flFklRvJu8feeRbIM/90ZRvWwfdipXSwUrjZXl8oP4tb6K
qnQchVcu+u33V/xFJ42jrbb4eaes/ceC0BoMOnAw6Dbaq2gEJiHmM9EFpyTBO3lqHN3p+bFAxMCD
3buSbqWBojFQphZq/AQddLqZSW5etYE1M9MDh/n/CzjuI6L/L3F6VHvy1UxCSH/Ng4rZhTi3464j
6Sdt9Mhz9PrJrgceBFWizcu2eoC48RlnpW9VXJRN6Sg2sZr9VODTfQYoGtRcUxHEQf1tddq5YqZG
KeV9Jo5YIkY6ZvbXVK+MA9oICGJxFGc3nwCkx6UtZRygYwJiLRI7+Tg3uTcoPVo2ymTF68PikaZs
s5YAO7xruOkTm0/xchtdhpgHmVh6I8GKveOMhrc8o/kad1RI47wth/Ttlh+Nlds5s7FWKOoriB1A
VZWEoAiy41qCv0MAYECs+7qm/5by+Q8tOO0TV1X1/cMnNdLdarLdPSh9QPsw1ylgT4/z/3Fi9/3H
1uPexxSGeuR4Aottjbg1/dcnMfkgI+/eF8wN8qicIs+WXjfPs0x3RG0qiidr+d0zTxQlIusOipql
LX7ERp6zp88wZqxk48b2dPMoTVRZWRzdCXnHcTJpbHs44BWDEW3okqBZlQC3dPpS5V9VrN51haF6
IAwhr6P2vnnxNKEXlgo0OFCr6fkq2oYWUyn6O0ajnx8WaeJ6fmF86aEtwfYHr+VqQWAvHGWTHSgW
B9IImsUVOAtlmIxvEAK2BYYYcEDX5g5y0akKu/O/ziC4Nr7Wtojh2c3kN0DqocHitDazx4xcKD9K
1MtmoJuY/Ca+turpOSA2A6fiYmNGxSHszgQHzrTIsRyggXBs0TqydqdtlEALT5ZeHNu0hHUAT+1f
WilnSUA9/mK0vYCDze7dTifeFgWko5Hf7ifFP9jvyzLuCqVGzzdpOL4XDqpyqu04SoyeHLYcYVBP
1dTIYrZimhzrkikC7tLSfXq86nSSu9e7pVlU/op0e1JyqLeJfaB8i0MMsyuhOLyeZPyHhknphAQ2
lDkz7GkRrAc2SLFImkYT0j/6iJiVg1/zS9rc/OdKl1bUQR83XCmptZtK/23yY2oVpXhoaqkMq3Ve
soUUY9K0MCKrHKwnhOKHjN1Pd5HbzczWeZcZfZj96wEsk34MZWJW+peipKYWExihlTp0k+3Qnb69
V2I4m6NnXRCOcKXTMMhxgfxsLTV/b1iopx65ooe4ITg757/VFcs0IUtaswtzkRdXXeKwX9FeIU2d
VhY7L/sjj/IYPTnpH51RpfXLOdeI/oBLw4RlYACnPifXF+4l+p7iuA19l/WzL6oUHVJpXmmPr09n
nbWmpQqS26Ovvb7L2hOHT5bwyljAu3WBn0b3IyeyN3oIOUOkF9Gh5TwA2G9tBllqrP2n//xs28tV
r4gNDHpYcncjIMHk0h7+0BpT4GMkfeoRsUWBhInRnV2oDjGOzjRxc1FYjcoiTyKSiy7GkLHbbV7+
KO2p2sH9Cdg27iAAGHBv5RPll9Q/PcwA3X73Sp0mTcyyUaI0LMdUbBm2QiBbT3cMZIZzGo9vyRle
ZW7jarYdhqi25QrbCepXlsoXMM2dhZMrffa6k50ktM07XCD12hjk4r/o9cROh7jLZFXQqIu+e9xe
aKx94hczizxh42bj/YdJSNbTpdum2kU9NYtFv0hV6xzUPDcztBEUSza83jWq5qF/WdB0r6uvQTw/
G3uDH1SjjhbuiDfAemARpra5xK0WEkDlipdaPL0cKpxMbMBAsEqiwHE+pFtBMdXAlT4Z4LnKm0/B
406dHcXlgmgxd7Sk7O2/c7+M0xSoaXnxA7BQGIQTH8tVog5TgsPd6AYo908neNrZ8ghLbgKGm5eA
G/kaUDdBHDGBeU/aqpFO6H+adBYXWq1ZwhVnuQmZWamHfsonscD/q3UyWexRtiSRz+rqWuBBjUNG
ODARZGWySTdrxB7MSFGEEtrVwrnKloXzevP/Fhxoxw8N3zafBRjZ8cmdwbpQQ4nqr/jM0NRDbWUg
MCY/8pb29BSkdvpIinfObPpPRkGZq5UStXjiXuWMC4gjZi6MZwipGFkaMFI0Aio9rW31isMbiZBS
Evnp5tUBBtrj/sjrA+DahJEekCgabUftyMD/AYfpM93/mtnWxKktlZL30skonQtqyXFbTSztB/s2
D+oRqHfupjYRAOwqZDLcBFZp0p0jF6r9T5BaWr2qg0Ci5moSoX0iLeSomX1z46W5T369jUb0Wss3
fodNwPQi/RCDrneEp1K9Jx629aYQUyuOpRlswu9klhQXpBLKTO6GyEwsnX1uEoFbEh9jGgVNIg7A
v7szqkiMj7jVz8FWCiPPPlJ/bPd93Y3XiSfXX7LqK26S18A8dgr54ks83vayRdgiwsJ7jK/sSOk8
lLbhyNIyJaCgajXCD+Cf5PSJGbnMD3i/rp4SNs/vpXWTATo+GsRWLUE6Oicy6E3mMAWcQIvG7JXV
Vc4mia8P1TB4UpXy8FGG6QnSsiKpc8opJpL35TKImmfqX+3HzEvrr8LpUJn6Q6wwSV+WltYCg4H/
5UPL1ftQcrQ7dijYqQQ3Dphbt8UieWe8z/gQ8RuaDPjB+di8+mnhIilOqKcukMj/6EObXg3JIV9M
ZI77Ew+r23bfbKdtcfVnAewUnytvKp8ISh72oZ3rLeBm1u+ukoWS3n+mJYnZdr2g9R72BnM4cGkU
H5eQ8d2LAhwQAtYHqaOQb/h3Oz62dUkfDj0rS0DP/8vqDXWOBhOfsFHvjVZtdjHWUYgMj0i+QhGo
PSbGmIapTCEPYAqgHpXLERG2M6w/82Nf0Jmum3OUYZoDtVYgR+5tw80hdYTC51Cko9BrADTqOWxH
kGf0ags7Uh5EGnUcwiGuxGGKFDKfKWmAnXWN19Wj7ZgLRS4DKUPa2MWMVZ3JCtKzXoOt2FHmr8nl
abXEUP0lCdBrRfXXLftOsjQuWu//ZM4AMZ30P5OgorldlboTZ8/ggdVz4Cf7oNaZ4QAiKMnMTIfX
0SmSRfHlohSiFkF6zQPgJcQDlthx0iK+X0IKtn0ooNtR16yEN496UqhxVeC7wtlvns5n83Tb40B7
O83r9GJAvVJXfydoleVSLpkM0CggInav1BU8ddE694+5xq/ad/P5qIpARJewfdb9vqlFLBb5MJGE
Caua4OxbzIw9vMRl5ADcFx93tMXmcBBZdwiH5VX1ZxQuKgRFGiwkAutAMNzQTgoQifRyIi+V5akB
3K6giIY2KJ15GaU7mk5ayR6rRKXJ42nJy4o7oc7a5awOVLmPGu0wpANIkv/uyImw/4NP5qyeW+PZ
3X0anKSO6w8Q2p272wV2YcGAzs6I80v0wgrhNFS53vZmQ4kiIqza1LKa+wuiH0N7hLq1DIcMY8d5
prexpwcGp+kMpozXftl56alSp3V19U2Vmy5SnmQdp5T+soQzK3t4nb5Pxqaav1Px/c8FcZ+lt1xe
DOtGoNL4bMbbVvx7NC9UA6lY+XveMCkOf9JGEY+kBqPrpI7Nv+L4tL+3rHtvXScNBPN1GrQeq0td
LRcy7MFCIwMcCBAaWOQ4bsJQDE+T3brAhTx7NQiKZLDTB9i+IJJePoAqIo63x698sRAoMNhTFvSo
FFo/F7l5NP34MULl42Edi0Uzk3+JPNQs6En67Xs1teORSjG8Vnrljv1JuUVcFtzthbJqqKQuBciN
uP6tzGNmf0L2AvESNVUlWkdxyHiudSEz/PeHfj2Xj4IM6w8IAZvQ2QOKZbUA5mB1xkuebrOIr6vx
FbQ5FAzWcHxPA4QVhsfRAwQPz/Z08jTw99sMmUuCT3r/V6cmNZwf+sth38nu3sWG/W6qTsu1wjtW
Aq//K+FGsnhFFmSjoqgg2AufC3DHrD4qKpJL20qCcr8GPxMSC4kKyIoGa5FKdEaOKr12Gd774G9B
oUjDF54BkHrKZeSudCFz0STR6ndiBLpZ77dfM4Xq1B5IL7st93vN+i/GO9Cv3CYYb8hrCohqO5xk
lKV8CGt3XNzuq02T8srUsCWUlVDS01UYqmFWsQmGFMGps6N1zTfB2MtinIWypt92PQp9VpUl9c9W
Miwe5sn8UAxCbm98UvbgkNEcr5VLPEkdxwdgYvirxx4cyqTykDWNSVyfLtsjr9sM7GRp21umtCBz
Y1PcQENsVgoU9+veKSvYiIsIUV0h1vsUJRuNObuwGcZzMZHCOWnJSH1lsaMpGhN8Yy174HwJCHCN
AHdfJ/wfkqKq48rV0bWLsmMDyjY6ATuu5oqB2enu5SazN71crY9InEiqKVCfyyJjUYGD7KCWCEhM
cmkLFlI1gUNnP77zmniDstsbzMmnswmC+GRVk6QdvJOlPcJ/cmuFElUsbES5MIUsWabvLu2x0Q1i
KgFCR+n6b5e1SBKQiodYtpPi97B+X8NaM3Kc/cp4u6ZHP1jwJ19KO2VdWm+hScx7ZCYwpwO1Skfl
LjC40hBBD9lTHjq2okShN0NwnKH6iErkyGZ2/nM9yDsxCdiT75jVS6vU45e4opU8GF9Z
`protect end_protected
