// BLH dynamic attribute configuration look-up table addresses
//
// Build Summary:
//    Built By:     mk_defines_vh 3.0001
//    Built On:     Tue Apr 16 13:43:06 2013
//    Bundle:       MMCME3
//    Architecture: olympus
//    Snapshot Dir: /tmp/JCf4HQIBFW
// Environment Variables:
//    XILENV="/build/xcoxfndry/P/env/"
//    MYXILENV=""
//

`ifdef B_MMCME3_ADV_DEFINES_VH
`else
`define B_MMCME3_ADV_DEFINES_VH

// Look-up table parameters
//

`define MMCME3_ADV_ADDR_N  57
`define MMCME3_ADV_ADDR_SZ 32
`define MMCME3_ADV_DATA_SZ 88

// Attribute addresses
//

`define MMCME3_ADV__BANDWIDTH   	32'h0000	// Type=STRING; Values=OPTIMIZED,HIGH,LOW
`define MMCME3_ADV__BANDWIDTH_SZ	72

`define MMCME3_ADV__CLKFBOUT_MULT_F   	32'h0001	// Type=FLOAT; Min=2.000, Max=64.000
`define MMCME3_ADV__CLKFBOUT_MULT_F_SZ	64

`define MMCME3_ADV__CLKFBOUT_PHASE   	32'h0002	// Type=FLOAT; Min=-360.000, Max=360.000
`define MMCME3_ADV__CLKFBOUT_PHASE_SZ	64

`define MMCME3_ADV__CLKFBOUT_USE_FINE_PS   	32'h0003	// Type=BOOLSTRING; Values=FALSE,TRUE
`define MMCME3_ADV__CLKFBOUT_USE_FINE_PS_SZ	40

`define MMCME3_ADV__CLKIN1_PERIOD   	32'h0004	// Type=FLOAT; Min=0.000, Max=100.000
`define MMCME3_ADV__CLKIN1_PERIOD_SZ	64

`define MMCME3_ADV__CLKIN2_PERIOD   	32'h0005	// Type=FLOAT; Min=0.000, Max=100.000
`define MMCME3_ADV__CLKIN2_PERIOD_SZ	64

`define MMCME3_ADV__CLKIN_FREQ_MAX   	32'h0006	// Type=FLOAT; Min=800.000, Max=1066.000
`define MMCME3_ADV__CLKIN_FREQ_MAX_SZ	64

`define MMCME3_ADV__CLKIN_FREQ_MIN   	32'h0007	// Type=FLOAT; Min=10.000, Max=10.000
`define MMCME3_ADV__CLKIN_FREQ_MIN_SZ	64

`define MMCME3_ADV__CLKOUT0_DIVIDE_F   	32'h0008	// Type=FLOAT; Min=1.000, Max=128.000
`define MMCME3_ADV__CLKOUT0_DIVIDE_F_SZ	64

`define MMCME3_ADV__CLKOUT0_DUTY_CYCLE   	32'h0009	// Type=FLOAT; Min=0.001, Max=0.999
`define MMCME3_ADV__CLKOUT0_DUTY_CYCLE_SZ	64

`define MMCME3_ADV__CLKOUT0_PHASE   	32'h000a	// Type=FLOAT; Min=-360.000, Max=360.000
`define MMCME3_ADV__CLKOUT0_PHASE_SZ	64

`define MMCME3_ADV__CLKOUT0_USE_FINE_PS   	32'h000b	// Type=BOOLSTRING; Values=FALSE,TRUE
`define MMCME3_ADV__CLKOUT0_USE_FINE_PS_SZ	40

`define MMCME3_ADV__CLKOUT1_DIVIDE   	32'h000c	// Type=DECIMAL; Min=1, Max=128
`define MMCME3_ADV__CLKOUT1_DIVIDE_SZ	32

`define MMCME3_ADV__CLKOUT1_DUTY_CYCLE   	32'h000d	// Type=FLOAT; Min=0.001, Max=0.999
`define MMCME3_ADV__CLKOUT1_DUTY_CYCLE_SZ	64

`define MMCME3_ADV__CLKOUT1_PHASE   	32'h000e	// Type=FLOAT; Min=-360.000, Max=360.000
`define MMCME3_ADV__CLKOUT1_PHASE_SZ	64

`define MMCME3_ADV__CLKOUT1_USE_FINE_PS   	32'h000f	// Type=BOOLSTRING; Values=FALSE,TRUE
`define MMCME3_ADV__CLKOUT1_USE_FINE_PS_SZ	40

`define MMCME3_ADV__CLKOUT2_DIVIDE   	32'h0010	// Type=DECIMAL; Min=1, Max=128
`define MMCME3_ADV__CLKOUT2_DIVIDE_SZ	32

`define MMCME3_ADV__CLKOUT2_DUTY_CYCLE   	32'h0011	// Type=FLOAT; Min=0.001, Max=0.999
`define MMCME3_ADV__CLKOUT2_DUTY_CYCLE_SZ	64

`define MMCME3_ADV__CLKOUT2_PHASE   	32'h0012	// Type=FLOAT; Min=-360.000, Max=360.000
`define MMCME3_ADV__CLKOUT2_PHASE_SZ	64

`define MMCME3_ADV__CLKOUT2_USE_FINE_PS   	32'h0013	// Type=BOOLSTRING; Values=FALSE,TRUE
`define MMCME3_ADV__CLKOUT2_USE_FINE_PS_SZ	40

`define MMCME3_ADV__CLKOUT3_DIVIDE   	32'h0014	// Type=DECIMAL; Min=1, Max=128
`define MMCME3_ADV__CLKOUT3_DIVIDE_SZ	32

`define MMCME3_ADV__CLKOUT3_DUTY_CYCLE   	32'h0015	// Type=FLOAT; Min=0.001, Max=0.999
`define MMCME3_ADV__CLKOUT3_DUTY_CYCLE_SZ	64

`define MMCME3_ADV__CLKOUT3_PHASE   	32'h0016	// Type=FLOAT; Min=-360.000, Max=360.000
`define MMCME3_ADV__CLKOUT3_PHASE_SZ	64

`define MMCME3_ADV__CLKOUT3_USE_FINE_PS   	32'h0017	// Type=BOOLSTRING; Values=FALSE,TRUE
`define MMCME3_ADV__CLKOUT3_USE_FINE_PS_SZ	40

`define MMCME3_ADV__CLKOUT4_CASCADE   	32'h0018	// Type=BOOLSTRING; Values=FALSE,TRUE
`define MMCME3_ADV__CLKOUT4_CASCADE_SZ	40

`define MMCME3_ADV__CLKOUT4_DIVIDE   	32'h0019	// Type=DECIMAL; Min=1, Max=128
`define MMCME3_ADV__CLKOUT4_DIVIDE_SZ	32

`define MMCME3_ADV__CLKOUT4_DUTY_CYCLE   	32'h001a	// Type=FLOAT; Min=0.001, Max=0.999
`define MMCME3_ADV__CLKOUT4_DUTY_CYCLE_SZ	64

`define MMCME3_ADV__CLKOUT4_PHASE   	32'h001b	// Type=FLOAT; Min=-360.000, Max=360.000
`define MMCME3_ADV__CLKOUT4_PHASE_SZ	64

`define MMCME3_ADV__CLKOUT4_USE_FINE_PS   	32'h001c	// Type=BOOLSTRING; Values=FALSE,TRUE
`define MMCME3_ADV__CLKOUT4_USE_FINE_PS_SZ	40

`define MMCME3_ADV__CLKOUT5_DIVIDE   	32'h001d	// Type=DECIMAL; Min=1, Max=128
`define MMCME3_ADV__CLKOUT5_DIVIDE_SZ	32

`define MMCME3_ADV__CLKOUT5_DUTY_CYCLE   	32'h001e	// Type=FLOAT; Min=0.001, Max=0.999
`define MMCME3_ADV__CLKOUT5_DUTY_CYCLE_SZ	64

`define MMCME3_ADV__CLKOUT5_PHASE   	32'h001f	// Type=FLOAT; Min=-360.000, Max=360.000
`define MMCME3_ADV__CLKOUT5_PHASE_SZ	64

`define MMCME3_ADV__CLKOUT5_USE_FINE_PS   	32'h0020	// Type=BOOLSTRING; Values=FALSE,TRUE
`define MMCME3_ADV__CLKOUT5_USE_FINE_PS_SZ	40

`define MMCME3_ADV__CLKOUT6_DIVIDE   	32'h0021	// Type=DECIMAL; Min=1, Max=128
`define MMCME3_ADV__CLKOUT6_DIVIDE_SZ	32

`define MMCME3_ADV__CLKOUT6_DUTY_CYCLE   	32'h0022	// Type=FLOAT; Min=0.001, Max=0.999
`define MMCME3_ADV__CLKOUT6_DUTY_CYCLE_SZ	64

`define MMCME3_ADV__CLKOUT6_PHASE   	32'h0023	// Type=FLOAT; Min=-360.000, Max=360.000
`define MMCME3_ADV__CLKOUT6_PHASE_SZ	64

`define MMCME3_ADV__CLKOUT6_USE_FINE_PS   	32'h0024	// Type=BOOLSTRING; Values=FALSE,TRUE
`define MMCME3_ADV__CLKOUT6_USE_FINE_PS_SZ	40

`define MMCME3_ADV__CLKPFD_FREQ_MAX   	32'h0025	// Type=FLOAT; Min=450.000, Max=550.000
`define MMCME3_ADV__CLKPFD_FREQ_MAX_SZ	64

`define MMCME3_ADV__CLKPFD_FREQ_MIN   	32'h0026	// Type=FLOAT; Min=10.000, Max=10.000
`define MMCME3_ADV__CLKPFD_FREQ_MIN_SZ	64

`define MMCME3_ADV__COMPENSATION   	32'h0027	// Type=STRING; Values=AUTO,BUF_IN,EXTERNAL,INTERNAL,ZHOLD
`define MMCME3_ADV__COMPENSATION_SZ	64

`define MMCME3_ADV__DIVCLK_DIVIDE   	32'h0028	// Type=DECIMAL; Min=1, Max=106
`define MMCME3_ADV__DIVCLK_DIVIDE_SZ	32

`define MMCME3_ADV__IS_CLKFBIN_INVERTED   	32'h0029	// Type=BINARY; Min=1'b0, Max=1'b1
`define MMCME3_ADV__IS_CLKFBIN_INVERTED_SZ	1

`define MMCME3_ADV__IS_CLKIN1_INVERTED   	32'h002a	// Type=BINARY; Min=1'b0, Max=1'b1
`define MMCME3_ADV__IS_CLKIN1_INVERTED_SZ	1

`define MMCME3_ADV__IS_CLKIN2_INVERTED   	32'h002b	// Type=BINARY; Min=1'b0, Max=1'b1
`define MMCME3_ADV__IS_CLKIN2_INVERTED_SZ	1

`define MMCME3_ADV__IS_CLKINSEL_INVERTED   	32'h002c	// Type=BINARY; Min=1'b0, Max=1'b1
`define MMCME3_ADV__IS_CLKINSEL_INVERTED_SZ	1

`define MMCME3_ADV__IS_PSEN_INVERTED   	32'h002d	// Type=BINARY; Min=1'b0, Max=1'b1
`define MMCME3_ADV__IS_PSEN_INVERTED_SZ	1

`define MMCME3_ADV__IS_PSINCDEC_INVERTED   	32'h002e	// Type=BINARY; Min=1'b0, Max=1'b1
`define MMCME3_ADV__IS_PSINCDEC_INVERTED_SZ	1

`define MMCME3_ADV__IS_PWRDWN_INVERTED   	32'h002f	// Type=BINARY; Min=1'b0, Max=1'b1
`define MMCME3_ADV__IS_PWRDWN_INVERTED_SZ	1

`define MMCME3_ADV__IS_RST_INVERTED   	32'h0030	// Type=BINARY; Min=1'b0, Max=1'b1
`define MMCME3_ADV__IS_RST_INVERTED_SZ	1

`define MMCME3_ADV__REF_JITTER1   	32'h0031	// Type=FLOAT; Min=0.000, Max=0.999
`define MMCME3_ADV__REF_JITTER1_SZ	64

`define MMCME3_ADV__REF_JITTER2   	32'h0032	// Type=FLOAT; Min=0.000, Max=0.999
`define MMCME3_ADV__REF_JITTER2_SZ	64

`define MMCME3_ADV__SS_EN   	32'h0033	// Type=BOOLSTRING; Values=FALSE,TRUE
`define MMCME3_ADV__SS_EN_SZ	40

`define MMCME3_ADV__SS_MODE   	32'h0034	// Type=STRING; Values=CENTER_HIGH,CENTER_LOW,DOWN_HIGH,DOWN_LOW
`define MMCME3_ADV__SS_MODE_SZ	88

`define MMCME3_ADV__SS_MOD_PERIOD   	32'h0035	// Type=DECIMAL; Min=4000, Max=40000
`define MMCME3_ADV__SS_MOD_PERIOD_SZ	32

`define MMCME3_ADV__STARTUP_WAIT   	32'h0036	// Type=BOOLSTRING; Values=FALSE,TRUE
`define MMCME3_ADV__STARTUP_WAIT_SZ	40

`define MMCME3_ADV__VCOCLK_FREQ_MAX   	32'h0037	// Type=FLOAT; Min=1200.000, Max=1600.000
`define MMCME3_ADV__VCOCLK_FREQ_MAX_SZ	64

`define MMCME3_ADV__VCOCLK_FREQ_MIN   	32'h0038	// Type=FLOAT; Min=600.000, Max=600.000
`define MMCME3_ADV__VCOCLK_FREQ_MIN_SZ	64

`endif  // B_MMCME3_ADV_DEFINES_VH
