///////////////////////////////////////////////////////////////////////////////
//  Copyright (c) 2011 Xilinx Inc.
//  All Right Reserved.
///////////////////////////////////////////////////////////////////////////////
//
//   ____   ___
//  /   /\/   / 
// /___/  \  /     Vendor      : Xilinx 
// \   \   \/      Version     : 2012.2
//  \   \          Description : Xilinx Unified Simulation Library Component
//  /   /                        
// /___/   /\      Filename    : PCIE_3_1.v
// \   \  /  \ 
//  \___\/\___\                    
//                                 
///////////////////////////////////////////////////////////////////////////////
//  Revision:
//
//  End Revision:
///////////////////////////////////////////////////////////////////////////////

`timescale 1 ps / 1 ps 

`celldefine
module PCIE_3_1 #(
  `ifdef XIL_TIMING //Simprim 
  parameter LOC = "UNPLACED",  
  `endif
  parameter ARI_CAP_ENABLE = "FALSE",
  parameter AXISTEN_IF_CC_ALIGNMENT_MODE = "FALSE",
  parameter AXISTEN_IF_CC_PARITY_CHK = "TRUE",
  parameter AXISTEN_IF_CQ_ALIGNMENT_MODE = "FALSE",
  parameter AXISTEN_IF_ENABLE_CLIENT_TAG = "FALSE",
  parameter [17:0] AXISTEN_IF_ENABLE_MSG_ROUTE = 18'h00000,
  parameter AXISTEN_IF_ENABLE_RX_MSG_INTFC = "FALSE",
  parameter AXISTEN_IF_RC_ALIGNMENT_MODE = "FALSE",
  parameter AXISTEN_IF_RC_STRADDLE = "FALSE",
  parameter AXISTEN_IF_RQ_ALIGNMENT_MODE = "FALSE",
  parameter AXISTEN_IF_RQ_PARITY_CHK = "TRUE",
  parameter [1:0] AXISTEN_IF_WIDTH = 2'h2,
  parameter CRM_CORE_CLK_FREQ_500 = "TRUE",
  parameter [1:0] CRM_USER_CLK_FREQ = 2'h2,
  parameter DEBUG_CFG_LOCAL_MGMT_REG_ACCESS_OVERRIDE = "FALSE",
  parameter DEBUG_PL_DISABLE_EI_INFER_IN_L0 = "FALSE",
  parameter DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS = "FALSE",
  parameter [7:0] DNSTREAM_LINK_NUM = 8'h00,
  parameter [8:0] LL_ACK_TIMEOUT = 9'h000,
  parameter LL_ACK_TIMEOUT_EN = "FALSE",
  parameter integer LL_ACK_TIMEOUT_FUNC = 0,
  parameter [15:0] LL_CPL_FC_UPDATE_TIMER = 16'h0000,
  parameter LL_CPL_FC_UPDATE_TIMER_OVERRIDE = "FALSE",
  parameter [15:0] LL_FC_UPDATE_TIMER = 16'h0000,
  parameter LL_FC_UPDATE_TIMER_OVERRIDE = "FALSE",
  parameter [15:0] LL_NP_FC_UPDATE_TIMER = 16'h0000,
  parameter LL_NP_FC_UPDATE_TIMER_OVERRIDE = "FALSE",
  parameter [15:0] LL_P_FC_UPDATE_TIMER = 16'h0000,
  parameter LL_P_FC_UPDATE_TIMER_OVERRIDE = "FALSE",
  parameter [8:0] LL_REPLAY_TIMEOUT = 9'h000,
  parameter LL_REPLAY_TIMEOUT_EN = "FALSE",
  parameter integer LL_REPLAY_TIMEOUT_FUNC = 0,
  parameter [9:0] LTR_TX_MESSAGE_MINIMUM_INTERVAL = 10'h0FA,
  parameter LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE = "FALSE",
  parameter LTR_TX_MESSAGE_ON_LTR_ENABLE = "FALSE",
  parameter [11:0] MCAP_CAP_NEXTPTR = 12'h000,
  parameter MCAP_CONFIGURE_OVERRIDE = "FALSE",
  parameter MCAP_ENABLE = "FALSE",
  parameter MCAP_EOS_DESIGN_SWITCH = "FALSE",
  parameter [31:0] MCAP_FPGA_BITSTREAM_VERSION = 32'h00000000,
  parameter MCAP_GATE_IO_ENABLE_DESIGN_SWITCH = "FALSE",
  parameter MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH = "FALSE",
  parameter MCAP_INPUT_GATE_DESIGN_SWITCH = "FALSE",
  parameter MCAP_INTERRUPT_ON_MCAP_EOS = "FALSE",
  parameter MCAP_INTERRUPT_ON_MCAP_ERROR = "FALSE",
  parameter [15:0] MCAP_VSEC_ID = 16'h0000,
  parameter [11:0] MCAP_VSEC_LEN = 12'h02C,
  parameter [3:0] MCAP_VSEC_REV = 4'h0,
  parameter PF0_AER_CAP_ECRC_CHECK_CAPABLE = "FALSE",
  parameter PF0_AER_CAP_ECRC_GEN_CAPABLE = "FALSE",
  parameter [11:0] PF0_AER_CAP_NEXTPTR = 12'h000,
  parameter [11:0] PF0_ARI_CAP_NEXTPTR = 12'h000,
  parameter [7:0] PF0_ARI_CAP_NEXT_FUNC = 8'h00,
  parameter [3:0] PF0_ARI_CAP_VER = 4'h1,
  parameter [5:0] PF0_BAR0_APERTURE_SIZE = 6'h03,
  parameter [2:0] PF0_BAR0_CONTROL = 3'h4,
  parameter [5:0] PF0_BAR1_APERTURE_SIZE = 6'h00,
  parameter [2:0] PF0_BAR1_CONTROL = 3'h0,
  parameter [4:0] PF0_BAR2_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF0_BAR2_CONTROL = 3'h4,
  parameter [4:0] PF0_BAR3_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF0_BAR3_CONTROL = 3'h0,
  parameter [4:0] PF0_BAR4_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF0_BAR4_CONTROL = 3'h4,
  parameter [4:0] PF0_BAR5_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF0_BAR5_CONTROL = 3'h0,
  parameter [7:0] PF0_BIST_REGISTER = 8'h00,
  parameter [7:0] PF0_CAPABILITY_POINTER = 8'h50,
  parameter [23:0] PF0_CLASS_CODE = 24'h000000,
  parameter [15:0] PF0_DEVICE_ID = 16'h0000,
  parameter PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT = "TRUE",
  parameter PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT = "TRUE",
  parameter PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT = "TRUE",
  parameter PF0_DEV_CAP2_ARI_FORWARD_ENABLE = "FALSE",
  parameter PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE = "TRUE",
  parameter PF0_DEV_CAP2_LTR_SUPPORT = "TRUE",
  parameter [1:0] PF0_DEV_CAP2_OBFF_SUPPORT = 2'h0,
  parameter PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT = "FALSE",
  parameter integer PF0_DEV_CAP_ENDPOINT_L0S_LATENCY = 0,
  parameter integer PF0_DEV_CAP_ENDPOINT_L1_LATENCY = 0,
  parameter PF0_DEV_CAP_EXT_TAG_SUPPORTED = "TRUE",
  parameter PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE = "TRUE",
  parameter [2:0] PF0_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3,
  parameter [11:0] PF0_DPA_CAP_NEXTPTR = 12'h000,
  parameter [4:0] PF0_DPA_CAP_SUB_STATE_CONTROL = 5'h00,
  parameter PF0_DPA_CAP_SUB_STATE_CONTROL_EN = "TRUE",
  parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 = 8'h00,
  parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 = 8'h00,
  parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 = 8'h00,
  parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 = 8'h00,
  parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 = 8'h00,
  parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 = 8'h00,
  parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 = 8'h00,
  parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 = 8'h00,
  parameter [3:0] PF0_DPA_CAP_VER = 4'h1,
  parameter [11:0] PF0_DSN_CAP_NEXTPTR = 12'h10C,
  parameter [4:0] PF0_EXPANSION_ROM_APERTURE_SIZE = 5'h03,
  parameter PF0_EXPANSION_ROM_ENABLE = "FALSE",
  parameter [7:0] PF0_INTERRUPT_LINE = 8'h00,
  parameter [2:0] PF0_INTERRUPT_PIN = 3'h1,
  parameter integer PF0_LINK_CAP_ASPM_SUPPORT = 0,
  parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 = 7,
  parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 = 7,
  parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3 = 7,
  parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1 = 7,
  parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2 = 7,
  parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3 = 7,
  parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 = 7,
  parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 = 7,
  parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3 = 7,
  parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1 = 7,
  parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2 = 7,
  parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3 = 7,
  parameter PF0_LINK_STATUS_SLOT_CLOCK_CONFIG = "TRUE",
  parameter [9:0] PF0_LTR_CAP_MAX_NOSNOOP_LAT = 10'h000,
  parameter [9:0] PF0_LTR_CAP_MAX_SNOOP_LAT = 10'h000,
  parameter [11:0] PF0_LTR_CAP_NEXTPTR = 12'h000,
  parameter [3:0] PF0_LTR_CAP_VER = 4'h1,
  parameter [7:0] PF0_MSIX_CAP_NEXTPTR = 8'h00,
  parameter integer PF0_MSIX_CAP_PBA_BIR = 0,
  parameter [28:0] PF0_MSIX_CAP_PBA_OFFSET = 29'h00000050,
  parameter integer PF0_MSIX_CAP_TABLE_BIR = 0,
  parameter [28:0] PF0_MSIX_CAP_TABLE_OFFSET = 29'h00000040,
  parameter [10:0] PF0_MSIX_CAP_TABLE_SIZE = 11'h000,
  parameter integer PF0_MSI_CAP_MULTIMSGCAP = 0,
  parameter [7:0] PF0_MSI_CAP_NEXTPTR = 8'h00,
  parameter PF0_MSI_CAP_PERVECMASKCAP = "FALSE",
  parameter [31:0] PF0_PB_CAP_DATA_REG_D0 = 32'h00000000,
  parameter [31:0] PF0_PB_CAP_DATA_REG_D0_SUSTAINED = 32'h00000000,
  parameter [31:0] PF0_PB_CAP_DATA_REG_D1 = 32'h00000000,
  parameter [31:0] PF0_PB_CAP_DATA_REG_D3HOT = 32'h00000000,
  parameter [11:0] PF0_PB_CAP_NEXTPTR = 12'h000,
  parameter PF0_PB_CAP_SYSTEM_ALLOCATED = "FALSE",
  parameter [3:0] PF0_PB_CAP_VER = 4'h1,
  parameter [7:0] PF0_PM_CAP_ID = 8'h01,
  parameter [7:0] PF0_PM_CAP_NEXTPTR = 8'h00,
  parameter PF0_PM_CAP_PMESUPPORT_D0 = "TRUE",
  parameter PF0_PM_CAP_PMESUPPORT_D1 = "TRUE",
  parameter PF0_PM_CAP_PMESUPPORT_D3HOT = "TRUE",
  parameter PF0_PM_CAP_SUPP_D1_STATE = "TRUE",
  parameter [2:0] PF0_PM_CAP_VER_ID = 3'h3,
  parameter PF0_PM_CSR_NOSOFTRESET = "TRUE",
  parameter PF0_RBAR_CAP_ENABLE = "FALSE",
  parameter [11:0] PF0_RBAR_CAP_NEXTPTR = 12'h000,
  parameter [19:0] PF0_RBAR_CAP_SIZE0 = 20'h00000,
  parameter [19:0] PF0_RBAR_CAP_SIZE1 = 20'h00000,
  parameter [19:0] PF0_RBAR_CAP_SIZE2 = 20'h00000,
  parameter [3:0] PF0_RBAR_CAP_VER = 4'h1,
  parameter [2:0] PF0_RBAR_CONTROL_INDEX0 = 3'h0,
  parameter [2:0] PF0_RBAR_CONTROL_INDEX1 = 3'h0,
  parameter [2:0] PF0_RBAR_CONTROL_INDEX2 = 3'h0,
  parameter [4:0] PF0_RBAR_CONTROL_SIZE0 = 5'h00,
  parameter [4:0] PF0_RBAR_CONTROL_SIZE1 = 5'h00,
  parameter [4:0] PF0_RBAR_CONTROL_SIZE2 = 5'h00,
  parameter [2:0] PF0_RBAR_NUM = 3'h1,
  parameter [7:0] PF0_REVISION_ID = 8'h00,
  parameter [11:0] PF0_SECONDARY_PCIE_CAP_NEXTPTR = 12'h000,
  parameter [4:0] PF0_SRIOV_BAR0_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF0_SRIOV_BAR0_CONTROL = 3'h4,
  parameter [4:0] PF0_SRIOV_BAR1_APERTURE_SIZE = 5'h00,
  parameter [2:0] PF0_SRIOV_BAR1_CONTROL = 3'h0,
  parameter [4:0] PF0_SRIOV_BAR2_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF0_SRIOV_BAR2_CONTROL = 3'h4,
  parameter [4:0] PF0_SRIOV_BAR3_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF0_SRIOV_BAR3_CONTROL = 3'h0,
  parameter [4:0] PF0_SRIOV_BAR4_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF0_SRIOV_BAR4_CONTROL = 3'h4,
  parameter [4:0] PF0_SRIOV_BAR5_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF0_SRIOV_BAR5_CONTROL = 3'h0,
  parameter [15:0] PF0_SRIOV_CAP_INITIAL_VF = 16'h0000,
  parameter [11:0] PF0_SRIOV_CAP_NEXTPTR = 12'h000,
  parameter [15:0] PF0_SRIOV_CAP_TOTAL_VF = 16'h0000,
  parameter [3:0] PF0_SRIOV_CAP_VER = 4'h1,
  parameter [15:0] PF0_SRIOV_FIRST_VF_OFFSET = 16'h0000,
  parameter [15:0] PF0_SRIOV_FUNC_DEP_LINK = 16'h0000,
  parameter [31:0] PF0_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000,
  parameter [15:0] PF0_SRIOV_VF_DEVICE_ID = 16'h0000,
  parameter [15:0] PF0_SUBSYSTEM_ID = 16'h0000,
  parameter PF0_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE",
  parameter PF0_TPHR_CAP_ENABLE = "FALSE",
  parameter PF0_TPHR_CAP_INT_VEC_MODE = "TRUE",
  parameter [11:0] PF0_TPHR_CAP_NEXTPTR = 12'h000,
  parameter [2:0] PF0_TPHR_CAP_ST_MODE_SEL = 3'h0,
  parameter [1:0] PF0_TPHR_CAP_ST_TABLE_LOC = 2'h0,
  parameter [10:0] PF0_TPHR_CAP_ST_TABLE_SIZE = 11'h000,
  parameter [3:0] PF0_TPHR_CAP_VER = 4'h1,
  parameter PF0_VC_CAP_ENABLE = "FALSE",
  parameter [11:0] PF0_VC_CAP_NEXTPTR = 12'h000,
  parameter [3:0] PF0_VC_CAP_VER = 4'h1,
  parameter PF1_AER_CAP_ECRC_CHECK_CAPABLE = "FALSE",
  parameter PF1_AER_CAP_ECRC_GEN_CAPABLE = "FALSE",
  parameter [11:0] PF1_AER_CAP_NEXTPTR = 12'h000,
  parameter [11:0] PF1_ARI_CAP_NEXTPTR = 12'h000,
  parameter [7:0] PF1_ARI_CAP_NEXT_FUNC = 8'h00,
  parameter [5:0] PF1_BAR0_APERTURE_SIZE = 6'h03,
  parameter [2:0] PF1_BAR0_CONTROL = 3'h4,
  parameter [5:0] PF1_BAR1_APERTURE_SIZE = 6'h00,
  parameter [2:0] PF1_BAR1_CONTROL = 3'h0,
  parameter [4:0] PF1_BAR2_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF1_BAR2_CONTROL = 3'h4,
  parameter [4:0] PF1_BAR3_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF1_BAR3_CONTROL = 3'h0,
  parameter [4:0] PF1_BAR4_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF1_BAR4_CONTROL = 3'h4,
  parameter [4:0] PF1_BAR5_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF1_BAR5_CONTROL = 3'h0,
  parameter [7:0] PF1_BIST_REGISTER = 8'h00,
  parameter [7:0] PF1_CAPABILITY_POINTER = 8'h50,
  parameter [23:0] PF1_CLASS_CODE = 24'h000000,
  parameter [15:0] PF1_DEVICE_ID = 16'h0000,
  parameter [2:0] PF1_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3,
  parameter [11:0] PF1_DPA_CAP_NEXTPTR = 12'h000,
  parameter [4:0] PF1_DPA_CAP_SUB_STATE_CONTROL = 5'h00,
  parameter PF1_DPA_CAP_SUB_STATE_CONTROL_EN = "TRUE",
  parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 = 8'h00,
  parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 = 8'h00,
  parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 = 8'h00,
  parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 = 8'h00,
  parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 = 8'h00,
  parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 = 8'h00,
  parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 = 8'h00,
  parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 = 8'h00,
  parameter [3:0] PF1_DPA_CAP_VER = 4'h1,
  parameter [11:0] PF1_DSN_CAP_NEXTPTR = 12'h10C,
  parameter [4:0] PF1_EXPANSION_ROM_APERTURE_SIZE = 5'h03,
  parameter PF1_EXPANSION_ROM_ENABLE = "FALSE",
  parameter [7:0] PF1_INTERRUPT_LINE = 8'h00,
  parameter [2:0] PF1_INTERRUPT_PIN = 3'h1,
  parameter [7:0] PF1_MSIX_CAP_NEXTPTR = 8'h00,
  parameter integer PF1_MSIX_CAP_PBA_BIR = 0,
  parameter [28:0] PF1_MSIX_CAP_PBA_OFFSET = 29'h00000050,
  parameter integer PF1_MSIX_CAP_TABLE_BIR = 0,
  parameter [28:0] PF1_MSIX_CAP_TABLE_OFFSET = 29'h00000040,
  parameter [10:0] PF1_MSIX_CAP_TABLE_SIZE = 11'h000,
  parameter integer PF1_MSI_CAP_MULTIMSGCAP = 0,
  parameter [7:0] PF1_MSI_CAP_NEXTPTR = 8'h00,
  parameter PF1_MSI_CAP_PERVECMASKCAP = "FALSE",
  parameter [31:0] PF1_PB_CAP_DATA_REG_D0 = 32'h00000000,
  parameter [31:0] PF1_PB_CAP_DATA_REG_D0_SUSTAINED = 32'h00000000,
  parameter [31:0] PF1_PB_CAP_DATA_REG_D1 = 32'h00000000,
  parameter [31:0] PF1_PB_CAP_DATA_REG_D3HOT = 32'h00000000,
  parameter [11:0] PF1_PB_CAP_NEXTPTR = 12'h000,
  parameter PF1_PB_CAP_SYSTEM_ALLOCATED = "FALSE",
  parameter [3:0] PF1_PB_CAP_VER = 4'h1,
  parameter [7:0] PF1_PM_CAP_ID = 8'h01,
  parameter [7:0] PF1_PM_CAP_NEXTPTR = 8'h00,
  parameter [2:0] PF1_PM_CAP_VER_ID = 3'h3,
  parameter PF1_RBAR_CAP_ENABLE = "FALSE",
  parameter [11:0] PF1_RBAR_CAP_NEXTPTR = 12'h000,
  parameter [19:0] PF1_RBAR_CAP_SIZE0 = 20'h00000,
  parameter [19:0] PF1_RBAR_CAP_SIZE1 = 20'h00000,
  parameter [19:0] PF1_RBAR_CAP_SIZE2 = 20'h00000,
  parameter [3:0] PF1_RBAR_CAP_VER = 4'h1,
  parameter [2:0] PF1_RBAR_CONTROL_INDEX0 = 3'h0,
  parameter [2:0] PF1_RBAR_CONTROL_INDEX1 = 3'h0,
  parameter [2:0] PF1_RBAR_CONTROL_INDEX2 = 3'h0,
  parameter [4:0] PF1_RBAR_CONTROL_SIZE0 = 5'h00,
  parameter [4:0] PF1_RBAR_CONTROL_SIZE1 = 5'h00,
  parameter [4:0] PF1_RBAR_CONTROL_SIZE2 = 5'h00,
  parameter [2:0] PF1_RBAR_NUM = 3'h1,
  parameter [7:0] PF1_REVISION_ID = 8'h00,
  parameter [4:0] PF1_SRIOV_BAR0_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF1_SRIOV_BAR0_CONTROL = 3'h4,
  parameter [4:0] PF1_SRIOV_BAR1_APERTURE_SIZE = 5'h00,
  parameter [2:0] PF1_SRIOV_BAR1_CONTROL = 3'h0,
  parameter [4:0] PF1_SRIOV_BAR2_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF1_SRIOV_BAR2_CONTROL = 3'h4,
  parameter [4:0] PF1_SRIOV_BAR3_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF1_SRIOV_BAR3_CONTROL = 3'h0,
  parameter [4:0] PF1_SRIOV_BAR4_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF1_SRIOV_BAR4_CONTROL = 3'h4,
  parameter [4:0] PF1_SRIOV_BAR5_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF1_SRIOV_BAR5_CONTROL = 3'h0,
  parameter [15:0] PF1_SRIOV_CAP_INITIAL_VF = 16'h0000,
  parameter [11:0] PF1_SRIOV_CAP_NEXTPTR = 12'h000,
  parameter [15:0] PF1_SRIOV_CAP_TOTAL_VF = 16'h0000,
  parameter [3:0] PF1_SRIOV_CAP_VER = 4'h1,
  parameter [15:0] PF1_SRIOV_FIRST_VF_OFFSET = 16'h0000,
  parameter [15:0] PF1_SRIOV_FUNC_DEP_LINK = 16'h0000,
  parameter [31:0] PF1_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000,
  parameter [15:0] PF1_SRIOV_VF_DEVICE_ID = 16'h0000,
  parameter [15:0] PF1_SUBSYSTEM_ID = 16'h0000,
  parameter PF1_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE",
  parameter PF1_TPHR_CAP_ENABLE = "FALSE",
  parameter PF1_TPHR_CAP_INT_VEC_MODE = "TRUE",
  parameter [11:0] PF1_TPHR_CAP_NEXTPTR = 12'h000,
  parameter [2:0] PF1_TPHR_CAP_ST_MODE_SEL = 3'h0,
  parameter [1:0] PF1_TPHR_CAP_ST_TABLE_LOC = 2'h0,
  parameter [10:0] PF1_TPHR_CAP_ST_TABLE_SIZE = 11'h000,
  parameter [3:0] PF1_TPHR_CAP_VER = 4'h1,
  parameter PF2_AER_CAP_ECRC_CHECK_CAPABLE = "FALSE",
  parameter PF2_AER_CAP_ECRC_GEN_CAPABLE = "FALSE",
  parameter [11:0] PF2_AER_CAP_NEXTPTR = 12'h000,
  parameter [11:0] PF2_ARI_CAP_NEXTPTR = 12'h000,
  parameter [7:0] PF2_ARI_CAP_NEXT_FUNC = 8'h00,
  parameter [5:0] PF2_BAR0_APERTURE_SIZE = 6'h03,
  parameter [2:0] PF2_BAR0_CONTROL = 3'h4,
  parameter [5:0] PF2_BAR1_APERTURE_SIZE = 6'h00,
  parameter [2:0] PF2_BAR1_CONTROL = 3'h0,
  parameter [4:0] PF2_BAR2_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF2_BAR2_CONTROL = 3'h4,
  parameter [4:0] PF2_BAR3_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF2_BAR3_CONTROL = 3'h0,
  parameter [4:0] PF2_BAR4_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF2_BAR4_CONTROL = 3'h4,
  parameter [4:0] PF2_BAR5_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF2_BAR5_CONTROL = 3'h0,
  parameter [7:0] PF2_BIST_REGISTER = 8'h00,
  parameter [7:0] PF2_CAPABILITY_POINTER = 8'h50,
  parameter [23:0] PF2_CLASS_CODE = 24'h000000,
  parameter [15:0] PF2_DEVICE_ID = 16'h0000,
  parameter [2:0] PF2_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3,
  parameter [11:0] PF2_DPA_CAP_NEXTPTR = 12'h000,
  parameter [4:0] PF2_DPA_CAP_SUB_STATE_CONTROL = 5'h00,
  parameter PF2_DPA_CAP_SUB_STATE_CONTROL_EN = "TRUE",
  parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 = 8'h00,
  parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 = 8'h00,
  parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 = 8'h00,
  parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 = 8'h00,
  parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 = 8'h00,
  parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 = 8'h00,
  parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 = 8'h00,
  parameter [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 = 8'h00,
  parameter [3:0] PF2_DPA_CAP_VER = 4'h1,
  parameter [11:0] PF2_DSN_CAP_NEXTPTR = 12'h10C,
  parameter [4:0] PF2_EXPANSION_ROM_APERTURE_SIZE = 5'h03,
  parameter PF2_EXPANSION_ROM_ENABLE = "FALSE",
  parameter [7:0] PF2_INTERRUPT_LINE = 8'h00,
  parameter [2:0] PF2_INTERRUPT_PIN = 3'h1,
  parameter [7:0] PF2_MSIX_CAP_NEXTPTR = 8'h00,
  parameter integer PF2_MSIX_CAP_PBA_BIR = 0,
  parameter [28:0] PF2_MSIX_CAP_PBA_OFFSET = 29'h00000050,
  parameter integer PF2_MSIX_CAP_TABLE_BIR = 0,
  parameter [28:0] PF2_MSIX_CAP_TABLE_OFFSET = 29'h00000040,
  parameter [10:0] PF2_MSIX_CAP_TABLE_SIZE = 11'h000,
  parameter integer PF2_MSI_CAP_MULTIMSGCAP = 0,
  parameter [7:0] PF2_MSI_CAP_NEXTPTR = 8'h00,
  parameter PF2_MSI_CAP_PERVECMASKCAP = "FALSE",
  parameter [31:0] PF2_PB_CAP_DATA_REG_D0 = 32'h00000000,
  parameter [31:0] PF2_PB_CAP_DATA_REG_D0_SUSTAINED = 32'h00000000,
  parameter [31:0] PF2_PB_CAP_DATA_REG_D1 = 32'h00000000,
  parameter [31:0] PF2_PB_CAP_DATA_REG_D3HOT = 32'h00000000,
  parameter [11:0] PF2_PB_CAP_NEXTPTR = 12'h000,
  parameter PF2_PB_CAP_SYSTEM_ALLOCATED = "FALSE",
  parameter [3:0] PF2_PB_CAP_VER = 4'h1,
  parameter [7:0] PF2_PM_CAP_ID = 8'h01,
  parameter [7:0] PF2_PM_CAP_NEXTPTR = 8'h00,
  parameter [2:0] PF2_PM_CAP_VER_ID = 3'h3,
  parameter PF2_RBAR_CAP_ENABLE = "FALSE",
  parameter [11:0] PF2_RBAR_CAP_NEXTPTR = 12'h000,
  parameter [19:0] PF2_RBAR_CAP_SIZE0 = 20'h00000,
  parameter [19:0] PF2_RBAR_CAP_SIZE1 = 20'h00000,
  parameter [19:0] PF2_RBAR_CAP_SIZE2 = 20'h00000,
  parameter [3:0] PF2_RBAR_CAP_VER = 4'h1,
  parameter [2:0] PF2_RBAR_CONTROL_INDEX0 = 3'h0,
  parameter [2:0] PF2_RBAR_CONTROL_INDEX1 = 3'h0,
  parameter [2:0] PF2_RBAR_CONTROL_INDEX2 = 3'h0,
  parameter [4:0] PF2_RBAR_CONTROL_SIZE0 = 5'h00,
  parameter [4:0] PF2_RBAR_CONTROL_SIZE1 = 5'h00,
  parameter [4:0] PF2_RBAR_CONTROL_SIZE2 = 5'h00,
  parameter [2:0] PF2_RBAR_NUM = 3'h1,
  parameter [7:0] PF2_REVISION_ID = 8'h00,
  parameter [4:0] PF2_SRIOV_BAR0_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF2_SRIOV_BAR0_CONTROL = 3'h4,
  parameter [4:0] PF2_SRIOV_BAR1_APERTURE_SIZE = 5'h00,
  parameter [2:0] PF2_SRIOV_BAR1_CONTROL = 3'h0,
  parameter [4:0] PF2_SRIOV_BAR2_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF2_SRIOV_BAR2_CONTROL = 3'h4,
  parameter [4:0] PF2_SRIOV_BAR3_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF2_SRIOV_BAR3_CONTROL = 3'h0,
  parameter [4:0] PF2_SRIOV_BAR4_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF2_SRIOV_BAR4_CONTROL = 3'h4,
  parameter [4:0] PF2_SRIOV_BAR5_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF2_SRIOV_BAR5_CONTROL = 3'h0,
  parameter [15:0] PF2_SRIOV_CAP_INITIAL_VF = 16'h0000,
  parameter [11:0] PF2_SRIOV_CAP_NEXTPTR = 12'h000,
  parameter [15:0] PF2_SRIOV_CAP_TOTAL_VF = 16'h0000,
  parameter [3:0] PF2_SRIOV_CAP_VER = 4'h1,
  parameter [15:0] PF2_SRIOV_FIRST_VF_OFFSET = 16'h0000,
  parameter [15:0] PF2_SRIOV_FUNC_DEP_LINK = 16'h0000,
  parameter [31:0] PF2_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000,
  parameter [15:0] PF2_SRIOV_VF_DEVICE_ID = 16'h0000,
  parameter [15:0] PF2_SUBSYSTEM_ID = 16'h0000,
  parameter PF2_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE",
  parameter PF2_TPHR_CAP_ENABLE = "FALSE",
  parameter PF2_TPHR_CAP_INT_VEC_MODE = "TRUE",
  parameter [11:0] PF2_TPHR_CAP_NEXTPTR = 12'h000,
  parameter [2:0] PF2_TPHR_CAP_ST_MODE_SEL = 3'h0,
  parameter [1:0] PF2_TPHR_CAP_ST_TABLE_LOC = 2'h0,
  parameter [10:0] PF2_TPHR_CAP_ST_TABLE_SIZE = 11'h000,
  parameter [3:0] PF2_TPHR_CAP_VER = 4'h1,
  parameter PF3_AER_CAP_ECRC_CHECK_CAPABLE = "FALSE",
  parameter PF3_AER_CAP_ECRC_GEN_CAPABLE = "FALSE",
  parameter [11:0] PF3_AER_CAP_NEXTPTR = 12'h000,
  parameter [11:0] PF3_ARI_CAP_NEXTPTR = 12'h000,
  parameter [7:0] PF3_ARI_CAP_NEXT_FUNC = 8'h00,
  parameter [5:0] PF3_BAR0_APERTURE_SIZE = 6'h03,
  parameter [2:0] PF3_BAR0_CONTROL = 3'h4,
  parameter [5:0] PF3_BAR1_APERTURE_SIZE = 6'h00,
  parameter [2:0] PF3_BAR1_CONTROL = 3'h0,
  parameter [4:0] PF3_BAR2_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF3_BAR2_CONTROL = 3'h4,
  parameter [4:0] PF3_BAR3_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF3_BAR3_CONTROL = 3'h0,
  parameter [4:0] PF3_BAR4_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF3_BAR4_CONTROL = 3'h4,
  parameter [4:0] PF3_BAR5_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF3_BAR5_CONTROL = 3'h0,
  parameter [7:0] PF3_BIST_REGISTER = 8'h00,
  parameter [7:0] PF3_CAPABILITY_POINTER = 8'h50,
  parameter [23:0] PF3_CLASS_CODE = 24'h000000,
  parameter [15:0] PF3_DEVICE_ID = 16'h0000,
  parameter [2:0] PF3_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3,
  parameter [11:0] PF3_DPA_CAP_NEXTPTR = 12'h000,
  parameter [4:0] PF3_DPA_CAP_SUB_STATE_CONTROL = 5'h00,
  parameter PF3_DPA_CAP_SUB_STATE_CONTROL_EN = "TRUE",
  parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 = 8'h00,
  parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 = 8'h00,
  parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 = 8'h00,
  parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 = 8'h00,
  parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 = 8'h00,
  parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 = 8'h00,
  parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 = 8'h00,
  parameter [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 = 8'h00,
  parameter [3:0] PF3_DPA_CAP_VER = 4'h1,
  parameter [11:0] PF3_DSN_CAP_NEXTPTR = 12'h10C,
  parameter [4:0] PF3_EXPANSION_ROM_APERTURE_SIZE = 5'h03,
  parameter PF3_EXPANSION_ROM_ENABLE = "FALSE",
  parameter [7:0] PF3_INTERRUPT_LINE = 8'h00,
  parameter [2:0] PF3_INTERRUPT_PIN = 3'h1,
  parameter [7:0] PF3_MSIX_CAP_NEXTPTR = 8'h00,
  parameter integer PF3_MSIX_CAP_PBA_BIR = 0,
  parameter [28:0] PF3_MSIX_CAP_PBA_OFFSET = 29'h00000050,
  parameter integer PF3_MSIX_CAP_TABLE_BIR = 0,
  parameter [28:0] PF3_MSIX_CAP_TABLE_OFFSET = 29'h00000040,
  parameter [10:0] PF3_MSIX_CAP_TABLE_SIZE = 11'h000,
  parameter integer PF3_MSI_CAP_MULTIMSGCAP = 0,
  parameter [7:0] PF3_MSI_CAP_NEXTPTR = 8'h00,
  parameter PF3_MSI_CAP_PERVECMASKCAP = "FALSE",
  parameter [31:0] PF3_PB_CAP_DATA_REG_D0 = 32'h00000000,
  parameter [31:0] PF3_PB_CAP_DATA_REG_D0_SUSTAINED = 32'h00000000,
  parameter [31:0] PF3_PB_CAP_DATA_REG_D1 = 32'h00000000,
  parameter [31:0] PF3_PB_CAP_DATA_REG_D3HOT = 32'h00000000,
  parameter [11:0] PF3_PB_CAP_NEXTPTR = 12'h000,
  parameter PF3_PB_CAP_SYSTEM_ALLOCATED = "FALSE",
  parameter [3:0] PF3_PB_CAP_VER = 4'h1,
  parameter [7:0] PF3_PM_CAP_ID = 8'h01,
  parameter [7:0] PF3_PM_CAP_NEXTPTR = 8'h00,
  parameter [2:0] PF3_PM_CAP_VER_ID = 3'h3,
  parameter PF3_RBAR_CAP_ENABLE = "FALSE",
  parameter [11:0] PF3_RBAR_CAP_NEXTPTR = 12'h000,
  parameter [19:0] PF3_RBAR_CAP_SIZE0 = 20'h00000,
  parameter [19:0] PF3_RBAR_CAP_SIZE1 = 20'h00000,
  parameter [19:0] PF3_RBAR_CAP_SIZE2 = 20'h00000,
  parameter [3:0] PF3_RBAR_CAP_VER = 4'h1,
  parameter [2:0] PF3_RBAR_CONTROL_INDEX0 = 3'h0,
  parameter [2:0] PF3_RBAR_CONTROL_INDEX1 = 3'h0,
  parameter [2:0] PF3_RBAR_CONTROL_INDEX2 = 3'h0,
  parameter [4:0] PF3_RBAR_CONTROL_SIZE0 = 5'h00,
  parameter [4:0] PF3_RBAR_CONTROL_SIZE1 = 5'h00,
  parameter [4:0] PF3_RBAR_CONTROL_SIZE2 = 5'h00,
  parameter [2:0] PF3_RBAR_NUM = 3'h1,
  parameter [7:0] PF3_REVISION_ID = 8'h00,
  parameter [4:0] PF3_SRIOV_BAR0_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF3_SRIOV_BAR0_CONTROL = 3'h4,
  parameter [4:0] PF3_SRIOV_BAR1_APERTURE_SIZE = 5'h00,
  parameter [2:0] PF3_SRIOV_BAR1_CONTROL = 3'h0,
  parameter [4:0] PF3_SRIOV_BAR2_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF3_SRIOV_BAR2_CONTROL = 3'h4,
  parameter [4:0] PF3_SRIOV_BAR3_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF3_SRIOV_BAR3_CONTROL = 3'h0,
  parameter [4:0] PF3_SRIOV_BAR4_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF3_SRIOV_BAR4_CONTROL = 3'h4,
  parameter [4:0] PF3_SRIOV_BAR5_APERTURE_SIZE = 5'h03,
  parameter [2:0] PF3_SRIOV_BAR5_CONTROL = 3'h0,
  parameter [15:0] PF3_SRIOV_CAP_INITIAL_VF = 16'h0000,
  parameter [11:0] PF3_SRIOV_CAP_NEXTPTR = 12'h000,
  parameter [15:0] PF3_SRIOV_CAP_TOTAL_VF = 16'h0000,
  parameter [3:0] PF3_SRIOV_CAP_VER = 4'h1,
  parameter [15:0] PF3_SRIOV_FIRST_VF_OFFSET = 16'h0000,
  parameter [15:0] PF3_SRIOV_FUNC_DEP_LINK = 16'h0000,
  parameter [31:0] PF3_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000,
  parameter [15:0] PF3_SRIOV_VF_DEVICE_ID = 16'h0000,
  parameter [15:0] PF3_SUBSYSTEM_ID = 16'h0000,
  parameter PF3_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE",
  parameter PF3_TPHR_CAP_ENABLE = "FALSE",
  parameter PF3_TPHR_CAP_INT_VEC_MODE = "TRUE",
  parameter [11:0] PF3_TPHR_CAP_NEXTPTR = 12'h000,
  parameter [2:0] PF3_TPHR_CAP_ST_MODE_SEL = 3'h0,
  parameter [1:0] PF3_TPHR_CAP_ST_TABLE_LOC = 2'h0,
  parameter [10:0] PF3_TPHR_CAP_ST_TABLE_SIZE = 11'h000,
  parameter [3:0] PF3_TPHR_CAP_VER = 4'h1,
  parameter PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3 = "FALSE",
  parameter PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2 = "FALSE",
  parameter PL_DISABLE_EI_INFER_IN_L0 = "FALSE",
  parameter PL_DISABLE_GEN3_DC_BALANCE = "FALSE",
  parameter PL_DISABLE_GEN3_LFSR_UPDATE_ON_SKP = "TRUE",
  parameter PL_DISABLE_RETRAIN_ON_FRAMING_ERROR = "FALSE",
  parameter PL_DISABLE_SCRAMBLING = "FALSE",
  parameter PL_DISABLE_SYNC_HEADER_FRAMING_ERROR = "FALSE",
  parameter PL_DISABLE_UPCONFIG_CAPABLE = "FALSE",
  parameter PL_EQ_ADAPT_DISABLE_COEFF_CHECK = "FALSE",
  parameter PL_EQ_ADAPT_DISABLE_PRESET_CHECK = "FALSE",
  parameter [4:0] PL_EQ_ADAPT_ITER_COUNT = 5'h02,
  parameter [1:0] PL_EQ_ADAPT_REJECT_RETRY_COUNT = 2'h1,
  parameter PL_EQ_BYPASS_PHASE23 = "FALSE",
  parameter [2:0] PL_EQ_DEFAULT_GEN3_RX_PRESET_HINT = 3'h3,
  parameter [3:0] PL_EQ_DEFAULT_GEN3_TX_PRESET = 4'h4,
  parameter PL_EQ_PHASE01_RX_ADAPT = "FALSE",
  parameter PL_EQ_SHORT_ADAPT_PHASE = "FALSE",
  parameter [15:0] PL_LANE0_EQ_CONTROL = 16'h3F00,
  parameter [15:0] PL_LANE1_EQ_CONTROL = 16'h3F00,
  parameter [15:0] PL_LANE2_EQ_CONTROL = 16'h3F00,
  parameter [15:0] PL_LANE3_EQ_CONTROL = 16'h3F00,
  parameter [15:0] PL_LANE4_EQ_CONTROL = 16'h3F00,
  parameter [15:0] PL_LANE5_EQ_CONTROL = 16'h3F00,
  parameter [15:0] PL_LANE6_EQ_CONTROL = 16'h3F00,
  parameter [15:0] PL_LANE7_EQ_CONTROL = 16'h3F00,
  parameter [2:0] PL_LINK_CAP_MAX_LINK_SPEED = 3'h4,
  parameter [3:0] PL_LINK_CAP_MAX_LINK_WIDTH = 4'h8,
  parameter integer PL_N_FTS_COMCLK_GEN1 = 255,
  parameter integer PL_N_FTS_COMCLK_GEN2 = 255,
  parameter integer PL_N_FTS_COMCLK_GEN3 = 255,
  parameter integer PL_N_FTS_GEN1 = 255,
  parameter integer PL_N_FTS_GEN2 = 255,
  parameter integer PL_N_FTS_GEN3 = 255,
  parameter PL_REPORT_ALL_PHY_ERRORS = "TRUE",
  parameter PL_SIM_FAST_LINK_TRAINING = "FALSE",
  parameter PL_UPSTREAM_FACING = "TRUE",
  parameter [15:0] PM_ASPML0S_TIMEOUT = 16'h05DC,
  parameter [19:0] PM_ASPML1_ENTRY_DELAY = 20'h00000,
  parameter PM_ENABLE_L23_ENTRY = "FALSE",
  parameter PM_ENABLE_SLOT_POWER_CAPTURE = "TRUE",
  parameter [31:0] PM_L1_REENTRY_DELAY = 32'h00000000,
  parameter [19:0] PM_PME_SERVICE_TIMEOUT_DELAY = 20'h186A0,
  parameter [15:0] PM_PME_TURNOFF_ACK_DELAY = 16'h0064,
  parameter [31:0] SIM_JTAG_IDCODE = 32'h00000000,
  parameter SIM_VERSION = "1.0",
  parameter integer SPARE_BIT0 = 0,
  parameter integer SPARE_BIT1 = 0,
  parameter integer SPARE_BIT2 = 0,
  parameter integer SPARE_BIT3 = 0,
  parameter integer SPARE_BIT4 = 0,
  parameter integer SPARE_BIT5 = 0,
  parameter integer SPARE_BIT6 = 0,
  parameter integer SPARE_BIT7 = 0,
  parameter integer SPARE_BIT8 = 0,
  parameter [7:0] SPARE_BYTE0 = 8'h00,
  parameter [7:0] SPARE_BYTE1 = 8'h00,
  parameter [7:0] SPARE_BYTE2 = 8'h00,
  parameter [7:0] SPARE_BYTE3 = 8'h00,
  parameter [31:0] SPARE_WORD0 = 32'h00000000,
  parameter [31:0] SPARE_WORD1 = 32'h00000000,
  parameter [31:0] SPARE_WORD2 = 32'h00000000,
  parameter [31:0] SPARE_WORD3 = 32'h00000000,
  parameter SRIOV_CAP_ENABLE = "FALSE",
  parameter TL_COMPLETION_RAM_SIZE_16K = "TRUE",
  parameter [23:0] TL_COMPL_TIMEOUT_REG0 = 24'hBEBC20,
  parameter [27:0] TL_COMPL_TIMEOUT_REG1 = 28'h2FAF080,
  parameter [11:0] TL_CREDITS_CD = 12'h3E0,
  parameter [7:0] TL_CREDITS_CH = 8'h20,
  parameter [11:0] TL_CREDITS_NPD = 12'h028,
  parameter [7:0] TL_CREDITS_NPH = 8'h20,
  parameter [11:0] TL_CREDITS_PD = 12'h198,
  parameter [7:0] TL_CREDITS_PH = 8'h20,
  parameter TL_ENABLE_MESSAGE_RID_CHECK_ENABLE = "TRUE",
  parameter TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE = "FALSE",
  parameter TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE = "FALSE",
  parameter TL_LEGACY_MODE_ENABLE = "FALSE",
  parameter [1:0] TL_PF_ENABLE_REG = 2'h0,
  parameter TL_TX_MUX_STRICT_PRIORITY = "TRUE",
  parameter TWO_LAYER_MODE_DLCMSM_ENABLE = "TRUE",
  parameter TWO_LAYER_MODE_ENABLE = "FALSE",
  parameter TWO_LAYER_MODE_WIDTH_256 = "TRUE",
  parameter [11:0] VF0_ARI_CAP_NEXTPTR = 12'h000,
  parameter [7:0] VF0_CAPABILITY_POINTER = 8'h50,
  parameter integer VF0_MSIX_CAP_PBA_BIR = 0,
  parameter [28:0] VF0_MSIX_CAP_PBA_OFFSET = 29'h00000050,
  parameter integer VF0_MSIX_CAP_TABLE_BIR = 0,
  parameter [28:0] VF0_MSIX_CAP_TABLE_OFFSET = 29'h00000040,
  parameter [10:0] VF0_MSIX_CAP_TABLE_SIZE = 11'h000,
  parameter integer VF0_MSI_CAP_MULTIMSGCAP = 0,
  parameter [7:0] VF0_PM_CAP_ID = 8'h01,
  parameter [7:0] VF0_PM_CAP_NEXTPTR = 8'h00,
  parameter [2:0] VF0_PM_CAP_VER_ID = 3'h3,
  parameter VF0_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE",
  parameter VF0_TPHR_CAP_ENABLE = "FALSE",
  parameter VF0_TPHR_CAP_INT_VEC_MODE = "TRUE",
  parameter [11:0] VF0_TPHR_CAP_NEXTPTR = 12'h000,
  parameter [2:0] VF0_TPHR_CAP_ST_MODE_SEL = 3'h0,
  parameter [1:0] VF0_TPHR_CAP_ST_TABLE_LOC = 2'h0,
  parameter [10:0] VF0_TPHR_CAP_ST_TABLE_SIZE = 11'h000,
  parameter [3:0] VF0_TPHR_CAP_VER = 4'h1,
  parameter [11:0] VF1_ARI_CAP_NEXTPTR = 12'h000,
  parameter integer VF1_MSIX_CAP_PBA_BIR = 0,
  parameter [28:0] VF1_MSIX_CAP_PBA_OFFSET = 29'h00000050,
  parameter integer VF1_MSIX_CAP_TABLE_BIR = 0,
  parameter [28:0] VF1_MSIX_CAP_TABLE_OFFSET = 29'h00000040,
  parameter [10:0] VF1_MSIX_CAP_TABLE_SIZE = 11'h000,
  parameter integer VF1_MSI_CAP_MULTIMSGCAP = 0,
  parameter [7:0] VF1_PM_CAP_ID = 8'h01,
  parameter [7:0] VF1_PM_CAP_NEXTPTR = 8'h00,
  parameter [2:0] VF1_PM_CAP_VER_ID = 3'h3,
  parameter VF1_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE",
  parameter VF1_TPHR_CAP_ENABLE = "FALSE",
  parameter VF1_TPHR_CAP_INT_VEC_MODE = "TRUE",
  parameter [11:0] VF1_TPHR_CAP_NEXTPTR = 12'h000,
  parameter [2:0] VF1_TPHR_CAP_ST_MODE_SEL = 3'h0,
  parameter [1:0] VF1_TPHR_CAP_ST_TABLE_LOC = 2'h0,
  parameter [10:0] VF1_TPHR_CAP_ST_TABLE_SIZE = 11'h000,
  parameter [3:0] VF1_TPHR_CAP_VER = 4'h1,
  parameter [11:0] VF2_ARI_CAP_NEXTPTR = 12'h000,
  parameter integer VF2_MSIX_CAP_PBA_BIR = 0,
  parameter [28:0] VF2_MSIX_CAP_PBA_OFFSET = 29'h00000050,
  parameter integer VF2_MSIX_CAP_TABLE_BIR = 0,
  parameter [28:0] VF2_MSIX_CAP_TABLE_OFFSET = 29'h00000040,
  parameter [10:0] VF2_MSIX_CAP_TABLE_SIZE = 11'h000,
  parameter integer VF2_MSI_CAP_MULTIMSGCAP = 0,
  parameter [7:0] VF2_PM_CAP_ID = 8'h01,
  parameter [7:0] VF2_PM_CAP_NEXTPTR = 8'h00,
  parameter [2:0] VF2_PM_CAP_VER_ID = 3'h3,
  parameter VF2_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE",
  parameter VF2_TPHR_CAP_ENABLE = "FALSE",
  parameter VF2_TPHR_CAP_INT_VEC_MODE = "TRUE",
  parameter [11:0] VF2_TPHR_CAP_NEXTPTR = 12'h000,
  parameter [2:0] VF2_TPHR_CAP_ST_MODE_SEL = 3'h0,
  parameter [1:0] VF2_TPHR_CAP_ST_TABLE_LOC = 2'h0,
  parameter [10:0] VF2_TPHR_CAP_ST_TABLE_SIZE = 11'h000,
  parameter [3:0] VF2_TPHR_CAP_VER = 4'h1,
  parameter [11:0] VF3_ARI_CAP_NEXTPTR = 12'h000,
  parameter integer VF3_MSIX_CAP_PBA_BIR = 0,
  parameter [28:0] VF3_MSIX_CAP_PBA_OFFSET = 29'h00000050,
  parameter integer VF3_MSIX_CAP_TABLE_BIR = 0,
  parameter [28:0] VF3_MSIX_CAP_TABLE_OFFSET = 29'h00000040,
  parameter [10:0] VF3_MSIX_CAP_TABLE_SIZE = 11'h000,
  parameter integer VF3_MSI_CAP_MULTIMSGCAP = 0,
  parameter [7:0] VF3_PM_CAP_ID = 8'h01,
  parameter [7:0] VF3_PM_CAP_NEXTPTR = 8'h00,
  parameter [2:0] VF3_PM_CAP_VER_ID = 3'h3,
  parameter VF3_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE",
  parameter VF3_TPHR_CAP_ENABLE = "FALSE",
  parameter VF3_TPHR_CAP_INT_VEC_MODE = "TRUE",
  parameter [11:0] VF3_TPHR_CAP_NEXTPTR = 12'h000,
  parameter [2:0] VF3_TPHR_CAP_ST_MODE_SEL = 3'h0,
  parameter [1:0] VF3_TPHR_CAP_ST_TABLE_LOC = 2'h0,
  parameter [10:0] VF3_TPHR_CAP_ST_TABLE_SIZE = 11'h000,
  parameter [3:0] VF3_TPHR_CAP_VER = 4'h1,
  parameter [11:0] VF4_ARI_CAP_NEXTPTR = 12'h000,
  parameter integer VF4_MSIX_CAP_PBA_BIR = 0,
  parameter [28:0] VF4_MSIX_CAP_PBA_OFFSET = 29'h00000050,
  parameter integer VF4_MSIX_CAP_TABLE_BIR = 0,
  parameter [28:0] VF4_MSIX_CAP_TABLE_OFFSET = 29'h00000040,
  parameter [10:0] VF4_MSIX_CAP_TABLE_SIZE = 11'h000,
  parameter integer VF4_MSI_CAP_MULTIMSGCAP = 0,
  parameter [7:0] VF4_PM_CAP_ID = 8'h01,
  parameter [7:0] VF4_PM_CAP_NEXTPTR = 8'h00,
  parameter [2:0] VF4_PM_CAP_VER_ID = 3'h3,
  parameter VF4_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE",
  parameter VF4_TPHR_CAP_ENABLE = "FALSE",
  parameter VF4_TPHR_CAP_INT_VEC_MODE = "TRUE",
  parameter [11:0] VF4_TPHR_CAP_NEXTPTR = 12'h000,
  parameter [2:0] VF4_TPHR_CAP_ST_MODE_SEL = 3'h0,
  parameter [1:0] VF4_TPHR_CAP_ST_TABLE_LOC = 2'h0,
  parameter [10:0] VF4_TPHR_CAP_ST_TABLE_SIZE = 11'h000,
  parameter [3:0] VF4_TPHR_CAP_VER = 4'h1,
  parameter [11:0] VF5_ARI_CAP_NEXTPTR = 12'h000,
  parameter integer VF5_MSIX_CAP_PBA_BIR = 0,
  parameter [28:0] VF5_MSIX_CAP_PBA_OFFSET = 29'h00000050,
  parameter integer VF5_MSIX_CAP_TABLE_BIR = 0,
  parameter [28:0] VF5_MSIX_CAP_TABLE_OFFSET = 29'h00000040,
  parameter [10:0] VF5_MSIX_CAP_TABLE_SIZE = 11'h000,
  parameter integer VF5_MSI_CAP_MULTIMSGCAP = 0,
  parameter [7:0] VF5_PM_CAP_ID = 8'h01,
  parameter [7:0] VF5_PM_CAP_NEXTPTR = 8'h00,
  parameter [2:0] VF5_PM_CAP_VER_ID = 3'h3,
  parameter VF5_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE",
  parameter VF5_TPHR_CAP_ENABLE = "FALSE",
  parameter VF5_TPHR_CAP_INT_VEC_MODE = "TRUE",
  parameter [11:0] VF5_TPHR_CAP_NEXTPTR = 12'h000,
  parameter [2:0] VF5_TPHR_CAP_ST_MODE_SEL = 3'h0,
  parameter [1:0] VF5_TPHR_CAP_ST_TABLE_LOC = 2'h0,
  parameter [10:0] VF5_TPHR_CAP_ST_TABLE_SIZE = 11'h000,
  parameter [3:0] VF5_TPHR_CAP_VER = 4'h1,
  parameter [11:0] VF6_ARI_CAP_NEXTPTR = 12'h000,
  parameter integer VF6_MSIX_CAP_PBA_BIR = 0,
  parameter [28:0] VF6_MSIX_CAP_PBA_OFFSET = 29'h00000050,
  parameter integer VF6_MSIX_CAP_TABLE_BIR = 0,
  parameter [28:0] VF6_MSIX_CAP_TABLE_OFFSET = 29'h00000040,
  parameter [10:0] VF6_MSIX_CAP_TABLE_SIZE = 11'h000,
  parameter integer VF6_MSI_CAP_MULTIMSGCAP = 0,
  parameter [7:0] VF6_PM_CAP_ID = 8'h01,
  parameter [7:0] VF6_PM_CAP_NEXTPTR = 8'h00,
  parameter [2:0] VF6_PM_CAP_VER_ID = 3'h3,
  parameter VF6_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE",
  parameter VF6_TPHR_CAP_ENABLE = "FALSE",
  parameter VF6_TPHR_CAP_INT_VEC_MODE = "TRUE",
  parameter [11:0] VF6_TPHR_CAP_NEXTPTR = 12'h000,
  parameter [2:0] VF6_TPHR_CAP_ST_MODE_SEL = 3'h0,
  parameter [1:0] VF6_TPHR_CAP_ST_TABLE_LOC = 2'h0,
  parameter [10:0] VF6_TPHR_CAP_ST_TABLE_SIZE = 11'h000,
  parameter [3:0] VF6_TPHR_CAP_VER = 4'h1,
  parameter [11:0] VF7_ARI_CAP_NEXTPTR = 12'h000,
  parameter integer VF7_MSIX_CAP_PBA_BIR = 0,
  parameter [28:0] VF7_MSIX_CAP_PBA_OFFSET = 29'h00000050,
  parameter integer VF7_MSIX_CAP_TABLE_BIR = 0,
  parameter [28:0] VF7_MSIX_CAP_TABLE_OFFSET = 29'h00000040,
  parameter [10:0] VF7_MSIX_CAP_TABLE_SIZE = 11'h000,
  parameter integer VF7_MSI_CAP_MULTIMSGCAP = 0,
  parameter [7:0] VF7_PM_CAP_ID = 8'h01,
  parameter [7:0] VF7_PM_CAP_NEXTPTR = 8'h00,
  parameter [2:0] VF7_PM_CAP_VER_ID = 3'h3,
  parameter VF7_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE",
  parameter VF7_TPHR_CAP_ENABLE = "FALSE",
  parameter VF7_TPHR_CAP_INT_VEC_MODE = "TRUE",
  parameter [11:0] VF7_TPHR_CAP_NEXTPTR = 12'h000,
  parameter [2:0] VF7_TPHR_CAP_ST_MODE_SEL = 3'h0,
  parameter [1:0] VF7_TPHR_CAP_ST_TABLE_LOC = 2'h0,
  parameter [10:0] VF7_TPHR_CAP_ST_TABLE_SIZE = 11'h000,
  parameter [3:0] VF7_TPHR_CAP_VER = 4'h1
)(
  output [2:0] CFGCURRENTSPEED,
  output [3:0] CFGDPASUBSTATECHANGE,
  output CFGERRCOROUT,
  output CFGERRFATALOUT,
  output CFGERRNONFATALOUT,
  output [7:0] CFGEXTFUNCTIONNUMBER,
  output CFGEXTREADRECEIVED,
  output [9:0] CFGEXTREGISTERNUMBER,
  output [3:0] CFGEXTWRITEBYTEENABLE,
  output [31:0] CFGEXTWRITEDATA,
  output CFGEXTWRITERECEIVED,
  output [11:0] CFGFCCPLD,
  output [7:0] CFGFCCPLH,
  output [11:0] CFGFCNPD,
  output [7:0] CFGFCNPH,
  output [11:0] CFGFCPD,
  output [7:0] CFGFCPH,
  output [3:0] CFGFLRINPROCESS,
  output [11:0] CFGFUNCTIONPOWERSTATE,
  output [15:0] CFGFUNCTIONSTATUS,
  output CFGHOTRESETOUT,
  output [31:0] CFGINTERRUPTMSIDATA,
  output [3:0] CFGINTERRUPTMSIENABLE,
  output CFGINTERRUPTMSIFAIL,
  output CFGINTERRUPTMSIMASKUPDATE,
  output [11:0] CFGINTERRUPTMSIMMENABLE,
  output CFGINTERRUPTMSISENT,
  output [7:0] CFGINTERRUPTMSIVFENABLE,
  output [3:0] CFGINTERRUPTMSIXENABLE,
  output CFGINTERRUPTMSIXFAIL,
  output [3:0] CFGINTERRUPTMSIXMASK,
  output CFGINTERRUPTMSIXSENT,
  output [7:0] CFGINTERRUPTMSIXVFENABLE,
  output [7:0] CFGINTERRUPTMSIXVFMASK,
  output CFGINTERRUPTSENT,
  output [1:0] CFGLINKPOWERSTATE,
  output CFGLOCALERROR,
  output CFGLTRENABLE,
  output [5:0] CFGLTSSMSTATE,
  output [2:0] CFGMAXPAYLOAD,
  output [2:0] CFGMAXREADREQ,
  output [31:0] CFGMGMTREADDATA,
  output CFGMGMTREADWRITEDONE,
  output CFGMSGRECEIVED,
  output [7:0] CFGMSGRECEIVEDDATA,
  output [4:0] CFGMSGRECEIVEDTYPE,
  output CFGMSGTRANSMITDONE,
  output [3:0] CFGNEGOTIATEDWIDTH,
  output [1:0] CFGOBFFENABLE,
  output [15:0] CFGPERFUNCSTATUSDATA,
  output CFGPERFUNCTIONUPDATEDONE,
  output CFGPHYLINKDOWN,
  output [1:0] CFGPHYLINKSTATUS,
  output CFGPLSTATUSCHANGE,
  output CFGPOWERSTATECHANGEINTERRUPT,
  output [3:0] CFGRCBSTATUS,
  output [3:0] CFGTPHFUNCTIONNUM,
  output [3:0] CFGTPHREQUESTERENABLE,
  output [11:0] CFGTPHSTMODE,
  output [4:0] CFGTPHSTTADDRESS,
  output CFGTPHSTTREADENABLE,
  output [3:0] CFGTPHSTTWRITEBYTEVALID,
  output [31:0] CFGTPHSTTWRITEDATA,
  output CFGTPHSTTWRITEENABLE,
  output [7:0] CFGVFFLRINPROCESS,
  output [23:0] CFGVFPOWERSTATE,
  output [15:0] CFGVFSTATUS,
  output [7:0] CFGVFTPHREQUESTERENABLE,
  output [23:0] CFGVFTPHSTMODE,
  output CONFMCAPDESIGNSWITCH,
  output CONFMCAPEOS,
  output CONFMCAPINUSEBYPCIE,
  output CONFREQREADY,
  output [31:0] CONFRESPRDATA,
  output CONFRESPVALID,
  output [15:0] DBGDATAOUT,
  output DBGMCAPCSB,
  output [31:0] DBGMCAPDATA,
  output DBGMCAPEOS,
  output DBGMCAPERROR,
  output DBGMCAPMODE,
  output DBGMCAPRDATAVALID,
  output DBGMCAPRDWRB,
  output DBGMCAPRESET,
  output DBGPLDATABLOCKRECEIVEDAFTEREDS,
  output DBGPLGEN3FRAMINGERRORDETECTED,
  output DBGPLGEN3SYNCHEADERERRORDETECTED,
  output [7:0] DBGPLINFERREDRXELECTRICALIDLE,
  output [15:0] DRPDO,
  output DRPRDY,
  output LL2LMMASTERTLPSENT0,
  output LL2LMMASTERTLPSENT1,
  output [3:0] LL2LMMASTERTLPSENTTLPID0,
  output [3:0] LL2LMMASTERTLPSENTTLPID1,
  output [255:0] LL2LMMAXISRXTDATA,
  output [17:0] LL2LMMAXISRXTUSER,
  output [7:0] LL2LMMAXISRXTVALID,
  output [7:0] LL2LMSAXISTXTREADY,
  output [255:0] MAXISCQTDATA,
  output [7:0] MAXISCQTKEEP,
  output MAXISCQTLAST,
  output [84:0] MAXISCQTUSER,
  output MAXISCQTVALID,
  output [255:0] MAXISRCTDATA,
  output [7:0] MAXISRCTKEEP,
  output MAXISRCTLAST,
  output [74:0] MAXISRCTUSER,
  output MAXISRCTVALID,
  output [9:0] MICOMPLETIONRAMREADADDRESSAL,
  output [9:0] MICOMPLETIONRAMREADADDRESSAU,
  output [9:0] MICOMPLETIONRAMREADADDRESSBL,
  output [9:0] MICOMPLETIONRAMREADADDRESSBU,
  output [3:0] MICOMPLETIONRAMREADENABLEL,
  output [3:0] MICOMPLETIONRAMREADENABLEU,
  output [9:0] MICOMPLETIONRAMWRITEADDRESSAL,
  output [9:0] MICOMPLETIONRAMWRITEADDRESSAU,
  output [9:0] MICOMPLETIONRAMWRITEADDRESSBL,
  output [9:0] MICOMPLETIONRAMWRITEADDRESSBU,
  output [71:0] MICOMPLETIONRAMWRITEDATAL,
  output [71:0] MICOMPLETIONRAMWRITEDATAU,
  output [3:0] MICOMPLETIONRAMWRITEENABLEL,
  output [3:0] MICOMPLETIONRAMWRITEENABLEU,
  output [8:0] MIREPLAYRAMADDRESS,
  output [1:0] MIREPLAYRAMREADENABLE,
  output [143:0] MIREPLAYRAMWRITEDATA,
  output [1:0] MIREPLAYRAMWRITEENABLE,
  output [8:0] MIREQUESTRAMREADADDRESSA,
  output [8:0] MIREQUESTRAMREADADDRESSB,
  output [3:0] MIREQUESTRAMREADENABLE,
  output [8:0] MIREQUESTRAMWRITEADDRESSA,
  output [8:0] MIREQUESTRAMWRITEADDRESSB,
  output [143:0] MIREQUESTRAMWRITEDATA,
  output [3:0] MIREQUESTRAMWRITEENABLE,
  output [5:0] PCIECQNPREQCOUNT,
  output PCIEPERST0B,
  output PCIEPERST1B,
  output [3:0] PCIERQSEQNUM,
  output PCIERQSEQNUMVLD,
  output [5:0] PCIERQTAG,
  output [1:0] PCIERQTAGAV,
  output PCIERQTAGVLD,
  output [1:0] PCIETFCNPDAV,
  output [1:0] PCIETFCNPHAV,
  output [1:0] PIPERX0EQCONTROL,
  output [5:0] PIPERX0EQLPLFFS,
  output [3:0] PIPERX0EQLPTXPRESET,
  output [2:0] PIPERX0EQPRESET,
  output PIPERX0POLARITY,
  output [1:0] PIPERX1EQCONTROL,
  output [5:0] PIPERX1EQLPLFFS,
  output [3:0] PIPERX1EQLPTXPRESET,
  output [2:0] PIPERX1EQPRESET,
  output PIPERX1POLARITY,
  output [1:0] PIPERX2EQCONTROL,
  output [5:0] PIPERX2EQLPLFFS,
  output [3:0] PIPERX2EQLPTXPRESET,
  output [2:0] PIPERX2EQPRESET,
  output PIPERX2POLARITY,
  output [1:0] PIPERX3EQCONTROL,
  output [5:0] PIPERX3EQLPLFFS,
  output [3:0] PIPERX3EQLPTXPRESET,
  output [2:0] PIPERX3EQPRESET,
  output PIPERX3POLARITY,
  output [1:0] PIPERX4EQCONTROL,
  output [5:0] PIPERX4EQLPLFFS,
  output [3:0] PIPERX4EQLPTXPRESET,
  output [2:0] PIPERX4EQPRESET,
  output PIPERX4POLARITY,
  output [1:0] PIPERX5EQCONTROL,
  output [5:0] PIPERX5EQLPLFFS,
  output [3:0] PIPERX5EQLPTXPRESET,
  output [2:0] PIPERX5EQPRESET,
  output PIPERX5POLARITY,
  output [1:0] PIPERX6EQCONTROL,
  output [5:0] PIPERX6EQLPLFFS,
  output [3:0] PIPERX6EQLPTXPRESET,
  output [2:0] PIPERX6EQPRESET,
  output PIPERX6POLARITY,
  output [1:0] PIPERX7EQCONTROL,
  output [5:0] PIPERX7EQLPLFFS,
  output [3:0] PIPERX7EQLPTXPRESET,
  output [2:0] PIPERX7EQPRESET,
  output PIPERX7POLARITY,
  output [1:0] PIPETX0CHARISK,
  output PIPETX0COMPLIANCE,
  output [31:0] PIPETX0DATA,
  output PIPETX0DATAVALID,
  output PIPETX0DEEMPH,
  output PIPETX0ELECIDLE,
  output [1:0] PIPETX0EQCONTROL,
  output [5:0] PIPETX0EQDEEMPH,
  output [3:0] PIPETX0EQPRESET,
  output [2:0] PIPETX0MARGIN,
  output [1:0] PIPETX0POWERDOWN,
  output [1:0] PIPETX0RATE,
  output PIPETX0RCVRDET,
  output PIPETX0RESET,
  output PIPETX0STARTBLOCK,
  output PIPETX0SWING,
  output [1:0] PIPETX0SYNCHEADER,
  output [1:0] PIPETX1CHARISK,
  output PIPETX1COMPLIANCE,
  output [31:0] PIPETX1DATA,
  output PIPETX1DATAVALID,
  output PIPETX1DEEMPH,
  output PIPETX1ELECIDLE,
  output [1:0] PIPETX1EQCONTROL,
  output [5:0] PIPETX1EQDEEMPH,
  output [3:0] PIPETX1EQPRESET,
  output [2:0] PIPETX1MARGIN,
  output [1:0] PIPETX1POWERDOWN,
  output [1:0] PIPETX1RATE,
  output PIPETX1RCVRDET,
  output PIPETX1RESET,
  output PIPETX1STARTBLOCK,
  output PIPETX1SWING,
  output [1:0] PIPETX1SYNCHEADER,
  output [1:0] PIPETX2CHARISK,
  output PIPETX2COMPLIANCE,
  output [31:0] PIPETX2DATA,
  output PIPETX2DATAVALID,
  output PIPETX2DEEMPH,
  output PIPETX2ELECIDLE,
  output [1:0] PIPETX2EQCONTROL,
  output [5:0] PIPETX2EQDEEMPH,
  output [3:0] PIPETX2EQPRESET,
  output [2:0] PIPETX2MARGIN,
  output [1:0] PIPETX2POWERDOWN,
  output [1:0] PIPETX2RATE,
  output PIPETX2RCVRDET,
  output PIPETX2RESET,
  output PIPETX2STARTBLOCK,
  output PIPETX2SWING,
  output [1:0] PIPETX2SYNCHEADER,
  output [1:0] PIPETX3CHARISK,
  output PIPETX3COMPLIANCE,
  output [31:0] PIPETX3DATA,
  output PIPETX3DATAVALID,
  output PIPETX3DEEMPH,
  output PIPETX3ELECIDLE,
  output [1:0] PIPETX3EQCONTROL,
  output [5:0] PIPETX3EQDEEMPH,
  output [3:0] PIPETX3EQPRESET,
  output [2:0] PIPETX3MARGIN,
  output [1:0] PIPETX3POWERDOWN,
  output [1:0] PIPETX3RATE,
  output PIPETX3RCVRDET,
  output PIPETX3RESET,
  output PIPETX3STARTBLOCK,
  output PIPETX3SWING,
  output [1:0] PIPETX3SYNCHEADER,
  output [1:0] PIPETX4CHARISK,
  output PIPETX4COMPLIANCE,
  output [31:0] PIPETX4DATA,
  output PIPETX4DATAVALID,
  output PIPETX4DEEMPH,
  output PIPETX4ELECIDLE,
  output [1:0] PIPETX4EQCONTROL,
  output [5:0] PIPETX4EQDEEMPH,
  output [3:0] PIPETX4EQPRESET,
  output [2:0] PIPETX4MARGIN,
  output [1:0] PIPETX4POWERDOWN,
  output [1:0] PIPETX4RATE,
  output PIPETX4RCVRDET,
  output PIPETX4RESET,
  output PIPETX4STARTBLOCK,
  output PIPETX4SWING,
  output [1:0] PIPETX4SYNCHEADER,
  output [1:0] PIPETX5CHARISK,
  output PIPETX5COMPLIANCE,
  output [31:0] PIPETX5DATA,
  output PIPETX5DATAVALID,
  output PIPETX5DEEMPH,
  output PIPETX5ELECIDLE,
  output [1:0] PIPETX5EQCONTROL,
  output [5:0] PIPETX5EQDEEMPH,
  output [3:0] PIPETX5EQPRESET,
  output [2:0] PIPETX5MARGIN,
  output [1:0] PIPETX5POWERDOWN,
  output [1:0] PIPETX5RATE,
  output PIPETX5RCVRDET,
  output PIPETX5RESET,
  output PIPETX5STARTBLOCK,
  output PIPETX5SWING,
  output [1:0] PIPETX5SYNCHEADER,
  output [1:0] PIPETX6CHARISK,
  output PIPETX6COMPLIANCE,
  output [31:0] PIPETX6DATA,
  output PIPETX6DATAVALID,
  output PIPETX6DEEMPH,
  output PIPETX6ELECIDLE,
  output [1:0] PIPETX6EQCONTROL,
  output [5:0] PIPETX6EQDEEMPH,
  output [3:0] PIPETX6EQPRESET,
  output [2:0] PIPETX6MARGIN,
  output [1:0] PIPETX6POWERDOWN,
  output [1:0] PIPETX6RATE,
  output PIPETX6RCVRDET,
  output PIPETX6RESET,
  output PIPETX6STARTBLOCK,
  output PIPETX6SWING,
  output [1:0] PIPETX6SYNCHEADER,
  output [1:0] PIPETX7CHARISK,
  output PIPETX7COMPLIANCE,
  output [31:0] PIPETX7DATA,
  output PIPETX7DATAVALID,
  output PIPETX7DEEMPH,
  output PIPETX7ELECIDLE,
  output [1:0] PIPETX7EQCONTROL,
  output [5:0] PIPETX7EQDEEMPH,
  output [3:0] PIPETX7EQPRESET,
  output [2:0] PIPETX7MARGIN,
  output [1:0] PIPETX7POWERDOWN,
  output [1:0] PIPETX7RATE,
  output PIPETX7RCVRDET,
  output PIPETX7RESET,
  output PIPETX7STARTBLOCK,
  output PIPETX7SWING,
  output [1:0] PIPETX7SYNCHEADER,
  output PLEQINPROGRESS,
  output [1:0] PLEQPHASE,
  output [3:0] SAXISCCTREADY,
  output [3:0] SAXISRQTREADY,
  output [31:0] SPAREOUT,

  input CFGCONFIGSPACEENABLE,
  input [15:0] CFGDEVID,
  input [7:0] CFGDSBUSNUMBER,
  input [4:0] CFGDSDEVICENUMBER,
  input [2:0] CFGDSFUNCTIONNUMBER,
  input [63:0] CFGDSN,
  input [7:0] CFGDSPORTNUMBER,
  input CFGERRCORIN,
  input CFGERRUNCORIN,
  input [31:0] CFGEXTREADDATA,
  input CFGEXTREADDATAVALID,
  input [2:0] CFGFCSEL,
  input [3:0] CFGFLRDONE,
  input CFGHOTRESETIN,
  input [3:0] CFGINTERRUPTINT,
  input [2:0] CFGINTERRUPTMSIATTR,
  input [3:0] CFGINTERRUPTMSIFUNCTIONNUMBER,
  input [31:0] CFGINTERRUPTMSIINT,
  input [31:0] CFGINTERRUPTMSIPENDINGSTATUS,
  input CFGINTERRUPTMSIPENDINGSTATUSDATAENABLE,
  input [3:0] CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM,
  input [3:0] CFGINTERRUPTMSISELECT,
  input CFGINTERRUPTMSITPHPRESENT,
  input [8:0] CFGINTERRUPTMSITPHSTTAG,
  input [1:0] CFGINTERRUPTMSITPHTYPE,
  input [63:0] CFGINTERRUPTMSIXADDRESS,
  input [31:0] CFGINTERRUPTMSIXDATA,
  input CFGINTERRUPTMSIXINT,
  input [3:0] CFGINTERRUPTPENDING,
  input CFGLINKTRAININGENABLE,
  input [18:0] CFGMGMTADDR,
  input [3:0] CFGMGMTBYTEENABLE,
  input CFGMGMTREAD,
  input CFGMGMTTYPE1CFGREGACCESS,
  input CFGMGMTWRITE,
  input [31:0] CFGMGMTWRITEDATA,
  input CFGMSGTRANSMIT,
  input [31:0] CFGMSGTRANSMITDATA,
  input [2:0] CFGMSGTRANSMITTYPE,
  input [2:0] CFGPERFUNCSTATUSCONTROL,
  input [3:0] CFGPERFUNCTIONNUMBER,
  input CFGPERFUNCTIONOUTPUTREQUEST,
  input CFGPOWERSTATECHANGEACK,
  input CFGREQPMTRANSITIONL23READY,
  input [7:0] CFGREVID,
  input [15:0] CFGSUBSYSID,
  input [15:0] CFGSUBSYSVENDID,
  input [31:0] CFGTPHSTTREADDATA,
  input CFGTPHSTTREADDATAVALID,
  input [15:0] CFGVENDID,
  input [7:0] CFGVFFLRDONE,
  input CONFMCAPREQUESTBYCONF,
  input [31:0] CONFREQDATA,
  input [3:0] CONFREQREGNUM,
  input [1:0] CONFREQTYPE,
  input CONFREQVALID,
  input CORECLK,
  input CORECLKMICOMPLETIONRAML,
  input CORECLKMICOMPLETIONRAMU,
  input CORECLKMIREPLAYRAM,
  input CORECLKMIREQUESTRAM,
  input DBGCFGLOCALMGMTREGOVERRIDE,
  input [3:0] DBGDATASEL,
  input [9:0] DRPADDR,
  input DRPCLK,
  input [15:0] DRPDI,
  input DRPEN,
  input DRPWE,
  input [13:0] LL2LMSAXISTXTUSER,
  input LL2LMSAXISTXTVALID,
  input [3:0] LL2LMTXTLPID0,
  input [3:0] LL2LMTXTLPID1,
  input [21:0] MAXISCQTREADY,
  input [21:0] MAXISRCTREADY,
  input MCAPCLK,
  input MCAPPERST0B,
  input MCAPPERST1B,
  input MGMTRESETN,
  input MGMTSTICKYRESETN,
  input [143:0] MICOMPLETIONRAMREADDATA,
  input [143:0] MIREPLAYRAMREADDATA,
  input [143:0] MIREQUESTRAMREADDATA,
  input PCIECQNPREQ,
  input PIPECLK,
  input [5:0] PIPEEQFS,
  input [5:0] PIPEEQLF,
  input PIPERESETN,
  input [1:0] PIPERX0CHARISK,
  input [31:0] PIPERX0DATA,
  input PIPERX0DATAVALID,
  input PIPERX0ELECIDLE,
  input PIPERX0EQDONE,
  input PIPERX0EQLPADAPTDONE,
  input PIPERX0EQLPLFFSSEL,
  input [17:0] PIPERX0EQLPNEWTXCOEFFORPRESET,
  input PIPERX0PHYSTATUS,
  input PIPERX0STARTBLOCK,
  input [2:0] PIPERX0STATUS,
  input [1:0] PIPERX0SYNCHEADER,
  input PIPERX0VALID,
  input [1:0] PIPERX1CHARISK,
  input [31:0] PIPERX1DATA,
  input PIPERX1DATAVALID,
  input PIPERX1ELECIDLE,
  input PIPERX1EQDONE,
  input PIPERX1EQLPADAPTDONE,
  input PIPERX1EQLPLFFSSEL,
  input [17:0] PIPERX1EQLPNEWTXCOEFFORPRESET,
  input PIPERX1PHYSTATUS,
  input PIPERX1STARTBLOCK,
  input [2:0] PIPERX1STATUS,
  input [1:0] PIPERX1SYNCHEADER,
  input PIPERX1VALID,
  input [1:0] PIPERX2CHARISK,
  input [31:0] PIPERX2DATA,
  input PIPERX2DATAVALID,
  input PIPERX2ELECIDLE,
  input PIPERX2EQDONE,
  input PIPERX2EQLPADAPTDONE,
  input PIPERX2EQLPLFFSSEL,
  input [17:0] PIPERX2EQLPNEWTXCOEFFORPRESET,
  input PIPERX2PHYSTATUS,
  input PIPERX2STARTBLOCK,
  input [2:0] PIPERX2STATUS,
  input [1:0] PIPERX2SYNCHEADER,
  input PIPERX2VALID,
  input [1:0] PIPERX3CHARISK,
  input [31:0] PIPERX3DATA,
  input PIPERX3DATAVALID,
  input PIPERX3ELECIDLE,
  input PIPERX3EQDONE,
  input PIPERX3EQLPADAPTDONE,
  input PIPERX3EQLPLFFSSEL,
  input [17:0] PIPERX3EQLPNEWTXCOEFFORPRESET,
  input PIPERX3PHYSTATUS,
  input PIPERX3STARTBLOCK,
  input [2:0] PIPERX3STATUS,
  input [1:0] PIPERX3SYNCHEADER,
  input PIPERX3VALID,
  input [1:0] PIPERX4CHARISK,
  input [31:0] PIPERX4DATA,
  input PIPERX4DATAVALID,
  input PIPERX4ELECIDLE,
  input PIPERX4EQDONE,
  input PIPERX4EQLPADAPTDONE,
  input PIPERX4EQLPLFFSSEL,
  input [17:0] PIPERX4EQLPNEWTXCOEFFORPRESET,
  input PIPERX4PHYSTATUS,
  input PIPERX4STARTBLOCK,
  input [2:0] PIPERX4STATUS,
  input [1:0] PIPERX4SYNCHEADER,
  input PIPERX4VALID,
  input [1:0] PIPERX5CHARISK,
  input [31:0] PIPERX5DATA,
  input PIPERX5DATAVALID,
  input PIPERX5ELECIDLE,
  input PIPERX5EQDONE,
  input PIPERX5EQLPADAPTDONE,
  input PIPERX5EQLPLFFSSEL,
  input [17:0] PIPERX5EQLPNEWTXCOEFFORPRESET,
  input PIPERX5PHYSTATUS,
  input PIPERX5STARTBLOCK,
  input [2:0] PIPERX5STATUS,
  input [1:0] PIPERX5SYNCHEADER,
  input PIPERX5VALID,
  input [1:0] PIPERX6CHARISK,
  input [31:0] PIPERX6DATA,
  input PIPERX6DATAVALID,
  input PIPERX6ELECIDLE,
  input PIPERX6EQDONE,
  input PIPERX6EQLPADAPTDONE,
  input PIPERX6EQLPLFFSSEL,
  input [17:0] PIPERX6EQLPNEWTXCOEFFORPRESET,
  input PIPERX6PHYSTATUS,
  input PIPERX6STARTBLOCK,
  input [2:0] PIPERX6STATUS,
  input [1:0] PIPERX6SYNCHEADER,
  input PIPERX6VALID,
  input [1:0] PIPERX7CHARISK,
  input [31:0] PIPERX7DATA,
  input PIPERX7DATAVALID,
  input PIPERX7ELECIDLE,
  input PIPERX7EQDONE,
  input PIPERX7EQLPADAPTDONE,
  input PIPERX7EQLPLFFSSEL,
  input [17:0] PIPERX7EQLPNEWTXCOEFFORPRESET,
  input PIPERX7PHYSTATUS,
  input PIPERX7STARTBLOCK,
  input [2:0] PIPERX7STATUS,
  input [1:0] PIPERX7SYNCHEADER,
  input PIPERX7VALID,
  input [17:0] PIPETX0EQCOEFF,
  input PIPETX0EQDONE,
  input [17:0] PIPETX1EQCOEFF,
  input PIPETX1EQDONE,
  input [17:0] PIPETX2EQCOEFF,
  input PIPETX2EQDONE,
  input [17:0] PIPETX3EQCOEFF,
  input PIPETX3EQDONE,
  input [17:0] PIPETX4EQCOEFF,
  input PIPETX4EQDONE,
  input [17:0] PIPETX5EQCOEFF,
  input PIPETX5EQDONE,
  input [17:0] PIPETX6EQCOEFF,
  input PIPETX6EQDONE,
  input [17:0] PIPETX7EQCOEFF,
  input PIPETX7EQDONE,
  input PLEQRESETEIEOSCOUNT,
  input PLGEN2UPSTREAMPREFERDEEMPH,
  input RESETN,
  input [255:0] SAXISCCTDATA,
  input [7:0] SAXISCCTKEEP,
  input SAXISCCTLAST,
  input [32:0] SAXISCCTUSER,
  input SAXISCCTVALID,
  input [255:0] SAXISRQTDATA,
  input [7:0] SAXISRQTKEEP,
  input SAXISRQTLAST,
  input [59:0] SAXISRQTUSER,
  input SAXISRQTVALID,
  input [31:0] SPAREIN,
  input USERCLK
);
  
// define constants
  localparam MODULE_NAME = "PCIE_3_1";
  localparam in_delay    = 0;
  localparam out_delay   = 0;
  localparam inclk_delay    = 0;
  localparam outclk_delay   = 0;

// Parameter encodings and registers

  `ifndef XIL_DR
  localparam [40:1] ARI_CAP_ENABLE_REG = ARI_CAP_ENABLE;
  localparam [40:1] AXISTEN_IF_CC_ALIGNMENT_MODE_REG = AXISTEN_IF_CC_ALIGNMENT_MODE;
  localparam [40:1] AXISTEN_IF_CC_PARITY_CHK_REG = AXISTEN_IF_CC_PARITY_CHK;
  localparam [40:1] AXISTEN_IF_CQ_ALIGNMENT_MODE_REG = AXISTEN_IF_CQ_ALIGNMENT_MODE;
  localparam [40:1] AXISTEN_IF_ENABLE_CLIENT_TAG_REG = AXISTEN_IF_ENABLE_CLIENT_TAG;
  localparam [17:0] AXISTEN_IF_ENABLE_MSG_ROUTE_REG = AXISTEN_IF_ENABLE_MSG_ROUTE;
  localparam [40:1] AXISTEN_IF_ENABLE_RX_MSG_INTFC_REG = AXISTEN_IF_ENABLE_RX_MSG_INTFC;
  localparam [40:1] AXISTEN_IF_RC_ALIGNMENT_MODE_REG = AXISTEN_IF_RC_ALIGNMENT_MODE;
  localparam [40:1] AXISTEN_IF_RC_STRADDLE_REG = AXISTEN_IF_RC_STRADDLE;
  localparam [40:1] AXISTEN_IF_RQ_ALIGNMENT_MODE_REG = AXISTEN_IF_RQ_ALIGNMENT_MODE;
  localparam [40:1] AXISTEN_IF_RQ_PARITY_CHK_REG = AXISTEN_IF_RQ_PARITY_CHK;
  localparam [1:0] AXISTEN_IF_WIDTH_REG = AXISTEN_IF_WIDTH;
  localparam [40:1] CRM_CORE_CLK_FREQ_500_REG = CRM_CORE_CLK_FREQ_500;
  localparam [1:0] CRM_USER_CLK_FREQ_REG = CRM_USER_CLK_FREQ;
  localparam [40:1] DEBUG_CFG_LOCAL_MGMT_REG_ACCESS_OVERRIDE_REG = DEBUG_CFG_LOCAL_MGMT_REG_ACCESS_OVERRIDE;
  localparam [40:1] DEBUG_PL_DISABLE_EI_INFER_IN_L0_REG = DEBUG_PL_DISABLE_EI_INFER_IN_L0;
  localparam [40:1] DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS_REG = DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS;
  localparam [7:0] DNSTREAM_LINK_NUM_REG = DNSTREAM_LINK_NUM;
  localparam [8:0] LL_ACK_TIMEOUT_REG = LL_ACK_TIMEOUT;
  localparam [40:1] LL_ACK_TIMEOUT_EN_REG = LL_ACK_TIMEOUT_EN;
  localparam [1:0] LL_ACK_TIMEOUT_FUNC_REG = LL_ACK_TIMEOUT_FUNC;
  localparam [15:0] LL_CPL_FC_UPDATE_TIMER_REG = LL_CPL_FC_UPDATE_TIMER;
  localparam [40:1] LL_CPL_FC_UPDATE_TIMER_OVERRIDE_REG = LL_CPL_FC_UPDATE_TIMER_OVERRIDE;
  localparam [15:0] LL_FC_UPDATE_TIMER_REG = LL_FC_UPDATE_TIMER;
  localparam [40:1] LL_FC_UPDATE_TIMER_OVERRIDE_REG = LL_FC_UPDATE_TIMER_OVERRIDE;
  localparam [15:0] LL_NP_FC_UPDATE_TIMER_REG = LL_NP_FC_UPDATE_TIMER;
  localparam [40:1] LL_NP_FC_UPDATE_TIMER_OVERRIDE_REG = LL_NP_FC_UPDATE_TIMER_OVERRIDE;
  localparam [15:0] LL_P_FC_UPDATE_TIMER_REG = LL_P_FC_UPDATE_TIMER;
  localparam [40:1] LL_P_FC_UPDATE_TIMER_OVERRIDE_REG = LL_P_FC_UPDATE_TIMER_OVERRIDE;
  localparam [8:0] LL_REPLAY_TIMEOUT_REG = LL_REPLAY_TIMEOUT;
  localparam [40:1] LL_REPLAY_TIMEOUT_EN_REG = LL_REPLAY_TIMEOUT_EN;
  localparam [1:0] LL_REPLAY_TIMEOUT_FUNC_REG = LL_REPLAY_TIMEOUT_FUNC;
  localparam [9:0] LTR_TX_MESSAGE_MINIMUM_INTERVAL_REG = LTR_TX_MESSAGE_MINIMUM_INTERVAL;
  localparam [40:1] LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE_REG = LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE;
  localparam [40:1] LTR_TX_MESSAGE_ON_LTR_ENABLE_REG = LTR_TX_MESSAGE_ON_LTR_ENABLE;
  localparam [11:0] MCAP_CAP_NEXTPTR_REG = MCAP_CAP_NEXTPTR;
  localparam [40:1] MCAP_CONFIGURE_OVERRIDE_REG = MCAP_CONFIGURE_OVERRIDE;
  localparam [40:1] MCAP_ENABLE_REG = MCAP_ENABLE;
  localparam [40:1] MCAP_EOS_DESIGN_SWITCH_REG = MCAP_EOS_DESIGN_SWITCH;
  localparam [31:0] MCAP_FPGA_BITSTREAM_VERSION_REG = MCAP_FPGA_BITSTREAM_VERSION;
  localparam [40:1] MCAP_GATE_IO_ENABLE_DESIGN_SWITCH_REG = MCAP_GATE_IO_ENABLE_DESIGN_SWITCH;
  localparam [40:1] MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH_REG = MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH;
  localparam [40:1] MCAP_INPUT_GATE_DESIGN_SWITCH_REG = MCAP_INPUT_GATE_DESIGN_SWITCH;
  localparam [40:1] MCAP_INTERRUPT_ON_MCAP_EOS_REG = MCAP_INTERRUPT_ON_MCAP_EOS;
  localparam [40:1] MCAP_INTERRUPT_ON_MCAP_ERROR_REG = MCAP_INTERRUPT_ON_MCAP_ERROR;
  localparam [15:0] MCAP_VSEC_ID_REG = MCAP_VSEC_ID;
  localparam [11:0] MCAP_VSEC_LEN_REG = MCAP_VSEC_LEN;
  localparam [3:0] MCAP_VSEC_REV_REG = MCAP_VSEC_REV;
  localparam [40:1] PF0_AER_CAP_ECRC_CHECK_CAPABLE_REG = PF0_AER_CAP_ECRC_CHECK_CAPABLE;
  localparam [40:1] PF0_AER_CAP_ECRC_GEN_CAPABLE_REG = PF0_AER_CAP_ECRC_GEN_CAPABLE;
  localparam [11:0] PF0_AER_CAP_NEXTPTR_REG = PF0_AER_CAP_NEXTPTR;
  localparam [11:0] PF0_ARI_CAP_NEXTPTR_REG = PF0_ARI_CAP_NEXTPTR;
  localparam [7:0] PF0_ARI_CAP_NEXT_FUNC_REG = PF0_ARI_CAP_NEXT_FUNC;
  localparam [3:0] PF0_ARI_CAP_VER_REG = PF0_ARI_CAP_VER;
  localparam [5:0] PF0_BAR0_APERTURE_SIZE_REG = PF0_BAR0_APERTURE_SIZE;
  localparam [2:0] PF0_BAR0_CONTROL_REG = PF0_BAR0_CONTROL;
  localparam [5:0] PF0_BAR1_APERTURE_SIZE_REG = PF0_BAR1_APERTURE_SIZE;
  localparam [2:0] PF0_BAR1_CONTROL_REG = PF0_BAR1_CONTROL;
  localparam [4:0] PF0_BAR2_APERTURE_SIZE_REG = PF0_BAR2_APERTURE_SIZE;
  localparam [2:0] PF0_BAR2_CONTROL_REG = PF0_BAR2_CONTROL;
  localparam [4:0] PF0_BAR3_APERTURE_SIZE_REG = PF0_BAR3_APERTURE_SIZE;
  localparam [2:0] PF0_BAR3_CONTROL_REG = PF0_BAR3_CONTROL;
  localparam [4:0] PF0_BAR4_APERTURE_SIZE_REG = PF0_BAR4_APERTURE_SIZE;
  localparam [2:0] PF0_BAR4_CONTROL_REG = PF0_BAR4_CONTROL;
  localparam [4:0] PF0_BAR5_APERTURE_SIZE_REG = PF0_BAR5_APERTURE_SIZE;
  localparam [2:0] PF0_BAR5_CONTROL_REG = PF0_BAR5_CONTROL;
  localparam [7:0] PF0_BIST_REGISTER_REG = PF0_BIST_REGISTER;
  localparam [7:0] PF0_CAPABILITY_POINTER_REG = PF0_CAPABILITY_POINTER;
  localparam [23:0] PF0_CLASS_CODE_REG = PF0_CLASS_CODE;
  localparam [15:0] PF0_DEVICE_ID_REG = PF0_DEVICE_ID;
  localparam [40:1] PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT_REG = PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT;
  localparam [40:1] PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT_REG = PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT;
  localparam [40:1] PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT_REG = PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT;
  localparam [40:1] PF0_DEV_CAP2_ARI_FORWARD_ENABLE_REG = PF0_DEV_CAP2_ARI_FORWARD_ENABLE;
  localparam [40:1] PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE_REG = PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE;
  localparam [40:1] PF0_DEV_CAP2_LTR_SUPPORT_REG = PF0_DEV_CAP2_LTR_SUPPORT;
  localparam [1:0] PF0_DEV_CAP2_OBFF_SUPPORT_REG = PF0_DEV_CAP2_OBFF_SUPPORT;
  localparam [40:1] PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT_REG = PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT;
  localparam [2:0] PF0_DEV_CAP_ENDPOINT_L0S_LATENCY_REG = PF0_DEV_CAP_ENDPOINT_L0S_LATENCY;
  localparam [2:0] PF0_DEV_CAP_ENDPOINT_L1_LATENCY_REG = PF0_DEV_CAP_ENDPOINT_L1_LATENCY;
  localparam [40:1] PF0_DEV_CAP_EXT_TAG_SUPPORTED_REG = PF0_DEV_CAP_EXT_TAG_SUPPORTED;
  localparam [40:1] PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE_REG = PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE;
  localparam [2:0] PF0_DEV_CAP_MAX_PAYLOAD_SIZE_REG = PF0_DEV_CAP_MAX_PAYLOAD_SIZE;
  localparam [11:0] PF0_DPA_CAP_NEXTPTR_REG = PF0_DPA_CAP_NEXTPTR;
  localparam [4:0] PF0_DPA_CAP_SUB_STATE_CONTROL_REG = PF0_DPA_CAP_SUB_STATE_CONTROL;
  localparam [40:1] PF0_DPA_CAP_SUB_STATE_CONTROL_EN_REG = PF0_DPA_CAP_SUB_STATE_CONTROL_EN;
  localparam [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION0_REG = PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION0;
  localparam [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION1_REG = PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION1;
  localparam [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION2_REG = PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION2;
  localparam [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION3_REG = PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION3;
  localparam [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION4_REG = PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION4;
  localparam [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION5_REG = PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION5;
  localparam [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION6_REG = PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION6;
  localparam [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION7_REG = PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION7;
  localparam [3:0] PF0_DPA_CAP_VER_REG = PF0_DPA_CAP_VER;
  localparam [11:0] PF0_DSN_CAP_NEXTPTR_REG = PF0_DSN_CAP_NEXTPTR;
  localparam [4:0] PF0_EXPANSION_ROM_APERTURE_SIZE_REG = PF0_EXPANSION_ROM_APERTURE_SIZE;
  localparam [40:1] PF0_EXPANSION_ROM_ENABLE_REG = PF0_EXPANSION_ROM_ENABLE;
  localparam [7:0] PF0_INTERRUPT_LINE_REG = PF0_INTERRUPT_LINE;
  localparam [2:0] PF0_INTERRUPT_PIN_REG = PF0_INTERRUPT_PIN;
  localparam [1:0] PF0_LINK_CAP_ASPM_SUPPORT_REG = PF0_LINK_CAP_ASPM_SUPPORT;
  localparam [2:0] PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1_REG = PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1;
  localparam [2:0] PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2_REG = PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2;
  localparam [2:0] PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3_REG = PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3;
  localparam [2:0] PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1_REG = PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1;
  localparam [2:0] PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2_REG = PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2;
  localparam [2:0] PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3_REG = PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3;
  localparam [2:0] PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1_REG = PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1;
  localparam [2:0] PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2_REG = PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2;
  localparam [2:0] PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3_REG = PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3;
  localparam [2:0] PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1_REG = PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1;
  localparam [2:0] PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2_REG = PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2;
  localparam [2:0] PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3_REG = PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3;
  localparam [40:1] PF0_LINK_STATUS_SLOT_CLOCK_CONFIG_REG = PF0_LINK_STATUS_SLOT_CLOCK_CONFIG;
  localparam [9:0] PF0_LTR_CAP_MAX_NOSNOOP_LAT_REG = PF0_LTR_CAP_MAX_NOSNOOP_LAT;
  localparam [9:0] PF0_LTR_CAP_MAX_SNOOP_LAT_REG = PF0_LTR_CAP_MAX_SNOOP_LAT;
  localparam [11:0] PF0_LTR_CAP_NEXTPTR_REG = PF0_LTR_CAP_NEXTPTR;
  localparam [3:0] PF0_LTR_CAP_VER_REG = PF0_LTR_CAP_VER;
  localparam [7:0] PF0_MSIX_CAP_NEXTPTR_REG = PF0_MSIX_CAP_NEXTPTR;
  localparam [2:0] PF0_MSIX_CAP_PBA_BIR_REG = PF0_MSIX_CAP_PBA_BIR;
  localparam [28:0] PF0_MSIX_CAP_PBA_OFFSET_REG = PF0_MSIX_CAP_PBA_OFFSET;
  localparam [2:0] PF0_MSIX_CAP_TABLE_BIR_REG = PF0_MSIX_CAP_TABLE_BIR;
  localparam [28:0] PF0_MSIX_CAP_TABLE_OFFSET_REG = PF0_MSIX_CAP_TABLE_OFFSET;
  localparam [10:0] PF0_MSIX_CAP_TABLE_SIZE_REG = PF0_MSIX_CAP_TABLE_SIZE;
  localparam [2:0] PF0_MSI_CAP_MULTIMSGCAP_REG = PF0_MSI_CAP_MULTIMSGCAP;
  localparam [7:0] PF0_MSI_CAP_NEXTPTR_REG = PF0_MSI_CAP_NEXTPTR;
  localparam [40:1] PF0_MSI_CAP_PERVECMASKCAP_REG = PF0_MSI_CAP_PERVECMASKCAP;
  localparam [31:0] PF0_PB_CAP_DATA_REG_D0_REG = PF0_PB_CAP_DATA_REG_D0;
  localparam [31:0] PF0_PB_CAP_DATA_REG_D0_SUSTAINED_REG = PF0_PB_CAP_DATA_REG_D0_SUSTAINED;
  localparam [31:0] PF0_PB_CAP_DATA_REG_D1_REG = PF0_PB_CAP_DATA_REG_D1;
  localparam [31:0] PF0_PB_CAP_DATA_REG_D3HOT_REG = PF0_PB_CAP_DATA_REG_D3HOT;
  localparam [11:0] PF0_PB_CAP_NEXTPTR_REG = PF0_PB_CAP_NEXTPTR;
  localparam [40:1] PF0_PB_CAP_SYSTEM_ALLOCATED_REG = PF0_PB_CAP_SYSTEM_ALLOCATED;
  localparam [3:0] PF0_PB_CAP_VER_REG = PF0_PB_CAP_VER;
  localparam [7:0] PF0_PM_CAP_ID_REG = PF0_PM_CAP_ID;
  localparam [7:0] PF0_PM_CAP_NEXTPTR_REG = PF0_PM_CAP_NEXTPTR;
  localparam [40:1] PF0_PM_CAP_PMESUPPORT_D0_REG = PF0_PM_CAP_PMESUPPORT_D0;
  localparam [40:1] PF0_PM_CAP_PMESUPPORT_D1_REG = PF0_PM_CAP_PMESUPPORT_D1;
  localparam [40:1] PF0_PM_CAP_PMESUPPORT_D3HOT_REG = PF0_PM_CAP_PMESUPPORT_D3HOT;
  localparam [40:1] PF0_PM_CAP_SUPP_D1_STATE_REG = PF0_PM_CAP_SUPP_D1_STATE;
  localparam [2:0] PF0_PM_CAP_VER_ID_REG = PF0_PM_CAP_VER_ID;
  localparam [40:1] PF0_PM_CSR_NOSOFTRESET_REG = PF0_PM_CSR_NOSOFTRESET;
  localparam [40:1] PF0_RBAR_CAP_ENABLE_REG = PF0_RBAR_CAP_ENABLE;
  localparam [11:0] PF0_RBAR_CAP_NEXTPTR_REG = PF0_RBAR_CAP_NEXTPTR;
  localparam [19:0] PF0_RBAR_CAP_SIZE0_REG = PF0_RBAR_CAP_SIZE0;
  localparam [19:0] PF0_RBAR_CAP_SIZE1_REG = PF0_RBAR_CAP_SIZE1;
  localparam [19:0] PF0_RBAR_CAP_SIZE2_REG = PF0_RBAR_CAP_SIZE2;
  localparam [3:0] PF0_RBAR_CAP_VER_REG = PF0_RBAR_CAP_VER;
  localparam [2:0] PF0_RBAR_CONTROL_INDEX0_REG = PF0_RBAR_CONTROL_INDEX0;
  localparam [2:0] PF0_RBAR_CONTROL_INDEX1_REG = PF0_RBAR_CONTROL_INDEX1;
  localparam [2:0] PF0_RBAR_CONTROL_INDEX2_REG = PF0_RBAR_CONTROL_INDEX2;
  localparam [4:0] PF0_RBAR_CONTROL_SIZE0_REG = PF0_RBAR_CONTROL_SIZE0;
  localparam [4:0] PF0_RBAR_CONTROL_SIZE1_REG = PF0_RBAR_CONTROL_SIZE1;
  localparam [4:0] PF0_RBAR_CONTROL_SIZE2_REG = PF0_RBAR_CONTROL_SIZE2;
  localparam [2:0] PF0_RBAR_NUM_REG = PF0_RBAR_NUM;
  localparam [7:0] PF0_REVISION_ID_REG = PF0_REVISION_ID;
  localparam [11:0] PF0_SECONDARY_PCIE_CAP_NEXTPTR_REG = PF0_SECONDARY_PCIE_CAP_NEXTPTR;
  localparam [4:0] PF0_SRIOV_BAR0_APERTURE_SIZE_REG = PF0_SRIOV_BAR0_APERTURE_SIZE;
  localparam [2:0] PF0_SRIOV_BAR0_CONTROL_REG = PF0_SRIOV_BAR0_CONTROL;
  localparam [4:0] PF0_SRIOV_BAR1_APERTURE_SIZE_REG = PF0_SRIOV_BAR1_APERTURE_SIZE;
  localparam [2:0] PF0_SRIOV_BAR1_CONTROL_REG = PF0_SRIOV_BAR1_CONTROL;
  localparam [4:0] PF0_SRIOV_BAR2_APERTURE_SIZE_REG = PF0_SRIOV_BAR2_APERTURE_SIZE;
  localparam [2:0] PF0_SRIOV_BAR2_CONTROL_REG = PF0_SRIOV_BAR2_CONTROL;
  localparam [4:0] PF0_SRIOV_BAR3_APERTURE_SIZE_REG = PF0_SRIOV_BAR3_APERTURE_SIZE;
  localparam [2:0] PF0_SRIOV_BAR3_CONTROL_REG = PF0_SRIOV_BAR3_CONTROL;
  localparam [4:0] PF0_SRIOV_BAR4_APERTURE_SIZE_REG = PF0_SRIOV_BAR4_APERTURE_SIZE;
  localparam [2:0] PF0_SRIOV_BAR4_CONTROL_REG = PF0_SRIOV_BAR4_CONTROL;
  localparam [4:0] PF0_SRIOV_BAR5_APERTURE_SIZE_REG = PF0_SRIOV_BAR5_APERTURE_SIZE;
  localparam [2:0] PF0_SRIOV_BAR5_CONTROL_REG = PF0_SRIOV_BAR5_CONTROL;
  localparam [15:0] PF0_SRIOV_CAP_INITIAL_VF_REG = PF0_SRIOV_CAP_INITIAL_VF;
  localparam [11:0] PF0_SRIOV_CAP_NEXTPTR_REG = PF0_SRIOV_CAP_NEXTPTR;
  localparam [15:0] PF0_SRIOV_CAP_TOTAL_VF_REG = PF0_SRIOV_CAP_TOTAL_VF;
  localparam [3:0] PF0_SRIOV_CAP_VER_REG = PF0_SRIOV_CAP_VER;
  localparam [15:0] PF0_SRIOV_FIRST_VF_OFFSET_REG = PF0_SRIOV_FIRST_VF_OFFSET;
  localparam [15:0] PF0_SRIOV_FUNC_DEP_LINK_REG = PF0_SRIOV_FUNC_DEP_LINK;
  localparam [31:0] PF0_SRIOV_SUPPORTED_PAGE_SIZE_REG = PF0_SRIOV_SUPPORTED_PAGE_SIZE;
  localparam [15:0] PF0_SRIOV_VF_DEVICE_ID_REG = PF0_SRIOV_VF_DEVICE_ID;
  localparam [15:0] PF0_SUBSYSTEM_ID_REG = PF0_SUBSYSTEM_ID;
  localparam [40:1] PF0_TPHR_CAP_DEV_SPECIFIC_MODE_REG = PF0_TPHR_CAP_DEV_SPECIFIC_MODE;
  localparam [40:1] PF0_TPHR_CAP_ENABLE_REG = PF0_TPHR_CAP_ENABLE;
  localparam [40:1] PF0_TPHR_CAP_INT_VEC_MODE_REG = PF0_TPHR_CAP_INT_VEC_MODE;
  localparam [11:0] PF0_TPHR_CAP_NEXTPTR_REG = PF0_TPHR_CAP_NEXTPTR;
  localparam [2:0] PF0_TPHR_CAP_ST_MODE_SEL_REG = PF0_TPHR_CAP_ST_MODE_SEL;
  localparam [1:0] PF0_TPHR_CAP_ST_TABLE_LOC_REG = PF0_TPHR_CAP_ST_TABLE_LOC;
  localparam [10:0] PF0_TPHR_CAP_ST_TABLE_SIZE_REG = PF0_TPHR_CAP_ST_TABLE_SIZE;
  localparam [3:0] PF0_TPHR_CAP_VER_REG = PF0_TPHR_CAP_VER;
  localparam [40:1] PF0_VC_CAP_ENABLE_REG = PF0_VC_CAP_ENABLE;
  localparam [11:0] PF0_VC_CAP_NEXTPTR_REG = PF0_VC_CAP_NEXTPTR;
  localparam [3:0] PF0_VC_CAP_VER_REG = PF0_VC_CAP_VER;
  localparam [40:1] PF1_AER_CAP_ECRC_CHECK_CAPABLE_REG = PF1_AER_CAP_ECRC_CHECK_CAPABLE;
  localparam [40:1] PF1_AER_CAP_ECRC_GEN_CAPABLE_REG = PF1_AER_CAP_ECRC_GEN_CAPABLE;
  localparam [11:0] PF1_AER_CAP_NEXTPTR_REG = PF1_AER_CAP_NEXTPTR;
  localparam [11:0] PF1_ARI_CAP_NEXTPTR_REG = PF1_ARI_CAP_NEXTPTR;
  localparam [7:0] PF1_ARI_CAP_NEXT_FUNC_REG = PF1_ARI_CAP_NEXT_FUNC;
  localparam [5:0] PF1_BAR0_APERTURE_SIZE_REG = PF1_BAR0_APERTURE_SIZE;
  localparam [2:0] PF1_BAR0_CONTROL_REG = PF1_BAR0_CONTROL;
  localparam [5:0] PF1_BAR1_APERTURE_SIZE_REG = PF1_BAR1_APERTURE_SIZE;
  localparam [2:0] PF1_BAR1_CONTROL_REG = PF1_BAR1_CONTROL;
  localparam [4:0] PF1_BAR2_APERTURE_SIZE_REG = PF1_BAR2_APERTURE_SIZE;
  localparam [2:0] PF1_BAR2_CONTROL_REG = PF1_BAR2_CONTROL;
  localparam [4:0] PF1_BAR3_APERTURE_SIZE_REG = PF1_BAR3_APERTURE_SIZE;
  localparam [2:0] PF1_BAR3_CONTROL_REG = PF1_BAR3_CONTROL;
  localparam [4:0] PF1_BAR4_APERTURE_SIZE_REG = PF1_BAR4_APERTURE_SIZE;
  localparam [2:0] PF1_BAR4_CONTROL_REG = PF1_BAR4_CONTROL;
  localparam [4:0] PF1_BAR5_APERTURE_SIZE_REG = PF1_BAR5_APERTURE_SIZE;
  localparam [2:0] PF1_BAR5_CONTROL_REG = PF1_BAR5_CONTROL;
  localparam [7:0] PF1_BIST_REGISTER_REG = PF1_BIST_REGISTER;
  localparam [7:0] PF1_CAPABILITY_POINTER_REG = PF1_CAPABILITY_POINTER;
  localparam [23:0] PF1_CLASS_CODE_REG = PF1_CLASS_CODE;
  localparam [15:0] PF1_DEVICE_ID_REG = PF1_DEVICE_ID;
  localparam [2:0] PF1_DEV_CAP_MAX_PAYLOAD_SIZE_REG = PF1_DEV_CAP_MAX_PAYLOAD_SIZE;
  localparam [11:0] PF1_DPA_CAP_NEXTPTR_REG = PF1_DPA_CAP_NEXTPTR;
  localparam [4:0] PF1_DPA_CAP_SUB_STATE_CONTROL_REG = PF1_DPA_CAP_SUB_STATE_CONTROL;
  localparam [40:1] PF1_DPA_CAP_SUB_STATE_CONTROL_EN_REG = PF1_DPA_CAP_SUB_STATE_CONTROL_EN;
  localparam [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION0_REG = PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION0;
  localparam [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION1_REG = PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION1;
  localparam [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION2_REG = PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION2;
  localparam [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION3_REG = PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION3;
  localparam [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION4_REG = PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION4;
  localparam [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION5_REG = PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION5;
  localparam [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION6_REG = PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION6;
  localparam [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION7_REG = PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION7;
  localparam [3:0] PF1_DPA_CAP_VER_REG = PF1_DPA_CAP_VER;
  localparam [11:0] PF1_DSN_CAP_NEXTPTR_REG = PF1_DSN_CAP_NEXTPTR;
  localparam [4:0] PF1_EXPANSION_ROM_APERTURE_SIZE_REG = PF1_EXPANSION_ROM_APERTURE_SIZE;
  localparam [40:1] PF1_EXPANSION_ROM_ENABLE_REG = PF1_EXPANSION_ROM_ENABLE;
  localparam [7:0] PF1_INTERRUPT_LINE_REG = PF1_INTERRUPT_LINE;
  localparam [2:0] PF1_INTERRUPT_PIN_REG = PF1_INTERRUPT_PIN;
  localparam [7:0] PF1_MSIX_CAP_NEXTPTR_REG = PF1_MSIX_CAP_NEXTPTR;
  localparam [2:0] PF1_MSIX_CAP_PBA_BIR_REG = PF1_MSIX_CAP_PBA_BIR;
  localparam [28:0] PF1_MSIX_CAP_PBA_OFFSET_REG = PF1_MSIX_CAP_PBA_OFFSET;
  localparam [2:0] PF1_MSIX_CAP_TABLE_BIR_REG = PF1_MSIX_CAP_TABLE_BIR;
  localparam [28:0] PF1_MSIX_CAP_TABLE_OFFSET_REG = PF1_MSIX_CAP_TABLE_OFFSET;
  localparam [10:0] PF1_MSIX_CAP_TABLE_SIZE_REG = PF1_MSIX_CAP_TABLE_SIZE;
  localparam [2:0] PF1_MSI_CAP_MULTIMSGCAP_REG = PF1_MSI_CAP_MULTIMSGCAP;
  localparam [7:0] PF1_MSI_CAP_NEXTPTR_REG = PF1_MSI_CAP_NEXTPTR;
  localparam [40:1] PF1_MSI_CAP_PERVECMASKCAP_REG = PF1_MSI_CAP_PERVECMASKCAP;
  localparam [31:0] PF1_PB_CAP_DATA_REG_D0_REG = PF1_PB_CAP_DATA_REG_D0;
  localparam [31:0] PF1_PB_CAP_DATA_REG_D0_SUSTAINED_REG = PF1_PB_CAP_DATA_REG_D0_SUSTAINED;
  localparam [31:0] PF1_PB_CAP_DATA_REG_D1_REG = PF1_PB_CAP_DATA_REG_D1;
  localparam [31:0] PF1_PB_CAP_DATA_REG_D3HOT_REG = PF1_PB_CAP_DATA_REG_D3HOT;
  localparam [11:0] PF1_PB_CAP_NEXTPTR_REG = PF1_PB_CAP_NEXTPTR;
  localparam [40:1] PF1_PB_CAP_SYSTEM_ALLOCATED_REG = PF1_PB_CAP_SYSTEM_ALLOCATED;
  localparam [3:0] PF1_PB_CAP_VER_REG = PF1_PB_CAP_VER;
  localparam [7:0] PF1_PM_CAP_ID_REG = PF1_PM_CAP_ID;
  localparam [7:0] PF1_PM_CAP_NEXTPTR_REG = PF1_PM_CAP_NEXTPTR;
  localparam [2:0] PF1_PM_CAP_VER_ID_REG = PF1_PM_CAP_VER_ID;
  localparam [40:1] PF1_RBAR_CAP_ENABLE_REG = PF1_RBAR_CAP_ENABLE;
  localparam [11:0] PF1_RBAR_CAP_NEXTPTR_REG = PF1_RBAR_CAP_NEXTPTR;
  localparam [19:0] PF1_RBAR_CAP_SIZE0_REG = PF1_RBAR_CAP_SIZE0;
  localparam [19:0] PF1_RBAR_CAP_SIZE1_REG = PF1_RBAR_CAP_SIZE1;
  localparam [19:0] PF1_RBAR_CAP_SIZE2_REG = PF1_RBAR_CAP_SIZE2;
  localparam [3:0] PF1_RBAR_CAP_VER_REG = PF1_RBAR_CAP_VER;
  localparam [2:0] PF1_RBAR_CONTROL_INDEX0_REG = PF1_RBAR_CONTROL_INDEX0;
  localparam [2:0] PF1_RBAR_CONTROL_INDEX1_REG = PF1_RBAR_CONTROL_INDEX1;
  localparam [2:0] PF1_RBAR_CONTROL_INDEX2_REG = PF1_RBAR_CONTROL_INDEX2;
  localparam [4:0] PF1_RBAR_CONTROL_SIZE0_REG = PF1_RBAR_CONTROL_SIZE0;
  localparam [4:0] PF1_RBAR_CONTROL_SIZE1_REG = PF1_RBAR_CONTROL_SIZE1;
  localparam [4:0] PF1_RBAR_CONTROL_SIZE2_REG = PF1_RBAR_CONTROL_SIZE2;
  localparam [2:0] PF1_RBAR_NUM_REG = PF1_RBAR_NUM;
  localparam [7:0] PF1_REVISION_ID_REG = PF1_REVISION_ID;
  localparam [4:0] PF1_SRIOV_BAR0_APERTURE_SIZE_REG = PF1_SRIOV_BAR0_APERTURE_SIZE;
  localparam [2:0] PF1_SRIOV_BAR0_CONTROL_REG = PF1_SRIOV_BAR0_CONTROL;
  localparam [4:0] PF1_SRIOV_BAR1_APERTURE_SIZE_REG = PF1_SRIOV_BAR1_APERTURE_SIZE;
  localparam [2:0] PF1_SRIOV_BAR1_CONTROL_REG = PF1_SRIOV_BAR1_CONTROL;
  localparam [4:0] PF1_SRIOV_BAR2_APERTURE_SIZE_REG = PF1_SRIOV_BAR2_APERTURE_SIZE;
  localparam [2:0] PF1_SRIOV_BAR2_CONTROL_REG = PF1_SRIOV_BAR2_CONTROL;
  localparam [4:0] PF1_SRIOV_BAR3_APERTURE_SIZE_REG = PF1_SRIOV_BAR3_APERTURE_SIZE;
  localparam [2:0] PF1_SRIOV_BAR3_CONTROL_REG = PF1_SRIOV_BAR3_CONTROL;
  localparam [4:0] PF1_SRIOV_BAR4_APERTURE_SIZE_REG = PF1_SRIOV_BAR4_APERTURE_SIZE;
  localparam [2:0] PF1_SRIOV_BAR4_CONTROL_REG = PF1_SRIOV_BAR4_CONTROL;
  localparam [4:0] PF1_SRIOV_BAR5_APERTURE_SIZE_REG = PF1_SRIOV_BAR5_APERTURE_SIZE;
  localparam [2:0] PF1_SRIOV_BAR5_CONTROL_REG = PF1_SRIOV_BAR5_CONTROL;
  localparam [15:0] PF1_SRIOV_CAP_INITIAL_VF_REG = PF1_SRIOV_CAP_INITIAL_VF;
  localparam [11:0] PF1_SRIOV_CAP_NEXTPTR_REG = PF1_SRIOV_CAP_NEXTPTR;
  localparam [15:0] PF1_SRIOV_CAP_TOTAL_VF_REG = PF1_SRIOV_CAP_TOTAL_VF;
  localparam [3:0] PF1_SRIOV_CAP_VER_REG = PF1_SRIOV_CAP_VER;
  localparam [15:0] PF1_SRIOV_FIRST_VF_OFFSET_REG = PF1_SRIOV_FIRST_VF_OFFSET;
  localparam [15:0] PF1_SRIOV_FUNC_DEP_LINK_REG = PF1_SRIOV_FUNC_DEP_LINK;
  localparam [31:0] PF1_SRIOV_SUPPORTED_PAGE_SIZE_REG = PF1_SRIOV_SUPPORTED_PAGE_SIZE;
  localparam [15:0] PF1_SRIOV_VF_DEVICE_ID_REG = PF1_SRIOV_VF_DEVICE_ID;
  localparam [15:0] PF1_SUBSYSTEM_ID_REG = PF1_SUBSYSTEM_ID;
  localparam [40:1] PF1_TPHR_CAP_DEV_SPECIFIC_MODE_REG = PF1_TPHR_CAP_DEV_SPECIFIC_MODE;
  localparam [40:1] PF1_TPHR_CAP_ENABLE_REG = PF1_TPHR_CAP_ENABLE;
  localparam [40:1] PF1_TPHR_CAP_INT_VEC_MODE_REG = PF1_TPHR_CAP_INT_VEC_MODE;
  localparam [11:0] PF1_TPHR_CAP_NEXTPTR_REG = PF1_TPHR_CAP_NEXTPTR;
  localparam [2:0] PF1_TPHR_CAP_ST_MODE_SEL_REG = PF1_TPHR_CAP_ST_MODE_SEL;
  localparam [1:0] PF1_TPHR_CAP_ST_TABLE_LOC_REG = PF1_TPHR_CAP_ST_TABLE_LOC;
  localparam [10:0] PF1_TPHR_CAP_ST_TABLE_SIZE_REG = PF1_TPHR_CAP_ST_TABLE_SIZE;
  localparam [3:0] PF1_TPHR_CAP_VER_REG = PF1_TPHR_CAP_VER;
  localparam [40:1] PF2_AER_CAP_ECRC_CHECK_CAPABLE_REG = PF2_AER_CAP_ECRC_CHECK_CAPABLE;
  localparam [40:1] PF2_AER_CAP_ECRC_GEN_CAPABLE_REG = PF2_AER_CAP_ECRC_GEN_CAPABLE;
  localparam [11:0] PF2_AER_CAP_NEXTPTR_REG = PF2_AER_CAP_NEXTPTR;
  localparam [11:0] PF2_ARI_CAP_NEXTPTR_REG = PF2_ARI_CAP_NEXTPTR;
  localparam [7:0] PF2_ARI_CAP_NEXT_FUNC_REG = PF2_ARI_CAP_NEXT_FUNC;
  localparam [5:0] PF2_BAR0_APERTURE_SIZE_REG = PF2_BAR0_APERTURE_SIZE;
  localparam [2:0] PF2_BAR0_CONTROL_REG = PF2_BAR0_CONTROL;
  localparam [5:0] PF2_BAR1_APERTURE_SIZE_REG = PF2_BAR1_APERTURE_SIZE;
  localparam [2:0] PF2_BAR1_CONTROL_REG = PF2_BAR1_CONTROL;
  localparam [4:0] PF2_BAR2_APERTURE_SIZE_REG = PF2_BAR2_APERTURE_SIZE;
  localparam [2:0] PF2_BAR2_CONTROL_REG = PF2_BAR2_CONTROL;
  localparam [4:0] PF2_BAR3_APERTURE_SIZE_REG = PF2_BAR3_APERTURE_SIZE;
  localparam [2:0] PF2_BAR3_CONTROL_REG = PF2_BAR3_CONTROL;
  localparam [4:0] PF2_BAR4_APERTURE_SIZE_REG = PF2_BAR4_APERTURE_SIZE;
  localparam [2:0] PF2_BAR4_CONTROL_REG = PF2_BAR4_CONTROL;
  localparam [4:0] PF2_BAR5_APERTURE_SIZE_REG = PF2_BAR5_APERTURE_SIZE;
  localparam [2:0] PF2_BAR5_CONTROL_REG = PF2_BAR5_CONTROL;
  localparam [7:0] PF2_BIST_REGISTER_REG = PF2_BIST_REGISTER;
  localparam [7:0] PF2_CAPABILITY_POINTER_REG = PF2_CAPABILITY_POINTER;
  localparam [23:0] PF2_CLASS_CODE_REG = PF2_CLASS_CODE;
  localparam [15:0] PF2_DEVICE_ID_REG = PF2_DEVICE_ID;
  localparam [2:0] PF2_DEV_CAP_MAX_PAYLOAD_SIZE_REG = PF2_DEV_CAP_MAX_PAYLOAD_SIZE;
  localparam [11:0] PF2_DPA_CAP_NEXTPTR_REG = PF2_DPA_CAP_NEXTPTR;
  localparam [4:0] PF2_DPA_CAP_SUB_STATE_CONTROL_REG = PF2_DPA_CAP_SUB_STATE_CONTROL;
  localparam [40:1] PF2_DPA_CAP_SUB_STATE_CONTROL_EN_REG = PF2_DPA_CAP_SUB_STATE_CONTROL_EN;
  localparam [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION0_REG = PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION0;
  localparam [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION1_REG = PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION1;
  localparam [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION2_REG = PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION2;
  localparam [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION3_REG = PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION3;
  localparam [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION4_REG = PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION4;
  localparam [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION5_REG = PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION5;
  localparam [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION6_REG = PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION6;
  localparam [7:0] PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION7_REG = PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION7;
  localparam [3:0] PF2_DPA_CAP_VER_REG = PF2_DPA_CAP_VER;
  localparam [11:0] PF2_DSN_CAP_NEXTPTR_REG = PF2_DSN_CAP_NEXTPTR;
  localparam [4:0] PF2_EXPANSION_ROM_APERTURE_SIZE_REG = PF2_EXPANSION_ROM_APERTURE_SIZE;
  localparam [40:1] PF2_EXPANSION_ROM_ENABLE_REG = PF2_EXPANSION_ROM_ENABLE;
  localparam [7:0] PF2_INTERRUPT_LINE_REG = PF2_INTERRUPT_LINE;
  localparam [2:0] PF2_INTERRUPT_PIN_REG = PF2_INTERRUPT_PIN;
  localparam [7:0] PF2_MSIX_CAP_NEXTPTR_REG = PF2_MSIX_CAP_NEXTPTR;
  localparam [2:0] PF2_MSIX_CAP_PBA_BIR_REG = PF2_MSIX_CAP_PBA_BIR;
  localparam [28:0] PF2_MSIX_CAP_PBA_OFFSET_REG = PF2_MSIX_CAP_PBA_OFFSET;
  localparam [2:0] PF2_MSIX_CAP_TABLE_BIR_REG = PF2_MSIX_CAP_TABLE_BIR;
  localparam [28:0] PF2_MSIX_CAP_TABLE_OFFSET_REG = PF2_MSIX_CAP_TABLE_OFFSET;
  localparam [10:0] PF2_MSIX_CAP_TABLE_SIZE_REG = PF2_MSIX_CAP_TABLE_SIZE;
  localparam [2:0] PF2_MSI_CAP_MULTIMSGCAP_REG = PF2_MSI_CAP_MULTIMSGCAP;
  localparam [7:0] PF2_MSI_CAP_NEXTPTR_REG = PF2_MSI_CAP_NEXTPTR;
  localparam [40:1] PF2_MSI_CAP_PERVECMASKCAP_REG = PF2_MSI_CAP_PERVECMASKCAP;
  localparam [31:0] PF2_PB_CAP_DATA_REG_D0_REG = PF2_PB_CAP_DATA_REG_D0;
  localparam [31:0] PF2_PB_CAP_DATA_REG_D0_SUSTAINED_REG = PF2_PB_CAP_DATA_REG_D0_SUSTAINED;
  localparam [31:0] PF2_PB_CAP_DATA_REG_D1_REG = PF2_PB_CAP_DATA_REG_D1;
  localparam [31:0] PF2_PB_CAP_DATA_REG_D3HOT_REG = PF2_PB_CAP_DATA_REG_D3HOT;
  localparam [11:0] PF2_PB_CAP_NEXTPTR_REG = PF2_PB_CAP_NEXTPTR;
  localparam [40:1] PF2_PB_CAP_SYSTEM_ALLOCATED_REG = PF2_PB_CAP_SYSTEM_ALLOCATED;
  localparam [3:0] PF2_PB_CAP_VER_REG = PF2_PB_CAP_VER;
  localparam [7:0] PF2_PM_CAP_ID_REG = PF2_PM_CAP_ID;
  localparam [7:0] PF2_PM_CAP_NEXTPTR_REG = PF2_PM_CAP_NEXTPTR;
  localparam [2:0] PF2_PM_CAP_VER_ID_REG = PF2_PM_CAP_VER_ID;
  localparam [40:1] PF2_RBAR_CAP_ENABLE_REG = PF2_RBAR_CAP_ENABLE;
  localparam [11:0] PF2_RBAR_CAP_NEXTPTR_REG = PF2_RBAR_CAP_NEXTPTR;
  localparam [19:0] PF2_RBAR_CAP_SIZE0_REG = PF2_RBAR_CAP_SIZE0;
  localparam [19:0] PF2_RBAR_CAP_SIZE1_REG = PF2_RBAR_CAP_SIZE1;
  localparam [19:0] PF2_RBAR_CAP_SIZE2_REG = PF2_RBAR_CAP_SIZE2;
  localparam [3:0] PF2_RBAR_CAP_VER_REG = PF2_RBAR_CAP_VER;
  localparam [2:0] PF2_RBAR_CONTROL_INDEX0_REG = PF2_RBAR_CONTROL_INDEX0;
  localparam [2:0] PF2_RBAR_CONTROL_INDEX1_REG = PF2_RBAR_CONTROL_INDEX1;
  localparam [2:0] PF2_RBAR_CONTROL_INDEX2_REG = PF2_RBAR_CONTROL_INDEX2;
  localparam [4:0] PF2_RBAR_CONTROL_SIZE0_REG = PF2_RBAR_CONTROL_SIZE0;
  localparam [4:0] PF2_RBAR_CONTROL_SIZE1_REG = PF2_RBAR_CONTROL_SIZE1;
  localparam [4:0] PF2_RBAR_CONTROL_SIZE2_REG = PF2_RBAR_CONTROL_SIZE2;
  localparam [2:0] PF2_RBAR_NUM_REG = PF2_RBAR_NUM;
  localparam [7:0] PF2_REVISION_ID_REG = PF2_REVISION_ID;
  localparam [4:0] PF2_SRIOV_BAR0_APERTURE_SIZE_REG = PF2_SRIOV_BAR0_APERTURE_SIZE;
  localparam [2:0] PF2_SRIOV_BAR0_CONTROL_REG = PF2_SRIOV_BAR0_CONTROL;
  localparam [4:0] PF2_SRIOV_BAR1_APERTURE_SIZE_REG = PF2_SRIOV_BAR1_APERTURE_SIZE;
  localparam [2:0] PF2_SRIOV_BAR1_CONTROL_REG = PF2_SRIOV_BAR1_CONTROL;
  localparam [4:0] PF2_SRIOV_BAR2_APERTURE_SIZE_REG = PF2_SRIOV_BAR2_APERTURE_SIZE;
  localparam [2:0] PF2_SRIOV_BAR2_CONTROL_REG = PF2_SRIOV_BAR2_CONTROL;
  localparam [4:0] PF2_SRIOV_BAR3_APERTURE_SIZE_REG = PF2_SRIOV_BAR3_APERTURE_SIZE;
  localparam [2:0] PF2_SRIOV_BAR3_CONTROL_REG = PF2_SRIOV_BAR3_CONTROL;
  localparam [4:0] PF2_SRIOV_BAR4_APERTURE_SIZE_REG = PF2_SRIOV_BAR4_APERTURE_SIZE;
  localparam [2:0] PF2_SRIOV_BAR4_CONTROL_REG = PF2_SRIOV_BAR4_CONTROL;
  localparam [4:0] PF2_SRIOV_BAR5_APERTURE_SIZE_REG = PF2_SRIOV_BAR5_APERTURE_SIZE;
  localparam [2:0] PF2_SRIOV_BAR5_CONTROL_REG = PF2_SRIOV_BAR5_CONTROL;
  localparam [15:0] PF2_SRIOV_CAP_INITIAL_VF_REG = PF2_SRIOV_CAP_INITIAL_VF;
  localparam [11:0] PF2_SRIOV_CAP_NEXTPTR_REG = PF2_SRIOV_CAP_NEXTPTR;
  localparam [15:0] PF2_SRIOV_CAP_TOTAL_VF_REG = PF2_SRIOV_CAP_TOTAL_VF;
  localparam [3:0] PF2_SRIOV_CAP_VER_REG = PF2_SRIOV_CAP_VER;
  localparam [15:0] PF2_SRIOV_FIRST_VF_OFFSET_REG = PF2_SRIOV_FIRST_VF_OFFSET;
  localparam [15:0] PF2_SRIOV_FUNC_DEP_LINK_REG = PF2_SRIOV_FUNC_DEP_LINK;
  localparam [31:0] PF2_SRIOV_SUPPORTED_PAGE_SIZE_REG = PF2_SRIOV_SUPPORTED_PAGE_SIZE;
  localparam [15:0] PF2_SRIOV_VF_DEVICE_ID_REG = PF2_SRIOV_VF_DEVICE_ID;
  localparam [15:0] PF2_SUBSYSTEM_ID_REG = PF2_SUBSYSTEM_ID;
  localparam [40:1] PF2_TPHR_CAP_DEV_SPECIFIC_MODE_REG = PF2_TPHR_CAP_DEV_SPECIFIC_MODE;
  localparam [40:1] PF2_TPHR_CAP_ENABLE_REG = PF2_TPHR_CAP_ENABLE;
  localparam [40:1] PF2_TPHR_CAP_INT_VEC_MODE_REG = PF2_TPHR_CAP_INT_VEC_MODE;
  localparam [11:0] PF2_TPHR_CAP_NEXTPTR_REG = PF2_TPHR_CAP_NEXTPTR;
  localparam [2:0] PF2_TPHR_CAP_ST_MODE_SEL_REG = PF2_TPHR_CAP_ST_MODE_SEL;
  localparam [1:0] PF2_TPHR_CAP_ST_TABLE_LOC_REG = PF2_TPHR_CAP_ST_TABLE_LOC;
  localparam [10:0] PF2_TPHR_CAP_ST_TABLE_SIZE_REG = PF2_TPHR_CAP_ST_TABLE_SIZE;
  localparam [3:0] PF2_TPHR_CAP_VER_REG = PF2_TPHR_CAP_VER;
  localparam [40:1] PF3_AER_CAP_ECRC_CHECK_CAPABLE_REG = PF3_AER_CAP_ECRC_CHECK_CAPABLE;
  localparam [40:1] PF3_AER_CAP_ECRC_GEN_CAPABLE_REG = PF3_AER_CAP_ECRC_GEN_CAPABLE;
  localparam [11:0] PF3_AER_CAP_NEXTPTR_REG = PF3_AER_CAP_NEXTPTR;
  localparam [11:0] PF3_ARI_CAP_NEXTPTR_REG = PF3_ARI_CAP_NEXTPTR;
  localparam [7:0] PF3_ARI_CAP_NEXT_FUNC_REG = PF3_ARI_CAP_NEXT_FUNC;
  localparam [5:0] PF3_BAR0_APERTURE_SIZE_REG = PF3_BAR0_APERTURE_SIZE;
  localparam [2:0] PF3_BAR0_CONTROL_REG = PF3_BAR0_CONTROL;
  localparam [5:0] PF3_BAR1_APERTURE_SIZE_REG = PF3_BAR1_APERTURE_SIZE;
  localparam [2:0] PF3_BAR1_CONTROL_REG = PF3_BAR1_CONTROL;
  localparam [4:0] PF3_BAR2_APERTURE_SIZE_REG = PF3_BAR2_APERTURE_SIZE;
  localparam [2:0] PF3_BAR2_CONTROL_REG = PF3_BAR2_CONTROL;
  localparam [4:0] PF3_BAR3_APERTURE_SIZE_REG = PF3_BAR3_APERTURE_SIZE;
  localparam [2:0] PF3_BAR3_CONTROL_REG = PF3_BAR3_CONTROL;
  localparam [4:0] PF3_BAR4_APERTURE_SIZE_REG = PF3_BAR4_APERTURE_SIZE;
  localparam [2:0] PF3_BAR4_CONTROL_REG = PF3_BAR4_CONTROL;
  localparam [4:0] PF3_BAR5_APERTURE_SIZE_REG = PF3_BAR5_APERTURE_SIZE;
  localparam [2:0] PF3_BAR5_CONTROL_REG = PF3_BAR5_CONTROL;
  localparam [7:0] PF3_BIST_REGISTER_REG = PF3_BIST_REGISTER;
  localparam [7:0] PF3_CAPABILITY_POINTER_REG = PF3_CAPABILITY_POINTER;
  localparam [23:0] PF3_CLASS_CODE_REG = PF3_CLASS_CODE;
  localparam [15:0] PF3_DEVICE_ID_REG = PF3_DEVICE_ID;
  localparam [2:0] PF3_DEV_CAP_MAX_PAYLOAD_SIZE_REG = PF3_DEV_CAP_MAX_PAYLOAD_SIZE;
  localparam [11:0] PF3_DPA_CAP_NEXTPTR_REG = PF3_DPA_CAP_NEXTPTR;
  localparam [4:0] PF3_DPA_CAP_SUB_STATE_CONTROL_REG = PF3_DPA_CAP_SUB_STATE_CONTROL;
  localparam [40:1] PF3_DPA_CAP_SUB_STATE_CONTROL_EN_REG = PF3_DPA_CAP_SUB_STATE_CONTROL_EN;
  localparam [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION0_REG = PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION0;
  localparam [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION1_REG = PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION1;
  localparam [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION2_REG = PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION2;
  localparam [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION3_REG = PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION3;
  localparam [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION4_REG = PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION4;
  localparam [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION5_REG = PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION5;
  localparam [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION6_REG = PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION6;
  localparam [7:0] PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION7_REG = PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION7;
  localparam [3:0] PF3_DPA_CAP_VER_REG = PF3_DPA_CAP_VER;
  localparam [11:0] PF3_DSN_CAP_NEXTPTR_REG = PF3_DSN_CAP_NEXTPTR;
  localparam [4:0] PF3_EXPANSION_ROM_APERTURE_SIZE_REG = PF3_EXPANSION_ROM_APERTURE_SIZE;
  localparam [40:1] PF3_EXPANSION_ROM_ENABLE_REG = PF3_EXPANSION_ROM_ENABLE;
  localparam [7:0] PF3_INTERRUPT_LINE_REG = PF3_INTERRUPT_LINE;
  localparam [2:0] PF3_INTERRUPT_PIN_REG = PF3_INTERRUPT_PIN;
  localparam [7:0] PF3_MSIX_CAP_NEXTPTR_REG = PF3_MSIX_CAP_NEXTPTR;
  localparam [2:0] PF3_MSIX_CAP_PBA_BIR_REG = PF3_MSIX_CAP_PBA_BIR;
  localparam [28:0] PF3_MSIX_CAP_PBA_OFFSET_REG = PF3_MSIX_CAP_PBA_OFFSET;
  localparam [2:0] PF3_MSIX_CAP_TABLE_BIR_REG = PF3_MSIX_CAP_TABLE_BIR;
  localparam [28:0] PF3_MSIX_CAP_TABLE_OFFSET_REG = PF3_MSIX_CAP_TABLE_OFFSET;
  localparam [10:0] PF3_MSIX_CAP_TABLE_SIZE_REG = PF3_MSIX_CAP_TABLE_SIZE;
  localparam [2:0] PF3_MSI_CAP_MULTIMSGCAP_REG = PF3_MSI_CAP_MULTIMSGCAP;
  localparam [7:0] PF3_MSI_CAP_NEXTPTR_REG = PF3_MSI_CAP_NEXTPTR;
  localparam [40:1] PF3_MSI_CAP_PERVECMASKCAP_REG = PF3_MSI_CAP_PERVECMASKCAP;
  localparam [31:0] PF3_PB_CAP_DATA_REG_D0_REG = PF3_PB_CAP_DATA_REG_D0;
  localparam [31:0] PF3_PB_CAP_DATA_REG_D0_SUSTAINED_REG = PF3_PB_CAP_DATA_REG_D0_SUSTAINED;
  localparam [31:0] PF3_PB_CAP_DATA_REG_D1_REG = PF3_PB_CAP_DATA_REG_D1;
  localparam [31:0] PF3_PB_CAP_DATA_REG_D3HOT_REG = PF3_PB_CAP_DATA_REG_D3HOT;
  localparam [11:0] PF3_PB_CAP_NEXTPTR_REG = PF3_PB_CAP_NEXTPTR;
  localparam [40:1] PF3_PB_CAP_SYSTEM_ALLOCATED_REG = PF3_PB_CAP_SYSTEM_ALLOCATED;
  localparam [3:0] PF3_PB_CAP_VER_REG = PF3_PB_CAP_VER;
  localparam [7:0] PF3_PM_CAP_ID_REG = PF3_PM_CAP_ID;
  localparam [7:0] PF3_PM_CAP_NEXTPTR_REG = PF3_PM_CAP_NEXTPTR;
  localparam [2:0] PF3_PM_CAP_VER_ID_REG = PF3_PM_CAP_VER_ID;
  localparam [40:1] PF3_RBAR_CAP_ENABLE_REG = PF3_RBAR_CAP_ENABLE;
  localparam [11:0] PF3_RBAR_CAP_NEXTPTR_REG = PF3_RBAR_CAP_NEXTPTR;
  localparam [19:0] PF3_RBAR_CAP_SIZE0_REG = PF3_RBAR_CAP_SIZE0;
  localparam [19:0] PF3_RBAR_CAP_SIZE1_REG = PF3_RBAR_CAP_SIZE1;
  localparam [19:0] PF3_RBAR_CAP_SIZE2_REG = PF3_RBAR_CAP_SIZE2;
  localparam [3:0] PF3_RBAR_CAP_VER_REG = PF3_RBAR_CAP_VER;
  localparam [2:0] PF3_RBAR_CONTROL_INDEX0_REG = PF3_RBAR_CONTROL_INDEX0;
  localparam [2:0] PF3_RBAR_CONTROL_INDEX1_REG = PF3_RBAR_CONTROL_INDEX1;
  localparam [2:0] PF3_RBAR_CONTROL_INDEX2_REG = PF3_RBAR_CONTROL_INDEX2;
  localparam [4:0] PF3_RBAR_CONTROL_SIZE0_REG = PF3_RBAR_CONTROL_SIZE0;
  localparam [4:0] PF3_RBAR_CONTROL_SIZE1_REG = PF3_RBAR_CONTROL_SIZE1;
  localparam [4:0] PF3_RBAR_CONTROL_SIZE2_REG = PF3_RBAR_CONTROL_SIZE2;
  localparam [2:0] PF3_RBAR_NUM_REG = PF3_RBAR_NUM;
  localparam [7:0] PF3_REVISION_ID_REG = PF3_REVISION_ID;
  localparam [4:0] PF3_SRIOV_BAR0_APERTURE_SIZE_REG = PF3_SRIOV_BAR0_APERTURE_SIZE;
  localparam [2:0] PF3_SRIOV_BAR0_CONTROL_REG = PF3_SRIOV_BAR0_CONTROL;
  localparam [4:0] PF3_SRIOV_BAR1_APERTURE_SIZE_REG = PF3_SRIOV_BAR1_APERTURE_SIZE;
  localparam [2:0] PF3_SRIOV_BAR1_CONTROL_REG = PF3_SRIOV_BAR1_CONTROL;
  localparam [4:0] PF3_SRIOV_BAR2_APERTURE_SIZE_REG = PF3_SRIOV_BAR2_APERTURE_SIZE;
  localparam [2:0] PF3_SRIOV_BAR2_CONTROL_REG = PF3_SRIOV_BAR2_CONTROL;
  localparam [4:0] PF3_SRIOV_BAR3_APERTURE_SIZE_REG = PF3_SRIOV_BAR3_APERTURE_SIZE;
  localparam [2:0] PF3_SRIOV_BAR3_CONTROL_REG = PF3_SRIOV_BAR3_CONTROL;
  localparam [4:0] PF3_SRIOV_BAR4_APERTURE_SIZE_REG = PF3_SRIOV_BAR4_APERTURE_SIZE;
  localparam [2:0] PF3_SRIOV_BAR4_CONTROL_REG = PF3_SRIOV_BAR4_CONTROL;
  localparam [4:0] PF3_SRIOV_BAR5_APERTURE_SIZE_REG = PF3_SRIOV_BAR5_APERTURE_SIZE;
  localparam [2:0] PF3_SRIOV_BAR5_CONTROL_REG = PF3_SRIOV_BAR5_CONTROL;
  localparam [15:0] PF3_SRIOV_CAP_INITIAL_VF_REG = PF3_SRIOV_CAP_INITIAL_VF;
  localparam [11:0] PF3_SRIOV_CAP_NEXTPTR_REG = PF3_SRIOV_CAP_NEXTPTR;
  localparam [15:0] PF3_SRIOV_CAP_TOTAL_VF_REG = PF3_SRIOV_CAP_TOTAL_VF;
  localparam [3:0] PF3_SRIOV_CAP_VER_REG = PF3_SRIOV_CAP_VER;
  localparam [15:0] PF3_SRIOV_FIRST_VF_OFFSET_REG = PF3_SRIOV_FIRST_VF_OFFSET;
  localparam [15:0] PF3_SRIOV_FUNC_DEP_LINK_REG = PF3_SRIOV_FUNC_DEP_LINK;
  localparam [31:0] PF3_SRIOV_SUPPORTED_PAGE_SIZE_REG = PF3_SRIOV_SUPPORTED_PAGE_SIZE;
  localparam [15:0] PF3_SRIOV_VF_DEVICE_ID_REG = PF3_SRIOV_VF_DEVICE_ID;
  localparam [15:0] PF3_SUBSYSTEM_ID_REG = PF3_SUBSYSTEM_ID;
  localparam [40:1] PF3_TPHR_CAP_DEV_SPECIFIC_MODE_REG = PF3_TPHR_CAP_DEV_SPECIFIC_MODE;
  localparam [40:1] PF3_TPHR_CAP_ENABLE_REG = PF3_TPHR_CAP_ENABLE;
  localparam [40:1] PF3_TPHR_CAP_INT_VEC_MODE_REG = PF3_TPHR_CAP_INT_VEC_MODE;
  localparam [11:0] PF3_TPHR_CAP_NEXTPTR_REG = PF3_TPHR_CAP_NEXTPTR;
  localparam [2:0] PF3_TPHR_CAP_ST_MODE_SEL_REG = PF3_TPHR_CAP_ST_MODE_SEL;
  localparam [1:0] PF3_TPHR_CAP_ST_TABLE_LOC_REG = PF3_TPHR_CAP_ST_TABLE_LOC;
  localparam [10:0] PF3_TPHR_CAP_ST_TABLE_SIZE_REG = PF3_TPHR_CAP_ST_TABLE_SIZE;
  localparam [3:0] PF3_TPHR_CAP_VER_REG = PF3_TPHR_CAP_VER;
  localparam [40:1] PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3_REG = PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3;
  localparam [40:1] PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2_REG = PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2;
  localparam [40:1] PL_DISABLE_EI_INFER_IN_L0_REG = PL_DISABLE_EI_INFER_IN_L0;
  localparam [40:1] PL_DISABLE_GEN3_DC_BALANCE_REG = PL_DISABLE_GEN3_DC_BALANCE;
  localparam [40:1] PL_DISABLE_GEN3_LFSR_UPDATE_ON_SKP_REG = PL_DISABLE_GEN3_LFSR_UPDATE_ON_SKP;
  localparam [40:1] PL_DISABLE_RETRAIN_ON_FRAMING_ERROR_REG = PL_DISABLE_RETRAIN_ON_FRAMING_ERROR;
  localparam [40:1] PL_DISABLE_SCRAMBLING_REG = PL_DISABLE_SCRAMBLING;
  localparam [40:1] PL_DISABLE_SYNC_HEADER_FRAMING_ERROR_REG = PL_DISABLE_SYNC_HEADER_FRAMING_ERROR;
  localparam [40:1] PL_DISABLE_UPCONFIG_CAPABLE_REG = PL_DISABLE_UPCONFIG_CAPABLE;
  localparam [40:1] PL_EQ_ADAPT_DISABLE_COEFF_CHECK_REG = PL_EQ_ADAPT_DISABLE_COEFF_CHECK;
  localparam [40:1] PL_EQ_ADAPT_DISABLE_PRESET_CHECK_REG = PL_EQ_ADAPT_DISABLE_PRESET_CHECK;
  localparam [4:0] PL_EQ_ADAPT_ITER_COUNT_REG = PL_EQ_ADAPT_ITER_COUNT;
  localparam [1:0] PL_EQ_ADAPT_REJECT_RETRY_COUNT_REG = PL_EQ_ADAPT_REJECT_RETRY_COUNT;
  localparam [40:1] PL_EQ_BYPASS_PHASE23_REG = PL_EQ_BYPASS_PHASE23;
  localparam [2:0] PL_EQ_DEFAULT_GEN3_RX_PRESET_HINT_REG = PL_EQ_DEFAULT_GEN3_RX_PRESET_HINT;
  localparam [3:0] PL_EQ_DEFAULT_GEN3_TX_PRESET_REG = PL_EQ_DEFAULT_GEN3_TX_PRESET;
  localparam [40:1] PL_EQ_PHASE01_RX_ADAPT_REG = PL_EQ_PHASE01_RX_ADAPT;
  localparam [40:1] PL_EQ_SHORT_ADAPT_PHASE_REG = PL_EQ_SHORT_ADAPT_PHASE;
  localparam [15:0] PL_LANE0_EQ_CONTROL_REG = PL_LANE0_EQ_CONTROL;
  localparam [15:0] PL_LANE1_EQ_CONTROL_REG = PL_LANE1_EQ_CONTROL;
  localparam [15:0] PL_LANE2_EQ_CONTROL_REG = PL_LANE2_EQ_CONTROL;
  localparam [15:0] PL_LANE3_EQ_CONTROL_REG = PL_LANE3_EQ_CONTROL;
  localparam [15:0] PL_LANE4_EQ_CONTROL_REG = PL_LANE4_EQ_CONTROL;
  localparam [15:0] PL_LANE5_EQ_CONTROL_REG = PL_LANE5_EQ_CONTROL;
  localparam [15:0] PL_LANE6_EQ_CONTROL_REG = PL_LANE6_EQ_CONTROL;
  localparam [15:0] PL_LANE7_EQ_CONTROL_REG = PL_LANE7_EQ_CONTROL;
  localparam [2:0] PL_LINK_CAP_MAX_LINK_SPEED_REG = PL_LINK_CAP_MAX_LINK_SPEED;
  localparam [3:0] PL_LINK_CAP_MAX_LINK_WIDTH_REG = PL_LINK_CAP_MAX_LINK_WIDTH;
  localparam [7:0] PL_N_FTS_COMCLK_GEN1_REG = PL_N_FTS_COMCLK_GEN1;
  localparam [7:0] PL_N_FTS_COMCLK_GEN2_REG = PL_N_FTS_COMCLK_GEN2;
  localparam [7:0] PL_N_FTS_COMCLK_GEN3_REG = PL_N_FTS_COMCLK_GEN3;
  localparam [7:0] PL_N_FTS_GEN1_REG = PL_N_FTS_GEN1;
  localparam [7:0] PL_N_FTS_GEN2_REG = PL_N_FTS_GEN2;
  localparam [7:0] PL_N_FTS_GEN3_REG = PL_N_FTS_GEN3;
  localparam [40:1] PL_REPORT_ALL_PHY_ERRORS_REG = PL_REPORT_ALL_PHY_ERRORS;
  localparam [40:1] PL_SIM_FAST_LINK_TRAINING_REG = PL_SIM_FAST_LINK_TRAINING;
  localparam [40:1] PL_UPSTREAM_FACING_REG = PL_UPSTREAM_FACING;
  localparam [15:0] PM_ASPML0S_TIMEOUT_REG = PM_ASPML0S_TIMEOUT;
  localparam [19:0] PM_ASPML1_ENTRY_DELAY_REG = PM_ASPML1_ENTRY_DELAY;
  localparam [40:1] PM_ENABLE_L23_ENTRY_REG = PM_ENABLE_L23_ENTRY;
  localparam [40:1] PM_ENABLE_SLOT_POWER_CAPTURE_REG = PM_ENABLE_SLOT_POWER_CAPTURE;
  localparam [31:0] PM_L1_REENTRY_DELAY_REG = PM_L1_REENTRY_DELAY;
  localparam [19:0] PM_PME_SERVICE_TIMEOUT_DELAY_REG = PM_PME_SERVICE_TIMEOUT_DELAY;
  localparam [15:0] PM_PME_TURNOFF_ACK_DELAY_REG = PM_PME_TURNOFF_ACK_DELAY;
  localparam [31:0] SIM_JTAG_IDCODE_REG = SIM_JTAG_IDCODE;
  localparam [24:1] SIM_VERSION_REG = SIM_VERSION;
  localparam [0:0] SPARE_BIT0_REG = SPARE_BIT0;
  localparam [0:0] SPARE_BIT1_REG = SPARE_BIT1;
  localparam [0:0] SPARE_BIT2_REG = SPARE_BIT2;
  localparam [0:0] SPARE_BIT3_REG = SPARE_BIT3;
  localparam [0:0] SPARE_BIT4_REG = SPARE_BIT4;
  localparam [0:0] SPARE_BIT5_REG = SPARE_BIT5;
  localparam [0:0] SPARE_BIT6_REG = SPARE_BIT6;
  localparam [0:0] SPARE_BIT7_REG = SPARE_BIT7;
  localparam [0:0] SPARE_BIT8_REG = SPARE_BIT8;
  localparam [7:0] SPARE_BYTE0_REG = SPARE_BYTE0;
  localparam [7:0] SPARE_BYTE1_REG = SPARE_BYTE1;
  localparam [7:0] SPARE_BYTE2_REG = SPARE_BYTE2;
  localparam [7:0] SPARE_BYTE3_REG = SPARE_BYTE3;
  localparam [31:0] SPARE_WORD0_REG = SPARE_WORD0;
  localparam [31:0] SPARE_WORD1_REG = SPARE_WORD1;
  localparam [31:0] SPARE_WORD2_REG = SPARE_WORD2;
  localparam [31:0] SPARE_WORD3_REG = SPARE_WORD3;
  localparam [40:1] SRIOV_CAP_ENABLE_REG = SRIOV_CAP_ENABLE;
  localparam [40:1] TL_COMPLETION_RAM_SIZE_16K_REG = TL_COMPLETION_RAM_SIZE_16K;
  localparam [23:0] TL_COMPL_TIMEOUT_REG0_REG = TL_COMPL_TIMEOUT_REG0;
  localparam [27:0] TL_COMPL_TIMEOUT_REG1_REG = TL_COMPL_TIMEOUT_REG1;
  localparam [11:0] TL_CREDITS_CD_REG = TL_CREDITS_CD;
  localparam [7:0] TL_CREDITS_CH_REG = TL_CREDITS_CH;
  localparam [11:0] TL_CREDITS_NPD_REG = TL_CREDITS_NPD;
  localparam [7:0] TL_CREDITS_NPH_REG = TL_CREDITS_NPH;
  localparam [11:0] TL_CREDITS_PD_REG = TL_CREDITS_PD;
  localparam [7:0] TL_CREDITS_PH_REG = TL_CREDITS_PH;
  localparam [40:1] TL_ENABLE_MESSAGE_RID_CHECK_ENABLE_REG = TL_ENABLE_MESSAGE_RID_CHECK_ENABLE;
  localparam [40:1] TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE_REG = TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE;
  localparam [40:1] TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE_REG = TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE;
  localparam [40:1] TL_LEGACY_MODE_ENABLE_REG = TL_LEGACY_MODE_ENABLE;
  localparam [1:0] TL_PF_ENABLE_REG_REG = TL_PF_ENABLE_REG;
  localparam [40:1] TL_TX_MUX_STRICT_PRIORITY_REG = TL_TX_MUX_STRICT_PRIORITY;
  localparam [40:1] TWO_LAYER_MODE_DLCMSM_ENABLE_REG = TWO_LAYER_MODE_DLCMSM_ENABLE;
  localparam [40:1] TWO_LAYER_MODE_ENABLE_REG = TWO_LAYER_MODE_ENABLE;
  localparam [40:1] TWO_LAYER_MODE_WIDTH_256_REG = TWO_LAYER_MODE_WIDTH_256;
  localparam [11:0] VF0_ARI_CAP_NEXTPTR_REG = VF0_ARI_CAP_NEXTPTR;
  localparam [7:0] VF0_CAPABILITY_POINTER_REG = VF0_CAPABILITY_POINTER;
  localparam [2:0] VF0_MSIX_CAP_PBA_BIR_REG = VF0_MSIX_CAP_PBA_BIR;
  localparam [28:0] VF0_MSIX_CAP_PBA_OFFSET_REG = VF0_MSIX_CAP_PBA_OFFSET;
  localparam [2:0] VF0_MSIX_CAP_TABLE_BIR_REG = VF0_MSIX_CAP_TABLE_BIR;
  localparam [28:0] VF0_MSIX_CAP_TABLE_OFFSET_REG = VF0_MSIX_CAP_TABLE_OFFSET;
  localparam [10:0] VF0_MSIX_CAP_TABLE_SIZE_REG = VF0_MSIX_CAP_TABLE_SIZE;
  localparam [2:0] VF0_MSI_CAP_MULTIMSGCAP_REG = VF0_MSI_CAP_MULTIMSGCAP;
  localparam [7:0] VF0_PM_CAP_ID_REG = VF0_PM_CAP_ID;
  localparam [7:0] VF0_PM_CAP_NEXTPTR_REG = VF0_PM_CAP_NEXTPTR;
  localparam [2:0] VF0_PM_CAP_VER_ID_REG = VF0_PM_CAP_VER_ID;
  localparam [40:1] VF0_TPHR_CAP_DEV_SPECIFIC_MODE_REG = VF0_TPHR_CAP_DEV_SPECIFIC_MODE;
  localparam [40:1] VF0_TPHR_CAP_ENABLE_REG = VF0_TPHR_CAP_ENABLE;
  localparam [40:1] VF0_TPHR_CAP_INT_VEC_MODE_REG = VF0_TPHR_CAP_INT_VEC_MODE;
  localparam [11:0] VF0_TPHR_CAP_NEXTPTR_REG = VF0_TPHR_CAP_NEXTPTR;
  localparam [2:0] VF0_TPHR_CAP_ST_MODE_SEL_REG = VF0_TPHR_CAP_ST_MODE_SEL;
  localparam [1:0] VF0_TPHR_CAP_ST_TABLE_LOC_REG = VF0_TPHR_CAP_ST_TABLE_LOC;
  localparam [10:0] VF0_TPHR_CAP_ST_TABLE_SIZE_REG = VF0_TPHR_CAP_ST_TABLE_SIZE;
  localparam [3:0] VF0_TPHR_CAP_VER_REG = VF0_TPHR_CAP_VER;
  localparam [11:0] VF1_ARI_CAP_NEXTPTR_REG = VF1_ARI_CAP_NEXTPTR;
  localparam [2:0] VF1_MSIX_CAP_PBA_BIR_REG = VF1_MSIX_CAP_PBA_BIR;
  localparam [28:0] VF1_MSIX_CAP_PBA_OFFSET_REG = VF1_MSIX_CAP_PBA_OFFSET;
  localparam [2:0] VF1_MSIX_CAP_TABLE_BIR_REG = VF1_MSIX_CAP_TABLE_BIR;
  localparam [28:0] VF1_MSIX_CAP_TABLE_OFFSET_REG = VF1_MSIX_CAP_TABLE_OFFSET;
  localparam [10:0] VF1_MSIX_CAP_TABLE_SIZE_REG = VF1_MSIX_CAP_TABLE_SIZE;
  localparam [2:0] VF1_MSI_CAP_MULTIMSGCAP_REG = VF1_MSI_CAP_MULTIMSGCAP;
  localparam [7:0] VF1_PM_CAP_ID_REG = VF1_PM_CAP_ID;
  localparam [7:0] VF1_PM_CAP_NEXTPTR_REG = VF1_PM_CAP_NEXTPTR;
  localparam [2:0] VF1_PM_CAP_VER_ID_REG = VF1_PM_CAP_VER_ID;
  localparam [40:1] VF1_TPHR_CAP_DEV_SPECIFIC_MODE_REG = VF1_TPHR_CAP_DEV_SPECIFIC_MODE;
  localparam [40:1] VF1_TPHR_CAP_ENABLE_REG = VF1_TPHR_CAP_ENABLE;
  localparam [40:1] VF1_TPHR_CAP_INT_VEC_MODE_REG = VF1_TPHR_CAP_INT_VEC_MODE;
  localparam [11:0] VF1_TPHR_CAP_NEXTPTR_REG = VF1_TPHR_CAP_NEXTPTR;
  localparam [2:0] VF1_TPHR_CAP_ST_MODE_SEL_REG = VF1_TPHR_CAP_ST_MODE_SEL;
  localparam [1:0] VF1_TPHR_CAP_ST_TABLE_LOC_REG = VF1_TPHR_CAP_ST_TABLE_LOC;
  localparam [10:0] VF1_TPHR_CAP_ST_TABLE_SIZE_REG = VF1_TPHR_CAP_ST_TABLE_SIZE;
  localparam [3:0] VF1_TPHR_CAP_VER_REG = VF1_TPHR_CAP_VER;
  localparam [11:0] VF2_ARI_CAP_NEXTPTR_REG = VF2_ARI_CAP_NEXTPTR;
  localparam [2:0] VF2_MSIX_CAP_PBA_BIR_REG = VF2_MSIX_CAP_PBA_BIR;
  localparam [28:0] VF2_MSIX_CAP_PBA_OFFSET_REG = VF2_MSIX_CAP_PBA_OFFSET;
  localparam [2:0] VF2_MSIX_CAP_TABLE_BIR_REG = VF2_MSIX_CAP_TABLE_BIR;
  localparam [28:0] VF2_MSIX_CAP_TABLE_OFFSET_REG = VF2_MSIX_CAP_TABLE_OFFSET;
  localparam [10:0] VF2_MSIX_CAP_TABLE_SIZE_REG = VF2_MSIX_CAP_TABLE_SIZE;
  localparam [2:0] VF2_MSI_CAP_MULTIMSGCAP_REG = VF2_MSI_CAP_MULTIMSGCAP;
  localparam [7:0] VF2_PM_CAP_ID_REG = VF2_PM_CAP_ID;
  localparam [7:0] VF2_PM_CAP_NEXTPTR_REG = VF2_PM_CAP_NEXTPTR;
  localparam [2:0] VF2_PM_CAP_VER_ID_REG = VF2_PM_CAP_VER_ID;
  localparam [40:1] VF2_TPHR_CAP_DEV_SPECIFIC_MODE_REG = VF2_TPHR_CAP_DEV_SPECIFIC_MODE;
  localparam [40:1] VF2_TPHR_CAP_ENABLE_REG = VF2_TPHR_CAP_ENABLE;
  localparam [40:1] VF2_TPHR_CAP_INT_VEC_MODE_REG = VF2_TPHR_CAP_INT_VEC_MODE;
  localparam [11:0] VF2_TPHR_CAP_NEXTPTR_REG = VF2_TPHR_CAP_NEXTPTR;
  localparam [2:0] VF2_TPHR_CAP_ST_MODE_SEL_REG = VF2_TPHR_CAP_ST_MODE_SEL;
  localparam [1:0] VF2_TPHR_CAP_ST_TABLE_LOC_REG = VF2_TPHR_CAP_ST_TABLE_LOC;
  localparam [10:0] VF2_TPHR_CAP_ST_TABLE_SIZE_REG = VF2_TPHR_CAP_ST_TABLE_SIZE;
  localparam [3:0] VF2_TPHR_CAP_VER_REG = VF2_TPHR_CAP_VER;
  localparam [11:0] VF3_ARI_CAP_NEXTPTR_REG = VF3_ARI_CAP_NEXTPTR;
  localparam [2:0] VF3_MSIX_CAP_PBA_BIR_REG = VF3_MSIX_CAP_PBA_BIR;
  localparam [28:0] VF3_MSIX_CAP_PBA_OFFSET_REG = VF3_MSIX_CAP_PBA_OFFSET;
  localparam [2:0] VF3_MSIX_CAP_TABLE_BIR_REG = VF3_MSIX_CAP_TABLE_BIR;
  localparam [28:0] VF3_MSIX_CAP_TABLE_OFFSET_REG = VF3_MSIX_CAP_TABLE_OFFSET;
  localparam [10:0] VF3_MSIX_CAP_TABLE_SIZE_REG = VF3_MSIX_CAP_TABLE_SIZE;
  localparam [2:0] VF3_MSI_CAP_MULTIMSGCAP_REG = VF3_MSI_CAP_MULTIMSGCAP;
  localparam [7:0] VF3_PM_CAP_ID_REG = VF3_PM_CAP_ID;
  localparam [7:0] VF3_PM_CAP_NEXTPTR_REG = VF3_PM_CAP_NEXTPTR;
  localparam [2:0] VF3_PM_CAP_VER_ID_REG = VF3_PM_CAP_VER_ID;
  localparam [40:1] VF3_TPHR_CAP_DEV_SPECIFIC_MODE_REG = VF3_TPHR_CAP_DEV_SPECIFIC_MODE;
  localparam [40:1] VF3_TPHR_CAP_ENABLE_REG = VF3_TPHR_CAP_ENABLE;
  localparam [40:1] VF3_TPHR_CAP_INT_VEC_MODE_REG = VF3_TPHR_CAP_INT_VEC_MODE;
  localparam [11:0] VF3_TPHR_CAP_NEXTPTR_REG = VF3_TPHR_CAP_NEXTPTR;
  localparam [2:0] VF3_TPHR_CAP_ST_MODE_SEL_REG = VF3_TPHR_CAP_ST_MODE_SEL;
  localparam [1:0] VF3_TPHR_CAP_ST_TABLE_LOC_REG = VF3_TPHR_CAP_ST_TABLE_LOC;
  localparam [10:0] VF3_TPHR_CAP_ST_TABLE_SIZE_REG = VF3_TPHR_CAP_ST_TABLE_SIZE;
  localparam [3:0] VF3_TPHR_CAP_VER_REG = VF3_TPHR_CAP_VER;
  localparam [11:0] VF4_ARI_CAP_NEXTPTR_REG = VF4_ARI_CAP_NEXTPTR;
  localparam [2:0] VF4_MSIX_CAP_PBA_BIR_REG = VF4_MSIX_CAP_PBA_BIR;
  localparam [28:0] VF4_MSIX_CAP_PBA_OFFSET_REG = VF4_MSIX_CAP_PBA_OFFSET;
  localparam [2:0] VF4_MSIX_CAP_TABLE_BIR_REG = VF4_MSIX_CAP_TABLE_BIR;
  localparam [28:0] VF4_MSIX_CAP_TABLE_OFFSET_REG = VF4_MSIX_CAP_TABLE_OFFSET;
  localparam [10:0] VF4_MSIX_CAP_TABLE_SIZE_REG = VF4_MSIX_CAP_TABLE_SIZE;
  localparam [2:0] VF4_MSI_CAP_MULTIMSGCAP_REG = VF4_MSI_CAP_MULTIMSGCAP;
  localparam [7:0] VF4_PM_CAP_ID_REG = VF4_PM_CAP_ID;
  localparam [7:0] VF4_PM_CAP_NEXTPTR_REG = VF4_PM_CAP_NEXTPTR;
  localparam [2:0] VF4_PM_CAP_VER_ID_REG = VF4_PM_CAP_VER_ID;
  localparam [40:1] VF4_TPHR_CAP_DEV_SPECIFIC_MODE_REG = VF4_TPHR_CAP_DEV_SPECIFIC_MODE;
  localparam [40:1] VF4_TPHR_CAP_ENABLE_REG = VF4_TPHR_CAP_ENABLE;
  localparam [40:1] VF4_TPHR_CAP_INT_VEC_MODE_REG = VF4_TPHR_CAP_INT_VEC_MODE;
  localparam [11:0] VF4_TPHR_CAP_NEXTPTR_REG = VF4_TPHR_CAP_NEXTPTR;
  localparam [2:0] VF4_TPHR_CAP_ST_MODE_SEL_REG = VF4_TPHR_CAP_ST_MODE_SEL;
  localparam [1:0] VF4_TPHR_CAP_ST_TABLE_LOC_REG = VF4_TPHR_CAP_ST_TABLE_LOC;
  localparam [10:0] VF4_TPHR_CAP_ST_TABLE_SIZE_REG = VF4_TPHR_CAP_ST_TABLE_SIZE;
  localparam [3:0] VF4_TPHR_CAP_VER_REG = VF4_TPHR_CAP_VER;
  localparam [11:0] VF5_ARI_CAP_NEXTPTR_REG = VF5_ARI_CAP_NEXTPTR;
  localparam [2:0] VF5_MSIX_CAP_PBA_BIR_REG = VF5_MSIX_CAP_PBA_BIR;
  localparam [28:0] VF5_MSIX_CAP_PBA_OFFSET_REG = VF5_MSIX_CAP_PBA_OFFSET;
  localparam [2:0] VF5_MSIX_CAP_TABLE_BIR_REG = VF5_MSIX_CAP_TABLE_BIR;
  localparam [28:0] VF5_MSIX_CAP_TABLE_OFFSET_REG = VF5_MSIX_CAP_TABLE_OFFSET;
  localparam [10:0] VF5_MSIX_CAP_TABLE_SIZE_REG = VF5_MSIX_CAP_TABLE_SIZE;
  localparam [2:0] VF5_MSI_CAP_MULTIMSGCAP_REG = VF5_MSI_CAP_MULTIMSGCAP;
  localparam [7:0] VF5_PM_CAP_ID_REG = VF5_PM_CAP_ID;
  localparam [7:0] VF5_PM_CAP_NEXTPTR_REG = VF5_PM_CAP_NEXTPTR;
  localparam [2:0] VF5_PM_CAP_VER_ID_REG = VF5_PM_CAP_VER_ID;
  localparam [40:1] VF5_TPHR_CAP_DEV_SPECIFIC_MODE_REG = VF5_TPHR_CAP_DEV_SPECIFIC_MODE;
  localparam [40:1] VF5_TPHR_CAP_ENABLE_REG = VF5_TPHR_CAP_ENABLE;
  localparam [40:1] VF5_TPHR_CAP_INT_VEC_MODE_REG = VF5_TPHR_CAP_INT_VEC_MODE;
  localparam [11:0] VF5_TPHR_CAP_NEXTPTR_REG = VF5_TPHR_CAP_NEXTPTR;
  localparam [2:0] VF5_TPHR_CAP_ST_MODE_SEL_REG = VF5_TPHR_CAP_ST_MODE_SEL;
  localparam [1:0] VF5_TPHR_CAP_ST_TABLE_LOC_REG = VF5_TPHR_CAP_ST_TABLE_LOC;
  localparam [10:0] VF5_TPHR_CAP_ST_TABLE_SIZE_REG = VF5_TPHR_CAP_ST_TABLE_SIZE;
  localparam [3:0] VF5_TPHR_CAP_VER_REG = VF5_TPHR_CAP_VER;
  localparam [11:0] VF6_ARI_CAP_NEXTPTR_REG = VF6_ARI_CAP_NEXTPTR;
  localparam [2:0] VF6_MSIX_CAP_PBA_BIR_REG = VF6_MSIX_CAP_PBA_BIR;
  localparam [28:0] VF6_MSIX_CAP_PBA_OFFSET_REG = VF6_MSIX_CAP_PBA_OFFSET;
  localparam [2:0] VF6_MSIX_CAP_TABLE_BIR_REG = VF6_MSIX_CAP_TABLE_BIR;
  localparam [28:0] VF6_MSIX_CAP_TABLE_OFFSET_REG = VF6_MSIX_CAP_TABLE_OFFSET;
  localparam [10:0] VF6_MSIX_CAP_TABLE_SIZE_REG = VF6_MSIX_CAP_TABLE_SIZE;
  localparam [2:0] VF6_MSI_CAP_MULTIMSGCAP_REG = VF6_MSI_CAP_MULTIMSGCAP;
  localparam [7:0] VF6_PM_CAP_ID_REG = VF6_PM_CAP_ID;
  localparam [7:0] VF6_PM_CAP_NEXTPTR_REG = VF6_PM_CAP_NEXTPTR;
  localparam [2:0] VF6_PM_CAP_VER_ID_REG = VF6_PM_CAP_VER_ID;
  localparam [40:1] VF6_TPHR_CAP_DEV_SPECIFIC_MODE_REG = VF6_TPHR_CAP_DEV_SPECIFIC_MODE;
  localparam [40:1] VF6_TPHR_CAP_ENABLE_REG = VF6_TPHR_CAP_ENABLE;
  localparam [40:1] VF6_TPHR_CAP_INT_VEC_MODE_REG = VF6_TPHR_CAP_INT_VEC_MODE;
  localparam [11:0] VF6_TPHR_CAP_NEXTPTR_REG = VF6_TPHR_CAP_NEXTPTR;
  localparam [2:0] VF6_TPHR_CAP_ST_MODE_SEL_REG = VF6_TPHR_CAP_ST_MODE_SEL;
  localparam [1:0] VF6_TPHR_CAP_ST_TABLE_LOC_REG = VF6_TPHR_CAP_ST_TABLE_LOC;
  localparam [10:0] VF6_TPHR_CAP_ST_TABLE_SIZE_REG = VF6_TPHR_CAP_ST_TABLE_SIZE;
  localparam [3:0] VF6_TPHR_CAP_VER_REG = VF6_TPHR_CAP_VER;
  localparam [11:0] VF7_ARI_CAP_NEXTPTR_REG = VF7_ARI_CAP_NEXTPTR;
  localparam [2:0] VF7_MSIX_CAP_PBA_BIR_REG = VF7_MSIX_CAP_PBA_BIR;
  localparam [28:0] VF7_MSIX_CAP_PBA_OFFSET_REG = VF7_MSIX_CAP_PBA_OFFSET;
  localparam [2:0] VF7_MSIX_CAP_TABLE_BIR_REG = VF7_MSIX_CAP_TABLE_BIR;
  localparam [28:0] VF7_MSIX_CAP_TABLE_OFFSET_REG = VF7_MSIX_CAP_TABLE_OFFSET;
  localparam [10:0] VF7_MSIX_CAP_TABLE_SIZE_REG = VF7_MSIX_CAP_TABLE_SIZE;
  localparam [2:0] VF7_MSI_CAP_MULTIMSGCAP_REG = VF7_MSI_CAP_MULTIMSGCAP;
  localparam [7:0] VF7_PM_CAP_ID_REG = VF7_PM_CAP_ID;
  localparam [7:0] VF7_PM_CAP_NEXTPTR_REG = VF7_PM_CAP_NEXTPTR;
  localparam [2:0] VF7_PM_CAP_VER_ID_REG = VF7_PM_CAP_VER_ID;
  localparam [40:1] VF7_TPHR_CAP_DEV_SPECIFIC_MODE_REG = VF7_TPHR_CAP_DEV_SPECIFIC_MODE;
  localparam [40:1] VF7_TPHR_CAP_ENABLE_REG = VF7_TPHR_CAP_ENABLE;
  localparam [40:1] VF7_TPHR_CAP_INT_VEC_MODE_REG = VF7_TPHR_CAP_INT_VEC_MODE;
  localparam [11:0] VF7_TPHR_CAP_NEXTPTR_REG = VF7_TPHR_CAP_NEXTPTR;
  localparam [2:0] VF7_TPHR_CAP_ST_MODE_SEL_REG = VF7_TPHR_CAP_ST_MODE_SEL;
  localparam [1:0] VF7_TPHR_CAP_ST_TABLE_LOC_REG = VF7_TPHR_CAP_ST_TABLE_LOC;
  localparam [10:0] VF7_TPHR_CAP_ST_TABLE_SIZE_REG = VF7_TPHR_CAP_ST_TABLE_SIZE;
  localparam [3:0] VF7_TPHR_CAP_VER_REG = VF7_TPHR_CAP_VER;
  `endif

  localparam [40:1] TEST_MODE_PIN_CHAR_REG = "FALSE";

  tri0 glblGSR = glbl.GSR;

  `ifdef XIL_TIMING //Simprim 
  reg notifier;
  `endif
  reg trig_attr = 1'b0;
  reg attr_err = 1'b0;
  
// include dynamic registers - XILINX test only
  `ifdef XIL_DR
  `include "PCIE_3_1_dr.v"
  `endif

  wire CFGERRCOROUT_out;
  wire CFGERRFATALOUT_out;
  wire CFGERRNONFATALOUT_out;
  wire CFGEXTREADRECEIVED_out;
  wire CFGEXTWRITERECEIVED_out;
  wire CFGHOTRESETOUT_out;
  wire CFGINTERRUPTMSIFAIL_out;
  wire CFGINTERRUPTMSIMASKUPDATE_out;
  wire CFGINTERRUPTMSISENT_out;
  wire CFGINTERRUPTMSIXFAIL_out;
  wire CFGINTERRUPTMSIXSENT_out;
  wire CFGINTERRUPTSENT_out;
  wire CFGLOCALERROR_out;
  wire CFGLTRENABLE_out;
  wire CFGMGMTREADWRITEDONE_out;
  wire CFGMSGRECEIVED_out;
  wire CFGMSGTRANSMITDONE_out;
  wire CFGPERFUNCTIONUPDATEDONE_out;
  wire CFGPHYLINKDOWN_out;
  wire CFGPLSTATUSCHANGE_out;
  wire CFGPOWERSTATECHANGEINTERRUPT_out;
  wire CFGTPHSTTREADENABLE_out;
  wire CFGTPHSTTWRITEENABLE_out;
  wire CONFMCAPDESIGNSWITCH_out;
  wire CONFMCAPEOS_out;
  wire CONFMCAPINUSEBYPCIE_out;
  wire CONFREQREADY_out;
  wire CONFRESPVALID_out;
  wire DBGMCAPCSB_out;
  wire DBGMCAPEOS_out;
  wire DBGMCAPERROR_out;
  wire DBGMCAPMODE_out;
  wire DBGMCAPRDATAVALID_out;
  wire DBGMCAPRDWRB_out;
  wire DBGMCAPRESET_out;
  wire DBGPLDATABLOCKRECEIVEDAFTEREDS_out;
  wire DBGPLGEN3FRAMINGERRORDETECTED_out;
  wire DBGPLGEN3SYNCHEADERERRORDETECTED_out;
  wire DRPRDY_out;
  wire LL2LMMASTERTLPSENT0_out;
  wire LL2LMMASTERTLPSENT1_out;
  wire MAXISCQTLAST_out;
  wire MAXISCQTVALID_out;
  wire MAXISRCTLAST_out;
  wire MAXISRCTVALID_out;
  wire PCIEPERST0B_out;
  wire PCIEPERST1B_out;
  wire PCIERQSEQNUMVLD_out;
  wire PCIERQTAGVLD_out;
  wire PIPERX0POLARITY_out;
  wire PIPERX1POLARITY_out;
  wire PIPERX2POLARITY_out;
  wire PIPERX3POLARITY_out;
  wire PIPERX4POLARITY_out;
  wire PIPERX5POLARITY_out;
  wire PIPERX6POLARITY_out;
  wire PIPERX7POLARITY_out;
  wire PIPETX0COMPLIANCE_out;
  wire PIPETX0DATAVALID_out;
  wire PIPETX0DEEMPH_out;
  wire PIPETX0ELECIDLE_out;
  wire PIPETX0RCVRDET_out;
  wire PIPETX0RESET_out;
  wire PIPETX0STARTBLOCK_out;
  wire PIPETX0SWING_out;
  wire PIPETX1COMPLIANCE_out;
  wire PIPETX1DATAVALID_out;
  wire PIPETX1DEEMPH_out;
  wire PIPETX1ELECIDLE_out;
  wire PIPETX1RCVRDET_out;
  wire PIPETX1RESET_out;
  wire PIPETX1STARTBLOCK_out;
  wire PIPETX1SWING_out;
  wire PIPETX2COMPLIANCE_out;
  wire PIPETX2DATAVALID_out;
  wire PIPETX2DEEMPH_out;
  wire PIPETX2ELECIDLE_out;
  wire PIPETX2RCVRDET_out;
  wire PIPETX2RESET_out;
  wire PIPETX2STARTBLOCK_out;
  wire PIPETX2SWING_out;
  wire PIPETX3COMPLIANCE_out;
  wire PIPETX3DATAVALID_out;
  wire PIPETX3DEEMPH_out;
  wire PIPETX3ELECIDLE_out;
  wire PIPETX3RCVRDET_out;
  wire PIPETX3RESET_out;
  wire PIPETX3STARTBLOCK_out;
  wire PIPETX3SWING_out;
  wire PIPETX4COMPLIANCE_out;
  wire PIPETX4DATAVALID_out;
  wire PIPETX4DEEMPH_out;
  wire PIPETX4ELECIDLE_out;
  wire PIPETX4RCVRDET_out;
  wire PIPETX4RESET_out;
  wire PIPETX4STARTBLOCK_out;
  wire PIPETX4SWING_out;
  wire PIPETX5COMPLIANCE_out;
  wire PIPETX5DATAVALID_out;
  wire PIPETX5DEEMPH_out;
  wire PIPETX5ELECIDLE_out;
  wire PIPETX5RCVRDET_out;
  wire PIPETX5RESET_out;
  wire PIPETX5STARTBLOCK_out;
  wire PIPETX5SWING_out;
  wire PIPETX6COMPLIANCE_out;
  wire PIPETX6DATAVALID_out;
  wire PIPETX6DEEMPH_out;
  wire PIPETX6ELECIDLE_out;
  wire PIPETX6RCVRDET_out;
  wire PIPETX6RESET_out;
  wire PIPETX6STARTBLOCK_out;
  wire PIPETX6SWING_out;
  wire PIPETX7COMPLIANCE_out;
  wire PIPETX7DATAVALID_out;
  wire PIPETX7DEEMPH_out;
  wire PIPETX7ELECIDLE_out;
  wire PIPETX7RCVRDET_out;
  wire PIPETX7RESET_out;
  wire PIPETX7STARTBLOCK_out;
  wire PIPETX7SWING_out;
  wire PLEQINPROGRESS_out;
  wire PMVOUT_out;
  wire [11:0] CFGFCCPLD_out;
  wire [11:0] CFGFCNPD_out;
  wire [11:0] CFGFCPD_out;
  wire [11:0] CFGFUNCTIONPOWERSTATE_out;
  wire [11:0] CFGINTERRUPTMSIMMENABLE_out;
  wire [11:0] CFGTPHSTMODE_out;
  wire [143:0] MIREPLAYRAMWRITEDATA_out;
  wire [143:0] MIREQUESTRAMWRITEDATA_out;
  wire [15:0] CFGFUNCTIONSTATUS_out;
  wire [15:0] CFGPERFUNCSTATUSDATA_out;
  wire [15:0] CFGVFSTATUS_out;
  wire [15:0] DBGDATAOUT_out;
  wire [15:0] DRPDO_out;
  wire [17:0] LL2LMMAXISRXTUSER_out;
  wire [1:0] CFGLINKPOWERSTATE_out;
  wire [1:0] CFGOBFFENABLE_out;
  wire [1:0] CFGPHYLINKSTATUS_out;
  wire [1:0] MIREPLAYRAMREADENABLE_out;
  wire [1:0] MIREPLAYRAMWRITEENABLE_out;
  wire [1:0] PCIERQTAGAV_out;
  wire [1:0] PCIETFCNPDAV_out;
  wire [1:0] PCIETFCNPHAV_out;
  wire [1:0] PIPERX0EQCONTROL_out;
  wire [1:0] PIPERX1EQCONTROL_out;
  wire [1:0] PIPERX2EQCONTROL_out;
  wire [1:0] PIPERX3EQCONTROL_out;
  wire [1:0] PIPERX4EQCONTROL_out;
  wire [1:0] PIPERX5EQCONTROL_out;
  wire [1:0] PIPERX6EQCONTROL_out;
  wire [1:0] PIPERX7EQCONTROL_out;
  wire [1:0] PIPETX0CHARISK_out;
  wire [1:0] PIPETX0EQCONTROL_out;
  wire [1:0] PIPETX0POWERDOWN_out;
  wire [1:0] PIPETX0RATE_out;
  wire [1:0] PIPETX0SYNCHEADER_out;
  wire [1:0] PIPETX1CHARISK_out;
  wire [1:0] PIPETX1EQCONTROL_out;
  wire [1:0] PIPETX1POWERDOWN_out;
  wire [1:0] PIPETX1RATE_out;
  wire [1:0] PIPETX1SYNCHEADER_out;
  wire [1:0] PIPETX2CHARISK_out;
  wire [1:0] PIPETX2EQCONTROL_out;
  wire [1:0] PIPETX2POWERDOWN_out;
  wire [1:0] PIPETX2RATE_out;
  wire [1:0] PIPETX2SYNCHEADER_out;
  wire [1:0] PIPETX3CHARISK_out;
  wire [1:0] PIPETX3EQCONTROL_out;
  wire [1:0] PIPETX3POWERDOWN_out;
  wire [1:0] PIPETX3RATE_out;
  wire [1:0] PIPETX3SYNCHEADER_out;
  wire [1:0] PIPETX4CHARISK_out;
  wire [1:0] PIPETX4EQCONTROL_out;
  wire [1:0] PIPETX4POWERDOWN_out;
  wire [1:0] PIPETX4RATE_out;
  wire [1:0] PIPETX4SYNCHEADER_out;
  wire [1:0] PIPETX5CHARISK_out;
  wire [1:0] PIPETX5EQCONTROL_out;
  wire [1:0] PIPETX5POWERDOWN_out;
  wire [1:0] PIPETX5RATE_out;
  wire [1:0] PIPETX5SYNCHEADER_out;
  wire [1:0] PIPETX6CHARISK_out;
  wire [1:0] PIPETX6EQCONTROL_out;
  wire [1:0] PIPETX6POWERDOWN_out;
  wire [1:0] PIPETX6RATE_out;
  wire [1:0] PIPETX6SYNCHEADER_out;
  wire [1:0] PIPETX7CHARISK_out;
  wire [1:0] PIPETX7EQCONTROL_out;
  wire [1:0] PIPETX7POWERDOWN_out;
  wire [1:0] PIPETX7RATE_out;
  wire [1:0] PIPETX7SYNCHEADER_out;
  wire [1:0] PLEQPHASE_out;
  wire [23:0] CFGVFPOWERSTATE_out;
  wire [23:0] CFGVFTPHSTMODE_out;
  wire [255:0] LL2LMMAXISRXTDATA_out;
  wire [255:0] MAXISCQTDATA_out;
  wire [255:0] MAXISRCTDATA_out;
  wire [2:0] CFGCURRENTSPEED_out;
  wire [2:0] CFGMAXPAYLOAD_out;
  wire [2:0] CFGMAXREADREQ_out;
  wire [2:0] PIPERX0EQPRESET_out;
  wire [2:0] PIPERX1EQPRESET_out;
  wire [2:0] PIPERX2EQPRESET_out;
  wire [2:0] PIPERX3EQPRESET_out;
  wire [2:0] PIPERX4EQPRESET_out;
  wire [2:0] PIPERX5EQPRESET_out;
  wire [2:0] PIPERX6EQPRESET_out;
  wire [2:0] PIPERX7EQPRESET_out;
  wire [2:0] PIPETX0MARGIN_out;
  wire [2:0] PIPETX1MARGIN_out;
  wire [2:0] PIPETX2MARGIN_out;
  wire [2:0] PIPETX3MARGIN_out;
  wire [2:0] PIPETX4MARGIN_out;
  wire [2:0] PIPETX5MARGIN_out;
  wire [2:0] PIPETX6MARGIN_out;
  wire [2:0] PIPETX7MARGIN_out;
  wire [31:0] CFGEXTWRITEDATA_out;
  wire [31:0] CFGINTERRUPTMSIDATA_out;
  wire [31:0] CFGMGMTREADDATA_out;
  wire [31:0] CFGTPHSTTWRITEDATA_out;
  wire [31:0] CONFRESPRDATA_out;
  wire [31:0] DBGMCAPDATA_out;
  wire [31:0] PIPETX0DATA_out;
  wire [31:0] PIPETX1DATA_out;
  wire [31:0] PIPETX2DATA_out;
  wire [31:0] PIPETX3DATA_out;
  wire [31:0] PIPETX4DATA_out;
  wire [31:0] PIPETX5DATA_out;
  wire [31:0] PIPETX6DATA_out;
  wire [31:0] PIPETX7DATA_out;
  wire [31:0] SPAREOUT_out;
  wire [3:0] CFGDPASUBSTATECHANGE_out;
  wire [3:0] CFGEXTWRITEBYTEENABLE_out;
  wire [3:0] CFGFLRINPROCESS_out;
  wire [3:0] CFGINTERRUPTMSIENABLE_out;
  wire [3:0] CFGINTERRUPTMSIXENABLE_out;
  wire [3:0] CFGINTERRUPTMSIXMASK_out;
  wire [3:0] CFGNEGOTIATEDWIDTH_out;
  wire [3:0] CFGRCBSTATUS_out;
  wire [3:0] CFGTPHFUNCTIONNUM_out;
  wire [3:0] CFGTPHREQUESTERENABLE_out;
  wire [3:0] CFGTPHSTTWRITEBYTEVALID_out;
  wire [3:0] LL2LMMASTERTLPSENTTLPID0_out;
  wire [3:0] LL2LMMASTERTLPSENTTLPID1_out;
  wire [3:0] MICOMPLETIONRAMREADENABLEL_out;
  wire [3:0] MICOMPLETIONRAMREADENABLEU_out;
  wire [3:0] MICOMPLETIONRAMWRITEENABLEL_out;
  wire [3:0] MICOMPLETIONRAMWRITEENABLEU_out;
  wire [3:0] MIREQUESTRAMREADENABLE_out;
  wire [3:0] MIREQUESTRAMWRITEENABLE_out;
  wire [3:0] PCIERQSEQNUM_out;
  wire [3:0] PIPERX0EQLPTXPRESET_out;
  wire [3:0] PIPERX1EQLPTXPRESET_out;
  wire [3:0] PIPERX2EQLPTXPRESET_out;
  wire [3:0] PIPERX3EQLPTXPRESET_out;
  wire [3:0] PIPERX4EQLPTXPRESET_out;
  wire [3:0] PIPERX5EQLPTXPRESET_out;
  wire [3:0] PIPERX6EQLPTXPRESET_out;
  wire [3:0] PIPERX7EQLPTXPRESET_out;
  wire [3:0] PIPETX0EQPRESET_out;
  wire [3:0] PIPETX1EQPRESET_out;
  wire [3:0] PIPETX2EQPRESET_out;
  wire [3:0] PIPETX3EQPRESET_out;
  wire [3:0] PIPETX4EQPRESET_out;
  wire [3:0] PIPETX5EQPRESET_out;
  wire [3:0] PIPETX6EQPRESET_out;
  wire [3:0] PIPETX7EQPRESET_out;
  wire [3:0] SAXISCCTREADY_out;
  wire [3:0] SAXISRQTREADY_out;
  wire [479:0] XILUNCONNBOUT_out;
  wire [4:0] CFGMSGRECEIVEDTYPE_out;
  wire [4:0] CFGTPHSTTADDRESS_out;
  wire [5:0] CFGLTSSMSTATE_out;
  wire [5:0] PCIECQNPREQCOUNT_out;
  wire [5:0] PCIERQTAG_out;
  wire [5:0] PIPERX0EQLPLFFS_out;
  wire [5:0] PIPERX1EQLPLFFS_out;
  wire [5:0] PIPERX2EQLPLFFS_out;
  wire [5:0] PIPERX3EQLPLFFS_out;
  wire [5:0] PIPERX4EQLPLFFS_out;
  wire [5:0] PIPERX5EQLPLFFS_out;
  wire [5:0] PIPERX6EQLPLFFS_out;
  wire [5:0] PIPERX7EQLPLFFS_out;
  wire [5:0] PIPETX0EQDEEMPH_out;
  wire [5:0] PIPETX1EQDEEMPH_out;
  wire [5:0] PIPETX2EQDEEMPH_out;
  wire [5:0] PIPETX3EQDEEMPH_out;
  wire [5:0] PIPETX4EQDEEMPH_out;
  wire [5:0] PIPETX5EQDEEMPH_out;
  wire [5:0] PIPETX6EQDEEMPH_out;
  wire [5:0] PIPETX7EQDEEMPH_out;
  wire [71:0] MICOMPLETIONRAMWRITEDATAL_out;
  wire [71:0] MICOMPLETIONRAMWRITEDATAU_out;
  wire [74:0] MAXISRCTUSER_out;
  wire [7:0] CFGEXTFUNCTIONNUMBER_out;
  wire [7:0] CFGFCCPLH_out;
  wire [7:0] CFGFCNPH_out;
  wire [7:0] CFGFCPH_out;
  wire [7:0] CFGINTERRUPTMSIVFENABLE_out;
  wire [7:0] CFGINTERRUPTMSIXVFENABLE_out;
  wire [7:0] CFGINTERRUPTMSIXVFMASK_out;
  wire [7:0] CFGMSGRECEIVEDDATA_out;
  wire [7:0] CFGVFFLRINPROCESS_out;
  wire [7:0] CFGVFTPHREQUESTERENABLE_out;
  wire [7:0] DBGPLINFERREDRXELECTRICALIDLE_out;
  wire [7:0] LL2LMMAXISRXTVALID_out;
  wire [7:0] LL2LMSAXISTXTREADY_out;
  wire [7:0] MAXISCQTKEEP_out;
  wire [7:0] MAXISRCTKEEP_out;
  wire [84:0] MAXISCQTUSER_out;
  wire [860:0] XILUNCONNOUT_out;
  wire [8:0] MIREPLAYRAMADDRESS_out;
  wire [8:0] MIREQUESTRAMREADADDRESSA_out;
  wire [8:0] MIREQUESTRAMREADADDRESSB_out;
  wire [8:0] MIREQUESTRAMWRITEADDRESSA_out;
  wire [8:0] MIREQUESTRAMWRITEADDRESSB_out;
  wire [95:0] SCANOUT_out;
  wire [9:0] CFGEXTREGISTERNUMBER_out;
  wire [9:0] MICOMPLETIONRAMREADADDRESSAL_out;
  wire [9:0] MICOMPLETIONRAMREADADDRESSAU_out;
  wire [9:0] MICOMPLETIONRAMREADADDRESSBL_out;
  wire [9:0] MICOMPLETIONRAMREADADDRESSBU_out;
  wire [9:0] MICOMPLETIONRAMWRITEADDRESSAL_out;
  wire [9:0] MICOMPLETIONRAMWRITEADDRESSAU_out;
  wire [9:0] MICOMPLETIONRAMWRITEADDRESSBL_out;
  wire [9:0] MICOMPLETIONRAMWRITEADDRESSBU_out;

  wire CFGERRCOROUT_delay;
  wire CFGERRFATALOUT_delay;
  wire CFGERRNONFATALOUT_delay;
  wire CFGEXTREADRECEIVED_delay;
  wire CFGEXTWRITERECEIVED_delay;
  wire CFGHOTRESETOUT_delay;
  wire CFGINTERRUPTMSIFAIL_delay;
  wire CFGINTERRUPTMSIMASKUPDATE_delay;
  wire CFGINTERRUPTMSISENT_delay;
  wire CFGINTERRUPTMSIXFAIL_delay;
  wire CFGINTERRUPTMSIXSENT_delay;
  wire CFGINTERRUPTSENT_delay;
  wire CFGLOCALERROR_delay;
  wire CFGLTRENABLE_delay;
  wire CFGMGMTREADWRITEDONE_delay;
  wire CFGMSGRECEIVED_delay;
  wire CFGMSGTRANSMITDONE_delay;
  wire CFGPERFUNCTIONUPDATEDONE_delay;
  wire CFGPHYLINKDOWN_delay;
  wire CFGPLSTATUSCHANGE_delay;
  wire CFGPOWERSTATECHANGEINTERRUPT_delay;
  wire CFGTPHSTTREADENABLE_delay;
  wire CFGTPHSTTWRITEENABLE_delay;
  wire CONFMCAPDESIGNSWITCH_delay;
  wire CONFMCAPEOS_delay;
  wire CONFMCAPINUSEBYPCIE_delay;
  wire CONFREQREADY_delay;
  wire CONFRESPVALID_delay;
  wire DBGMCAPCSB_delay;
  wire DBGMCAPEOS_delay;
  wire DBGMCAPERROR_delay;
  wire DBGMCAPMODE_delay;
  wire DBGMCAPRDATAVALID_delay;
  wire DBGMCAPRDWRB_delay;
  wire DBGMCAPRESET_delay;
  wire DBGPLDATABLOCKRECEIVEDAFTEREDS_delay;
  wire DBGPLGEN3FRAMINGERRORDETECTED_delay;
  wire DBGPLGEN3SYNCHEADERERRORDETECTED_delay;
  wire DRPRDY_delay;
  wire LL2LMMASTERTLPSENT0_delay;
  wire LL2LMMASTERTLPSENT1_delay;
  wire MAXISCQTLAST_delay;
  wire MAXISCQTVALID_delay;
  wire MAXISRCTLAST_delay;
  wire MAXISRCTVALID_delay;
  wire PCIEPERST0B_delay;
  wire PCIEPERST1B_delay;
  wire PCIERQSEQNUMVLD_delay;
  wire PCIERQTAGVLD_delay;
  wire PIPERX0POLARITY_delay;
  wire PIPERX1POLARITY_delay;
  wire PIPERX2POLARITY_delay;
  wire PIPERX3POLARITY_delay;
  wire PIPERX4POLARITY_delay;
  wire PIPERX5POLARITY_delay;
  wire PIPERX6POLARITY_delay;
  wire PIPERX7POLARITY_delay;
  wire PIPETX0COMPLIANCE_delay;
  wire PIPETX0DATAVALID_delay;
  wire PIPETX0DEEMPH_delay;
  wire PIPETX0ELECIDLE_delay;
  wire PIPETX0RCVRDET_delay;
  wire PIPETX0RESET_delay;
  wire PIPETX0STARTBLOCK_delay;
  wire PIPETX0SWING_delay;
  wire PIPETX1COMPLIANCE_delay;
  wire PIPETX1DATAVALID_delay;
  wire PIPETX1DEEMPH_delay;
  wire PIPETX1ELECIDLE_delay;
  wire PIPETX1RCVRDET_delay;
  wire PIPETX1RESET_delay;
  wire PIPETX1STARTBLOCK_delay;
  wire PIPETX1SWING_delay;
  wire PIPETX2COMPLIANCE_delay;
  wire PIPETX2DATAVALID_delay;
  wire PIPETX2DEEMPH_delay;
  wire PIPETX2ELECIDLE_delay;
  wire PIPETX2RCVRDET_delay;
  wire PIPETX2RESET_delay;
  wire PIPETX2STARTBLOCK_delay;
  wire PIPETX2SWING_delay;
  wire PIPETX3COMPLIANCE_delay;
  wire PIPETX3DATAVALID_delay;
  wire PIPETX3DEEMPH_delay;
  wire PIPETX3ELECIDLE_delay;
  wire PIPETX3RCVRDET_delay;
  wire PIPETX3RESET_delay;
  wire PIPETX3STARTBLOCK_delay;
  wire PIPETX3SWING_delay;
  wire PIPETX4COMPLIANCE_delay;
  wire PIPETX4DATAVALID_delay;
  wire PIPETX4DEEMPH_delay;
  wire PIPETX4ELECIDLE_delay;
  wire PIPETX4RCVRDET_delay;
  wire PIPETX4RESET_delay;
  wire PIPETX4STARTBLOCK_delay;
  wire PIPETX4SWING_delay;
  wire PIPETX5COMPLIANCE_delay;
  wire PIPETX5DATAVALID_delay;
  wire PIPETX5DEEMPH_delay;
  wire PIPETX5ELECIDLE_delay;
  wire PIPETX5RCVRDET_delay;
  wire PIPETX5RESET_delay;
  wire PIPETX5STARTBLOCK_delay;
  wire PIPETX5SWING_delay;
  wire PIPETX6COMPLIANCE_delay;
  wire PIPETX6DATAVALID_delay;
  wire PIPETX6DEEMPH_delay;
  wire PIPETX6ELECIDLE_delay;
  wire PIPETX6RCVRDET_delay;
  wire PIPETX6RESET_delay;
  wire PIPETX6STARTBLOCK_delay;
  wire PIPETX6SWING_delay;
  wire PIPETX7COMPLIANCE_delay;
  wire PIPETX7DATAVALID_delay;
  wire PIPETX7DEEMPH_delay;
  wire PIPETX7ELECIDLE_delay;
  wire PIPETX7RCVRDET_delay;
  wire PIPETX7RESET_delay;
  wire PIPETX7STARTBLOCK_delay;
  wire PIPETX7SWING_delay;
  wire PLEQINPROGRESS_delay;
  wire [11:0] CFGFCCPLD_delay;
  wire [11:0] CFGFCNPD_delay;
  wire [11:0] CFGFCPD_delay;
  wire [11:0] CFGFUNCTIONPOWERSTATE_delay;
  wire [11:0] CFGINTERRUPTMSIMMENABLE_delay;
  wire [11:0] CFGTPHSTMODE_delay;
  wire [143:0] MIREPLAYRAMWRITEDATA_delay;
  wire [143:0] MIREQUESTRAMWRITEDATA_delay;
  wire [15:0] CFGFUNCTIONSTATUS_delay;
  wire [15:0] CFGPERFUNCSTATUSDATA_delay;
  wire [15:0] CFGVFSTATUS_delay;
  wire [15:0] DBGDATAOUT_delay;
  wire [15:0] DRPDO_delay;
  wire [17:0] LL2LMMAXISRXTUSER_delay;
  wire [1:0] CFGLINKPOWERSTATE_delay;
  wire [1:0] CFGOBFFENABLE_delay;
  wire [1:0] CFGPHYLINKSTATUS_delay;
  wire [1:0] MIREPLAYRAMREADENABLE_delay;
  wire [1:0] MIREPLAYRAMWRITEENABLE_delay;
  wire [1:0] PCIERQTAGAV_delay;
  wire [1:0] PCIETFCNPDAV_delay;
  wire [1:0] PCIETFCNPHAV_delay;
  wire [1:0] PIPERX0EQCONTROL_delay;
  wire [1:0] PIPERX1EQCONTROL_delay;
  wire [1:0] PIPERX2EQCONTROL_delay;
  wire [1:0] PIPERX3EQCONTROL_delay;
  wire [1:0] PIPERX4EQCONTROL_delay;
  wire [1:0] PIPERX5EQCONTROL_delay;
  wire [1:0] PIPERX6EQCONTROL_delay;
  wire [1:0] PIPERX7EQCONTROL_delay;
  wire [1:0] PIPETX0CHARISK_delay;
  wire [1:0] PIPETX0EQCONTROL_delay;
  wire [1:0] PIPETX0POWERDOWN_delay;
  wire [1:0] PIPETX0RATE_delay;
  wire [1:0] PIPETX0SYNCHEADER_delay;
  wire [1:0] PIPETX1CHARISK_delay;
  wire [1:0] PIPETX1EQCONTROL_delay;
  wire [1:0] PIPETX1POWERDOWN_delay;
  wire [1:0] PIPETX1RATE_delay;
  wire [1:0] PIPETX1SYNCHEADER_delay;
  wire [1:0] PIPETX2CHARISK_delay;
  wire [1:0] PIPETX2EQCONTROL_delay;
  wire [1:0] PIPETX2POWERDOWN_delay;
  wire [1:0] PIPETX2RATE_delay;
  wire [1:0] PIPETX2SYNCHEADER_delay;
  wire [1:0] PIPETX3CHARISK_delay;
  wire [1:0] PIPETX3EQCONTROL_delay;
  wire [1:0] PIPETX3POWERDOWN_delay;
  wire [1:0] PIPETX3RATE_delay;
  wire [1:0] PIPETX3SYNCHEADER_delay;
  wire [1:0] PIPETX4CHARISK_delay;
  wire [1:0] PIPETX4EQCONTROL_delay;
  wire [1:0] PIPETX4POWERDOWN_delay;
  wire [1:0] PIPETX4RATE_delay;
  wire [1:0] PIPETX4SYNCHEADER_delay;
  wire [1:0] PIPETX5CHARISK_delay;
  wire [1:0] PIPETX5EQCONTROL_delay;
  wire [1:0] PIPETX5POWERDOWN_delay;
  wire [1:0] PIPETX5RATE_delay;
  wire [1:0] PIPETX5SYNCHEADER_delay;
  wire [1:0] PIPETX6CHARISK_delay;
  wire [1:0] PIPETX6EQCONTROL_delay;
  wire [1:0] PIPETX6POWERDOWN_delay;
  wire [1:0] PIPETX6RATE_delay;
  wire [1:0] PIPETX6SYNCHEADER_delay;
  wire [1:0] PIPETX7CHARISK_delay;
  wire [1:0] PIPETX7EQCONTROL_delay;
  wire [1:0] PIPETX7POWERDOWN_delay;
  wire [1:0] PIPETX7RATE_delay;
  wire [1:0] PIPETX7SYNCHEADER_delay;
  wire [1:0] PLEQPHASE_delay;
  wire [23:0] CFGVFPOWERSTATE_delay;
  wire [23:0] CFGVFTPHSTMODE_delay;
  wire [255:0] LL2LMMAXISRXTDATA_delay;
  wire [255:0] MAXISCQTDATA_delay;
  wire [255:0] MAXISRCTDATA_delay;
  wire [2:0] CFGCURRENTSPEED_delay;
  wire [2:0] CFGMAXPAYLOAD_delay;
  wire [2:0] CFGMAXREADREQ_delay;
  wire [2:0] PIPERX0EQPRESET_delay;
  wire [2:0] PIPERX1EQPRESET_delay;
  wire [2:0] PIPERX2EQPRESET_delay;
  wire [2:0] PIPERX3EQPRESET_delay;
  wire [2:0] PIPERX4EQPRESET_delay;
  wire [2:0] PIPERX5EQPRESET_delay;
  wire [2:0] PIPERX6EQPRESET_delay;
  wire [2:0] PIPERX7EQPRESET_delay;
  wire [2:0] PIPETX0MARGIN_delay;
  wire [2:0] PIPETX1MARGIN_delay;
  wire [2:0] PIPETX2MARGIN_delay;
  wire [2:0] PIPETX3MARGIN_delay;
  wire [2:0] PIPETX4MARGIN_delay;
  wire [2:0] PIPETX5MARGIN_delay;
  wire [2:0] PIPETX6MARGIN_delay;
  wire [2:0] PIPETX7MARGIN_delay;
  wire [31:0] CFGEXTWRITEDATA_delay;
  wire [31:0] CFGINTERRUPTMSIDATA_delay;
  wire [31:0] CFGMGMTREADDATA_delay;
  wire [31:0] CFGTPHSTTWRITEDATA_delay;
  wire [31:0] CONFRESPRDATA_delay;
  wire [31:0] DBGMCAPDATA_delay;
  wire [31:0] PIPETX0DATA_delay;
  wire [31:0] PIPETX1DATA_delay;
  wire [31:0] PIPETX2DATA_delay;
  wire [31:0] PIPETX3DATA_delay;
  wire [31:0] PIPETX4DATA_delay;
  wire [31:0] PIPETX5DATA_delay;
  wire [31:0] PIPETX6DATA_delay;
  wire [31:0] PIPETX7DATA_delay;
  wire [31:0] SPAREOUT_delay;
  wire [3:0] CFGDPASUBSTATECHANGE_delay;
  wire [3:0] CFGEXTWRITEBYTEENABLE_delay;
  wire [3:0] CFGFLRINPROCESS_delay;
  wire [3:0] CFGINTERRUPTMSIENABLE_delay;
  wire [3:0] CFGINTERRUPTMSIXENABLE_delay;
  wire [3:0] CFGINTERRUPTMSIXMASK_delay;
  wire [3:0] CFGNEGOTIATEDWIDTH_delay;
  wire [3:0] CFGRCBSTATUS_delay;
  wire [3:0] CFGTPHFUNCTIONNUM_delay;
  wire [3:0] CFGTPHREQUESTERENABLE_delay;
  wire [3:0] CFGTPHSTTWRITEBYTEVALID_delay;
  wire [3:0] LL2LMMASTERTLPSENTTLPID0_delay;
  wire [3:0] LL2LMMASTERTLPSENTTLPID1_delay;
  wire [3:0] MICOMPLETIONRAMREADENABLEL_delay;
  wire [3:0] MICOMPLETIONRAMREADENABLEU_delay;
  wire [3:0] MICOMPLETIONRAMWRITEENABLEL_delay;
  wire [3:0] MICOMPLETIONRAMWRITEENABLEU_delay;
  wire [3:0] MIREQUESTRAMREADENABLE_delay;
  wire [3:0] MIREQUESTRAMWRITEENABLE_delay;
  wire [3:0] PCIERQSEQNUM_delay;
  wire [3:0] PIPERX0EQLPTXPRESET_delay;
  wire [3:0] PIPERX1EQLPTXPRESET_delay;
  wire [3:0] PIPERX2EQLPTXPRESET_delay;
  wire [3:0] PIPERX3EQLPTXPRESET_delay;
  wire [3:0] PIPERX4EQLPTXPRESET_delay;
  wire [3:0] PIPERX5EQLPTXPRESET_delay;
  wire [3:0] PIPERX6EQLPTXPRESET_delay;
  wire [3:0] PIPERX7EQLPTXPRESET_delay;
  wire [3:0] PIPETX0EQPRESET_delay;
  wire [3:0] PIPETX1EQPRESET_delay;
  wire [3:0] PIPETX2EQPRESET_delay;
  wire [3:0] PIPETX3EQPRESET_delay;
  wire [3:0] PIPETX4EQPRESET_delay;
  wire [3:0] PIPETX5EQPRESET_delay;
  wire [3:0] PIPETX6EQPRESET_delay;
  wire [3:0] PIPETX7EQPRESET_delay;
  wire [3:0] SAXISCCTREADY_delay;
  wire [3:0] SAXISRQTREADY_delay;
  wire [4:0] CFGMSGRECEIVEDTYPE_delay;
  wire [4:0] CFGTPHSTTADDRESS_delay;
  wire [5:0] CFGLTSSMSTATE_delay;
  wire [5:0] PCIECQNPREQCOUNT_delay;
  wire [5:0] PCIERQTAG_delay;
  wire [5:0] PIPERX0EQLPLFFS_delay;
  wire [5:0] PIPERX1EQLPLFFS_delay;
  wire [5:0] PIPERX2EQLPLFFS_delay;
  wire [5:0] PIPERX3EQLPLFFS_delay;
  wire [5:0] PIPERX4EQLPLFFS_delay;
  wire [5:0] PIPERX5EQLPLFFS_delay;
  wire [5:0] PIPERX6EQLPLFFS_delay;
  wire [5:0] PIPERX7EQLPLFFS_delay;
  wire [5:0] PIPETX0EQDEEMPH_delay;
  wire [5:0] PIPETX1EQDEEMPH_delay;
  wire [5:0] PIPETX2EQDEEMPH_delay;
  wire [5:0] PIPETX3EQDEEMPH_delay;
  wire [5:0] PIPETX4EQDEEMPH_delay;
  wire [5:0] PIPETX5EQDEEMPH_delay;
  wire [5:0] PIPETX6EQDEEMPH_delay;
  wire [5:0] PIPETX7EQDEEMPH_delay;
  wire [71:0] MICOMPLETIONRAMWRITEDATAL_delay;
  wire [71:0] MICOMPLETIONRAMWRITEDATAU_delay;
  wire [74:0] MAXISRCTUSER_delay;
  wire [7:0] CFGEXTFUNCTIONNUMBER_delay;
  wire [7:0] CFGFCCPLH_delay;
  wire [7:0] CFGFCNPH_delay;
  wire [7:0] CFGFCPH_delay;
  wire [7:0] CFGINTERRUPTMSIVFENABLE_delay;
  wire [7:0] CFGINTERRUPTMSIXVFENABLE_delay;
  wire [7:0] CFGINTERRUPTMSIXVFMASK_delay;
  wire [7:0] CFGMSGRECEIVEDDATA_delay;
  wire [7:0] CFGVFFLRINPROCESS_delay;
  wire [7:0] CFGVFTPHREQUESTERENABLE_delay;
  wire [7:0] DBGPLINFERREDRXELECTRICALIDLE_delay;
  wire [7:0] LL2LMMAXISRXTVALID_delay;
  wire [7:0] LL2LMSAXISTXTREADY_delay;
  wire [7:0] MAXISCQTKEEP_delay;
  wire [7:0] MAXISRCTKEEP_delay;
  wire [84:0] MAXISCQTUSER_delay;
  wire [8:0] MIREPLAYRAMADDRESS_delay;
  wire [8:0] MIREQUESTRAMREADADDRESSA_delay;
  wire [8:0] MIREQUESTRAMREADADDRESSB_delay;
  wire [8:0] MIREQUESTRAMWRITEADDRESSA_delay;
  wire [8:0] MIREQUESTRAMWRITEADDRESSB_delay;
  wire [9:0] CFGEXTREGISTERNUMBER_delay;
  wire [9:0] MICOMPLETIONRAMREADADDRESSAL_delay;
  wire [9:0] MICOMPLETIONRAMREADADDRESSAU_delay;
  wire [9:0] MICOMPLETIONRAMREADADDRESSBL_delay;
  wire [9:0] MICOMPLETIONRAMREADADDRESSBU_delay;
  wire [9:0] MICOMPLETIONRAMWRITEADDRESSAL_delay;
  wire [9:0] MICOMPLETIONRAMWRITEADDRESSAU_delay;
  wire [9:0] MICOMPLETIONRAMWRITEADDRESSBL_delay;
  wire [9:0] MICOMPLETIONRAMWRITEADDRESSBU_delay;

  wire CFGCONFIGSPACEENABLE_in;
  wire CFGERRCORIN_in;
  wire CFGERRUNCORIN_in;
  wire CFGEXTREADDATAVALID_in;
  wire CFGHOTRESETIN_in;
  wire CFGINTERRUPTMSIPENDINGSTATUSDATAENABLE_in;
  wire CFGINTERRUPTMSITPHPRESENT_in;
  wire CFGINTERRUPTMSIXINT_in;
  wire CFGLINKTRAININGENABLE_in;
  wire CFGMGMTREAD_in;
  wire CFGMGMTTYPE1CFGREGACCESS_in;
  wire CFGMGMTWRITE_in;
  wire CFGMSGTRANSMIT_in;
  wire CFGPERFUNCTIONOUTPUTREQUEST_in;
  wire CFGPOWERSTATECHANGEACK_in;
  wire CFGREQPMTRANSITIONL23READY_in;
  wire CFGTPHSTTREADDATAVALID_in;
  wire CONFMCAPREQUESTBYCONF_in;
  wire CONFREQVALID_in;
  wire CORECLKMICOMPLETIONRAML_in;
  wire CORECLKMICOMPLETIONRAMU_in;
  wire CORECLKMIREPLAYRAM_in;
  wire CORECLKMIREQUESTRAM_in;
  wire CORECLK_in;
  wire DBGCFGLOCALMGMTREGOVERRIDE_in;
  wire DRPCLK_in;
  wire DRPEN_in;
  wire DRPWE_in;
  wire LL2LMSAXISTXTVALID_in;
  wire MCAPCLK_in;
  wire MCAPPERST0B_in;
  wire MCAPPERST1B_in;
  wire MGMTRESETN_in;
  wire MGMTSTICKYRESETN_in;
  wire PCIECQNPREQ_in;
  wire PIPECLK_in;
  wire PIPERESETN_in;
  wire PIPERX0DATAVALID_in;
  wire PIPERX0ELECIDLE_in;
  wire PIPERX0EQDONE_in;
  wire PIPERX0EQLPADAPTDONE_in;
  wire PIPERX0EQLPLFFSSEL_in;
  wire PIPERX0PHYSTATUS_in;
  wire PIPERX0STARTBLOCK_in;
  wire PIPERX0VALID_in;
  wire PIPERX1DATAVALID_in;
  wire PIPERX1ELECIDLE_in;
  wire PIPERX1EQDONE_in;
  wire PIPERX1EQLPADAPTDONE_in;
  wire PIPERX1EQLPLFFSSEL_in;
  wire PIPERX1PHYSTATUS_in;
  wire PIPERX1STARTBLOCK_in;
  wire PIPERX1VALID_in;
  wire PIPERX2DATAVALID_in;
  wire PIPERX2ELECIDLE_in;
  wire PIPERX2EQDONE_in;
  wire PIPERX2EQLPADAPTDONE_in;
  wire PIPERX2EQLPLFFSSEL_in;
  wire PIPERX2PHYSTATUS_in;
  wire PIPERX2STARTBLOCK_in;
  wire PIPERX2VALID_in;
  wire PIPERX3DATAVALID_in;
  wire PIPERX3ELECIDLE_in;
  wire PIPERX3EQDONE_in;
  wire PIPERX3EQLPADAPTDONE_in;
  wire PIPERX3EQLPLFFSSEL_in;
  wire PIPERX3PHYSTATUS_in;
  wire PIPERX3STARTBLOCK_in;
  wire PIPERX3VALID_in;
  wire PIPERX4DATAVALID_in;
  wire PIPERX4ELECIDLE_in;
  wire PIPERX4EQDONE_in;
  wire PIPERX4EQLPADAPTDONE_in;
  wire PIPERX4EQLPLFFSSEL_in;
  wire PIPERX4PHYSTATUS_in;
  wire PIPERX4STARTBLOCK_in;
  wire PIPERX4VALID_in;
  wire PIPERX5DATAVALID_in;
  wire PIPERX5ELECIDLE_in;
  wire PIPERX5EQDONE_in;
  wire PIPERX5EQLPADAPTDONE_in;
  wire PIPERX5EQLPLFFSSEL_in;
  wire PIPERX5PHYSTATUS_in;
  wire PIPERX5STARTBLOCK_in;
  wire PIPERX5VALID_in;
  wire PIPERX6DATAVALID_in;
  wire PIPERX6ELECIDLE_in;
  wire PIPERX6EQDONE_in;
  wire PIPERX6EQLPADAPTDONE_in;
  wire PIPERX6EQLPLFFSSEL_in;
  wire PIPERX6PHYSTATUS_in;
  wire PIPERX6STARTBLOCK_in;
  wire PIPERX6VALID_in;
  wire PIPERX7DATAVALID_in;
  wire PIPERX7ELECIDLE_in;
  wire PIPERX7EQDONE_in;
  wire PIPERX7EQLPADAPTDONE_in;
  wire PIPERX7EQLPLFFSSEL_in;
  wire PIPERX7PHYSTATUS_in;
  wire PIPERX7STARTBLOCK_in;
  wire PIPERX7VALID_in;
  wire PIPETX0EQDONE_in;
  wire PIPETX1EQDONE_in;
  wire PIPETX2EQDONE_in;
  wire PIPETX3EQDONE_in;
  wire PIPETX4EQDONE_in;
  wire PIPETX5EQDONE_in;
  wire PIPETX6EQDONE_in;
  wire PIPETX7EQDONE_in;
  wire PLEQRESETEIEOSCOUNT_in;
  wire PLGEN2UPSTREAMPREFERDEEMPH_in;
  wire PMVENABLEN_in;
  wire RESETN_in;
  wire SAXISCCTLAST_in;
  wire SAXISCCTVALID_in;
  wire SAXISRQTLAST_in;
  wire SAXISRQTVALID_in;
  wire SCANENABLEN_in;
  wire SCANMODEN_in;
  wire USERCLK_in;
  wire [13:0] LL2LMSAXISTXTUSER_in;
  wire [143:0] MICOMPLETIONRAMREADDATA_in;
  wire [143:0] MIREPLAYRAMREADDATA_in;
  wire [143:0] MIREQUESTRAMREADDATA_in;
  wire [15:0] CFGDEVID_in;
  wire [15:0] CFGSUBSYSID_in;
  wire [15:0] CFGSUBSYSVENDID_in;
  wire [15:0] CFGVENDID_in;
  wire [15:0] DRPDI_in;
  wire [17:0] PIPERX0EQLPNEWTXCOEFFORPRESET_in;
  wire [17:0] PIPERX1EQLPNEWTXCOEFFORPRESET_in;
  wire [17:0] PIPERX2EQLPNEWTXCOEFFORPRESET_in;
  wire [17:0] PIPERX3EQLPNEWTXCOEFFORPRESET_in;
  wire [17:0] PIPERX4EQLPNEWTXCOEFFORPRESET_in;
  wire [17:0] PIPERX5EQLPNEWTXCOEFFORPRESET_in;
  wire [17:0] PIPERX6EQLPNEWTXCOEFFORPRESET_in;
  wire [17:0] PIPERX7EQLPNEWTXCOEFFORPRESET_in;
  wire [17:0] PIPETX0EQCOEFF_in;
  wire [17:0] PIPETX1EQCOEFF_in;
  wire [17:0] PIPETX2EQCOEFF_in;
  wire [17:0] PIPETX3EQCOEFF_in;
  wire [17:0] PIPETX4EQCOEFF_in;
  wire [17:0] PIPETX5EQCOEFF_in;
  wire [17:0] PIPETX6EQCOEFF_in;
  wire [17:0] PIPETX7EQCOEFF_in;
  wire [18:0] CFGMGMTADDR_in;
  wire [1919:0] XILUNCONNBYP_in;
  wire [1:0] CFGINTERRUPTMSITPHTYPE_in;
  wire [1:0] CONFREQTYPE_in;
  wire [1:0] PIPERX0CHARISK_in;
  wire [1:0] PIPERX0SYNCHEADER_in;
  wire [1:0] PIPERX1CHARISK_in;
  wire [1:0] PIPERX1SYNCHEADER_in;
  wire [1:0] PIPERX2CHARISK_in;
  wire [1:0] PIPERX2SYNCHEADER_in;
  wire [1:0] PIPERX3CHARISK_in;
  wire [1:0] PIPERX3SYNCHEADER_in;
  wire [1:0] PIPERX4CHARISK_in;
  wire [1:0] PIPERX4SYNCHEADER_in;
  wire [1:0] PIPERX5CHARISK_in;
  wire [1:0] PIPERX5SYNCHEADER_in;
  wire [1:0] PIPERX6CHARISK_in;
  wire [1:0] PIPERX6SYNCHEADER_in;
  wire [1:0] PIPERX7CHARISK_in;
  wire [1:0] PIPERX7SYNCHEADER_in;
  wire [1:0] PMVDIVIDE_in;
  wire [21:0] MAXISCQTREADY_in;
  wire [21:0] MAXISRCTREADY_in;
  wire [255:0] SAXISCCTDATA_in;
  wire [255:0] SAXISRQTDATA_in;
  wire [2:0] CFGDSFUNCTIONNUMBER_in;
  wire [2:0] CFGFCSEL_in;
  wire [2:0] CFGINTERRUPTMSIATTR_in;
  wire [2:0] CFGMSGTRANSMITTYPE_in;
  wire [2:0] CFGPERFUNCSTATUSCONTROL_in;
  wire [2:0] PIPERX0STATUS_in;
  wire [2:0] PIPERX1STATUS_in;
  wire [2:0] PIPERX2STATUS_in;
  wire [2:0] PIPERX3STATUS_in;
  wire [2:0] PIPERX4STATUS_in;
  wire [2:0] PIPERX5STATUS_in;
  wire [2:0] PIPERX6STATUS_in;
  wire [2:0] PIPERX7STATUS_in;
  wire [2:0] PMVSELECT_in;
  wire [3188:0] XILUNCONNIN_in;
  wire [31:0] CFGEXTREADDATA_in;
  wire [31:0] CFGINTERRUPTMSIINT_in;
  wire [31:0] CFGINTERRUPTMSIPENDINGSTATUS_in;
  wire [31:0] CFGINTERRUPTMSIXDATA_in;
  wire [31:0] CFGMGMTWRITEDATA_in;
  wire [31:0] CFGMSGTRANSMITDATA_in;
  wire [31:0] CFGTPHSTTREADDATA_in;
  wire [31:0] CONFREQDATA_in;
  wire [31:0] PIPERX0DATA_in;
  wire [31:0] PIPERX1DATA_in;
  wire [31:0] PIPERX2DATA_in;
  wire [31:0] PIPERX3DATA_in;
  wire [31:0] PIPERX4DATA_in;
  wire [31:0] PIPERX5DATA_in;
  wire [31:0] PIPERX6DATA_in;
  wire [31:0] PIPERX7DATA_in;
  wire [31:0] SPAREIN_in;
  wire [32:0] SAXISCCTUSER_in;
  wire [3:0] CFGFLRDONE_in;
  wire [3:0] CFGINTERRUPTINT_in;
  wire [3:0] CFGINTERRUPTMSIFUNCTIONNUMBER_in;
  wire [3:0] CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM_in;
  wire [3:0] CFGINTERRUPTMSISELECT_in;
  wire [3:0] CFGINTERRUPTPENDING_in;
  wire [3:0] CFGMGMTBYTEENABLE_in;
  wire [3:0] CFGPERFUNCTIONNUMBER_in;
  wire [3:0] CONFREQREGNUM_in;
  wire [3:0] DBGDATASEL_in;
  wire [3:0] LL2LMTXTLPID0_in;
  wire [3:0] LL2LMTXTLPID1_in;
  wire [4:0] CFGDSDEVICENUMBER_in;
  wire [59:0] SAXISRQTUSER_in;
  wire [5:0] PIPEEQFS_in;
  wire [5:0] PIPEEQLF_in;
  wire [63:0] CFGDSN_in;
  wire [63:0] CFGINTERRUPTMSIXADDRESS_in;
  wire [7:0] CFGDSBUSNUMBER_in;
  wire [7:0] CFGDSPORTNUMBER_in;
  wire [7:0] CFGREVID_in;
  wire [7:0] CFGVFFLRDONE_in;
  wire [7:0] SAXISCCTKEEP_in;
  wire [7:0] SAXISRQTKEEP_in;
  wire [8:0] CFGINTERRUPTMSITPHSTTAG_in;
  wire [950:0] XILUNCONNCLK_in;
  wire [95:0] SCANIN_in;
  wire [9:0] DRPADDR_in;

  wire CFGCONFIGSPACEENABLE_delay;
  wire CFGERRCORIN_delay;
  wire CFGERRUNCORIN_delay;
  wire CFGEXTREADDATAVALID_delay;
  wire CFGHOTRESETIN_delay;
  wire CFGINTERRUPTMSIPENDINGSTATUSDATAENABLE_delay;
  wire CFGINTERRUPTMSITPHPRESENT_delay;
  wire CFGINTERRUPTMSIXINT_delay;
  wire CFGLINKTRAININGENABLE_delay;
  wire CFGMGMTREAD_delay;
  wire CFGMGMTTYPE1CFGREGACCESS_delay;
  wire CFGMGMTWRITE_delay;
  wire CFGMSGTRANSMIT_delay;
  wire CFGPERFUNCTIONOUTPUTREQUEST_delay;
  wire CFGPOWERSTATECHANGEACK_delay;
  wire CFGREQPMTRANSITIONL23READY_delay;
  wire CFGTPHSTTREADDATAVALID_delay;
  wire CONFMCAPREQUESTBYCONF_delay;
  wire CONFREQVALID_delay;
  wire CORECLKMICOMPLETIONRAML_delay;
  wire CORECLKMICOMPLETIONRAMU_delay;
  wire CORECLKMIREPLAYRAM_delay;
  wire CORECLKMIREQUESTRAM_delay;
  wire CORECLK_delay;
  wire DBGCFGLOCALMGMTREGOVERRIDE_delay;
  wire DRPCLK_delay;
  wire DRPEN_delay;
  wire DRPWE_delay;
  wire LL2LMSAXISTXTVALID_delay;
  wire MCAPCLK_delay;
  wire MCAPPERST0B_delay;
  wire MCAPPERST1B_delay;
  wire MGMTRESETN_delay;
  wire MGMTSTICKYRESETN_delay;
  wire PCIECQNPREQ_delay;
  wire PIPECLK_delay;
  wire PIPERESETN_delay;
  wire PIPERX0DATAVALID_delay;
  wire PIPERX0ELECIDLE_delay;
  wire PIPERX0EQDONE_delay;
  wire PIPERX0EQLPADAPTDONE_delay;
  wire PIPERX0EQLPLFFSSEL_delay;
  wire PIPERX0PHYSTATUS_delay;
  wire PIPERX0STARTBLOCK_delay;
  wire PIPERX0VALID_delay;
  wire PIPERX1DATAVALID_delay;
  wire PIPERX1ELECIDLE_delay;
  wire PIPERX1EQDONE_delay;
  wire PIPERX1EQLPADAPTDONE_delay;
  wire PIPERX1EQLPLFFSSEL_delay;
  wire PIPERX1PHYSTATUS_delay;
  wire PIPERX1STARTBLOCK_delay;
  wire PIPERX1VALID_delay;
  wire PIPERX2DATAVALID_delay;
  wire PIPERX2ELECIDLE_delay;
  wire PIPERX2EQDONE_delay;
  wire PIPERX2EQLPADAPTDONE_delay;
  wire PIPERX2EQLPLFFSSEL_delay;
  wire PIPERX2PHYSTATUS_delay;
  wire PIPERX2STARTBLOCK_delay;
  wire PIPERX2VALID_delay;
  wire PIPERX3DATAVALID_delay;
  wire PIPERX3ELECIDLE_delay;
  wire PIPERX3EQDONE_delay;
  wire PIPERX3EQLPADAPTDONE_delay;
  wire PIPERX3EQLPLFFSSEL_delay;
  wire PIPERX3PHYSTATUS_delay;
  wire PIPERX3STARTBLOCK_delay;
  wire PIPERX3VALID_delay;
  wire PIPERX4DATAVALID_delay;
  wire PIPERX4ELECIDLE_delay;
  wire PIPERX4EQDONE_delay;
  wire PIPERX4EQLPADAPTDONE_delay;
  wire PIPERX4EQLPLFFSSEL_delay;
  wire PIPERX4PHYSTATUS_delay;
  wire PIPERX4STARTBLOCK_delay;
  wire PIPERX4VALID_delay;
  wire PIPERX5DATAVALID_delay;
  wire PIPERX5ELECIDLE_delay;
  wire PIPERX5EQDONE_delay;
  wire PIPERX5EQLPADAPTDONE_delay;
  wire PIPERX5EQLPLFFSSEL_delay;
  wire PIPERX5PHYSTATUS_delay;
  wire PIPERX5STARTBLOCK_delay;
  wire PIPERX5VALID_delay;
  wire PIPERX6DATAVALID_delay;
  wire PIPERX6ELECIDLE_delay;
  wire PIPERX6EQDONE_delay;
  wire PIPERX6EQLPADAPTDONE_delay;
  wire PIPERX6EQLPLFFSSEL_delay;
  wire PIPERX6PHYSTATUS_delay;
  wire PIPERX6STARTBLOCK_delay;
  wire PIPERX6VALID_delay;
  wire PIPERX7DATAVALID_delay;
  wire PIPERX7ELECIDLE_delay;
  wire PIPERX7EQDONE_delay;
  wire PIPERX7EQLPADAPTDONE_delay;
  wire PIPERX7EQLPLFFSSEL_delay;
  wire PIPERX7PHYSTATUS_delay;
  wire PIPERX7STARTBLOCK_delay;
  wire PIPERX7VALID_delay;
  wire PIPETX0EQDONE_delay;
  wire PIPETX1EQDONE_delay;
  wire PIPETX2EQDONE_delay;
  wire PIPETX3EQDONE_delay;
  wire PIPETX4EQDONE_delay;
  wire PIPETX5EQDONE_delay;
  wire PIPETX6EQDONE_delay;
  wire PIPETX7EQDONE_delay;
  wire PLEQRESETEIEOSCOUNT_delay;
  wire PLGEN2UPSTREAMPREFERDEEMPH_delay;
  wire RESETN_delay;
  wire SAXISCCTLAST_delay;
  wire SAXISCCTVALID_delay;
  wire SAXISRQTLAST_delay;
  wire SAXISRQTVALID_delay;
  wire USERCLK_delay;
  wire [13:0] LL2LMSAXISTXTUSER_delay;
  wire [143:0] MICOMPLETIONRAMREADDATA_delay;
  wire [143:0] MIREPLAYRAMREADDATA_delay;
  wire [143:0] MIREQUESTRAMREADDATA_delay;
  wire [15:0] CFGDEVID_delay;
  wire [15:0] CFGSUBSYSID_delay;
  wire [15:0] CFGSUBSYSVENDID_delay;
  wire [15:0] CFGVENDID_delay;
  wire [15:0] DRPDI_delay;
  wire [17:0] PIPERX0EQLPNEWTXCOEFFORPRESET_delay;
  wire [17:0] PIPERX1EQLPNEWTXCOEFFORPRESET_delay;
  wire [17:0] PIPERX2EQLPNEWTXCOEFFORPRESET_delay;
  wire [17:0] PIPERX3EQLPNEWTXCOEFFORPRESET_delay;
  wire [17:0] PIPERX4EQLPNEWTXCOEFFORPRESET_delay;
  wire [17:0] PIPERX5EQLPNEWTXCOEFFORPRESET_delay;
  wire [17:0] PIPERX6EQLPNEWTXCOEFFORPRESET_delay;
  wire [17:0] PIPERX7EQLPNEWTXCOEFFORPRESET_delay;
  wire [17:0] PIPETX0EQCOEFF_delay;
  wire [17:0] PIPETX1EQCOEFF_delay;
  wire [17:0] PIPETX2EQCOEFF_delay;
  wire [17:0] PIPETX3EQCOEFF_delay;
  wire [17:0] PIPETX4EQCOEFF_delay;
  wire [17:0] PIPETX5EQCOEFF_delay;
  wire [17:0] PIPETX6EQCOEFF_delay;
  wire [17:0] PIPETX7EQCOEFF_delay;
  wire [18:0] CFGMGMTADDR_delay;
  wire [1:0] CFGINTERRUPTMSITPHTYPE_delay;
  wire [1:0] CONFREQTYPE_delay;
  wire [1:0] PIPERX0CHARISK_delay;
  wire [1:0] PIPERX0SYNCHEADER_delay;
  wire [1:0] PIPERX1CHARISK_delay;
  wire [1:0] PIPERX1SYNCHEADER_delay;
  wire [1:0] PIPERX2CHARISK_delay;
  wire [1:0] PIPERX2SYNCHEADER_delay;
  wire [1:0] PIPERX3CHARISK_delay;
  wire [1:0] PIPERX3SYNCHEADER_delay;
  wire [1:0] PIPERX4CHARISK_delay;
  wire [1:0] PIPERX4SYNCHEADER_delay;
  wire [1:0] PIPERX5CHARISK_delay;
  wire [1:0] PIPERX5SYNCHEADER_delay;
  wire [1:0] PIPERX6CHARISK_delay;
  wire [1:0] PIPERX6SYNCHEADER_delay;
  wire [1:0] PIPERX7CHARISK_delay;
  wire [1:0] PIPERX7SYNCHEADER_delay;
  wire [21:0] MAXISCQTREADY_delay;
  wire [21:0] MAXISRCTREADY_delay;
  wire [255:0] SAXISCCTDATA_delay;
  wire [255:0] SAXISRQTDATA_delay;
  wire [2:0] CFGDSFUNCTIONNUMBER_delay;
  wire [2:0] CFGFCSEL_delay;
  wire [2:0] CFGINTERRUPTMSIATTR_delay;
  wire [2:0] CFGMSGTRANSMITTYPE_delay;
  wire [2:0] CFGPERFUNCSTATUSCONTROL_delay;
  wire [2:0] PIPERX0STATUS_delay;
  wire [2:0] PIPERX1STATUS_delay;
  wire [2:0] PIPERX2STATUS_delay;
  wire [2:0] PIPERX3STATUS_delay;
  wire [2:0] PIPERX4STATUS_delay;
  wire [2:0] PIPERX5STATUS_delay;
  wire [2:0] PIPERX6STATUS_delay;
  wire [2:0] PIPERX7STATUS_delay;
  wire [31:0] CFGEXTREADDATA_delay;
  wire [31:0] CFGINTERRUPTMSIINT_delay;
  wire [31:0] CFGINTERRUPTMSIPENDINGSTATUS_delay;
  wire [31:0] CFGINTERRUPTMSIXDATA_delay;
  wire [31:0] CFGMGMTWRITEDATA_delay;
  wire [31:0] CFGMSGTRANSMITDATA_delay;
  wire [31:0] CFGTPHSTTREADDATA_delay;
  wire [31:0] CONFREQDATA_delay;
  wire [31:0] PIPERX0DATA_delay;
  wire [31:0] PIPERX1DATA_delay;
  wire [31:0] PIPERX2DATA_delay;
  wire [31:0] PIPERX3DATA_delay;
  wire [31:0] PIPERX4DATA_delay;
  wire [31:0] PIPERX5DATA_delay;
  wire [31:0] PIPERX6DATA_delay;
  wire [31:0] PIPERX7DATA_delay;
  wire [31:0] SPAREIN_delay;
  wire [32:0] SAXISCCTUSER_delay;
  wire [3:0] CFGFLRDONE_delay;
  wire [3:0] CFGINTERRUPTINT_delay;
  wire [3:0] CFGINTERRUPTMSIFUNCTIONNUMBER_delay;
  wire [3:0] CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM_delay;
  wire [3:0] CFGINTERRUPTMSISELECT_delay;
  wire [3:0] CFGINTERRUPTPENDING_delay;
  wire [3:0] CFGMGMTBYTEENABLE_delay;
  wire [3:0] CFGPERFUNCTIONNUMBER_delay;
  wire [3:0] CONFREQREGNUM_delay;
  wire [3:0] DBGDATASEL_delay;
  wire [3:0] LL2LMTXTLPID0_delay;
  wire [3:0] LL2LMTXTLPID1_delay;
  wire [4:0] CFGDSDEVICENUMBER_delay;
  wire [59:0] SAXISRQTUSER_delay;
  wire [5:0] PIPEEQFS_delay;
  wire [5:0] PIPEEQLF_delay;
  wire [63:0] CFGDSN_delay;
  wire [63:0] CFGINTERRUPTMSIXADDRESS_delay;
  wire [7:0] CFGDSBUSNUMBER_delay;
  wire [7:0] CFGDSPORTNUMBER_delay;
  wire [7:0] CFGREVID_delay;
  wire [7:0] CFGVFFLRDONE_delay;
  wire [7:0] SAXISCCTKEEP_delay;
  wire [7:0] SAXISRQTKEEP_delay;
  wire [8:0] CFGINTERRUPTMSITPHSTTAG_delay;
  wire [9:0] DRPADDR_delay;

  
  assign #(out_delay) CFGCURRENTSPEED = CFGCURRENTSPEED_delay;
  assign #(out_delay) CFGDPASUBSTATECHANGE = CFGDPASUBSTATECHANGE_delay;
  assign #(out_delay) CFGERRCOROUT = CFGERRCOROUT_delay;
  assign #(out_delay) CFGERRFATALOUT = CFGERRFATALOUT_delay;
  assign #(out_delay) CFGERRNONFATALOUT = CFGERRNONFATALOUT_delay;
  assign #(out_delay) CFGEXTFUNCTIONNUMBER = CFGEXTFUNCTIONNUMBER_delay;
  assign #(out_delay) CFGEXTREADRECEIVED = CFGEXTREADRECEIVED_delay;
  assign #(out_delay) CFGEXTREGISTERNUMBER = CFGEXTREGISTERNUMBER_delay;
  assign #(out_delay) CFGEXTWRITEBYTEENABLE = CFGEXTWRITEBYTEENABLE_delay;
  assign #(out_delay) CFGEXTWRITEDATA = CFGEXTWRITEDATA_delay;
  assign #(out_delay) CFGEXTWRITERECEIVED = CFGEXTWRITERECEIVED_delay;
  assign #(out_delay) CFGFCCPLD = CFGFCCPLD_delay;
  assign #(out_delay) CFGFCCPLH = CFGFCCPLH_delay;
  assign #(out_delay) CFGFCNPD = CFGFCNPD_delay;
  assign #(out_delay) CFGFCNPH = CFGFCNPH_delay;
  assign #(out_delay) CFGFCPD = CFGFCPD_delay;
  assign #(out_delay) CFGFCPH = CFGFCPH_delay;
  assign #(out_delay) CFGFLRINPROCESS = CFGFLRINPROCESS_delay;
  assign #(out_delay) CFGFUNCTIONPOWERSTATE = CFGFUNCTIONPOWERSTATE_delay;
  assign #(out_delay) CFGFUNCTIONSTATUS = CFGFUNCTIONSTATUS_delay;
  assign #(out_delay) CFGHOTRESETOUT = CFGHOTRESETOUT_delay;
  assign #(out_delay) CFGINTERRUPTMSIDATA = CFGINTERRUPTMSIDATA_delay;
  assign #(out_delay) CFGINTERRUPTMSIENABLE = CFGINTERRUPTMSIENABLE_delay;
  assign #(out_delay) CFGINTERRUPTMSIFAIL = CFGINTERRUPTMSIFAIL_delay;
  assign #(out_delay) CFGINTERRUPTMSIMASKUPDATE = CFGINTERRUPTMSIMASKUPDATE_delay;
  assign #(out_delay) CFGINTERRUPTMSIMMENABLE = CFGINTERRUPTMSIMMENABLE_delay;
  assign #(out_delay) CFGINTERRUPTMSISENT = CFGINTERRUPTMSISENT_delay;
  assign #(out_delay) CFGINTERRUPTMSIVFENABLE = CFGINTERRUPTMSIVFENABLE_delay;
  assign #(out_delay) CFGINTERRUPTMSIXENABLE = CFGINTERRUPTMSIXENABLE_delay;
  assign #(out_delay) CFGINTERRUPTMSIXFAIL = CFGINTERRUPTMSIXFAIL_delay;
  assign #(out_delay) CFGINTERRUPTMSIXMASK = CFGINTERRUPTMSIXMASK_delay;
  assign #(out_delay) CFGINTERRUPTMSIXSENT = CFGINTERRUPTMSIXSENT_delay;
  assign #(out_delay) CFGINTERRUPTMSIXVFENABLE = CFGINTERRUPTMSIXVFENABLE_delay;
  assign #(out_delay) CFGINTERRUPTMSIXVFMASK = CFGINTERRUPTMSIXVFMASK_delay;
  assign #(out_delay) CFGINTERRUPTSENT = CFGINTERRUPTSENT_delay;
  assign #(out_delay) CFGLINKPOWERSTATE = CFGLINKPOWERSTATE_delay;
  assign #(out_delay) CFGLOCALERROR = CFGLOCALERROR_delay;
  assign #(out_delay) CFGLTRENABLE = CFGLTRENABLE_delay;
  assign #(out_delay) CFGLTSSMSTATE = CFGLTSSMSTATE_delay;
  assign #(out_delay) CFGMAXPAYLOAD = CFGMAXPAYLOAD_delay;
  assign #(out_delay) CFGMAXREADREQ = CFGMAXREADREQ_delay;
  assign #(out_delay) CFGMGMTREADDATA = CFGMGMTREADDATA_delay;
  assign #(out_delay) CFGMGMTREADWRITEDONE = CFGMGMTREADWRITEDONE_delay;
  assign #(out_delay) CFGMSGRECEIVED = CFGMSGRECEIVED_delay;
  assign #(out_delay) CFGMSGRECEIVEDDATA = CFGMSGRECEIVEDDATA_delay;
  assign #(out_delay) CFGMSGRECEIVEDTYPE = CFGMSGRECEIVEDTYPE_delay;
  assign #(out_delay) CFGMSGTRANSMITDONE = CFGMSGTRANSMITDONE_delay;
  assign #(out_delay) CFGNEGOTIATEDWIDTH = CFGNEGOTIATEDWIDTH_delay;
  assign #(out_delay) CFGOBFFENABLE = CFGOBFFENABLE_delay;
  assign #(out_delay) CFGPERFUNCSTATUSDATA = CFGPERFUNCSTATUSDATA_delay;
  assign #(out_delay) CFGPERFUNCTIONUPDATEDONE = CFGPERFUNCTIONUPDATEDONE_delay;
  assign #(out_delay) CFGPHYLINKDOWN = CFGPHYLINKDOWN_delay;
  assign #(out_delay) CFGPHYLINKSTATUS = CFGPHYLINKSTATUS_delay;
  assign #(out_delay) CFGPLSTATUSCHANGE = CFGPLSTATUSCHANGE_delay;
  assign #(out_delay) CFGPOWERSTATECHANGEINTERRUPT = CFGPOWERSTATECHANGEINTERRUPT_delay;
  assign #(out_delay) CFGRCBSTATUS = CFGRCBSTATUS_delay;
  assign #(out_delay) CFGTPHFUNCTIONNUM = CFGTPHFUNCTIONNUM_delay;
  assign #(out_delay) CFGTPHREQUESTERENABLE = CFGTPHREQUESTERENABLE_delay;
  assign #(out_delay) CFGTPHSTMODE = CFGTPHSTMODE_delay;
  assign #(out_delay) CFGTPHSTTADDRESS = CFGTPHSTTADDRESS_delay;
  assign #(out_delay) CFGTPHSTTREADENABLE = CFGTPHSTTREADENABLE_delay;
  assign #(out_delay) CFGTPHSTTWRITEBYTEVALID = CFGTPHSTTWRITEBYTEVALID_delay;
  assign #(out_delay) CFGTPHSTTWRITEDATA = CFGTPHSTTWRITEDATA_delay;
  assign #(out_delay) CFGTPHSTTWRITEENABLE = CFGTPHSTTWRITEENABLE_delay;
  assign #(out_delay) CFGVFFLRINPROCESS = CFGVFFLRINPROCESS_delay;
  assign #(out_delay) CFGVFPOWERSTATE = CFGVFPOWERSTATE_delay;
  assign #(out_delay) CFGVFSTATUS = CFGVFSTATUS_delay;
  assign #(out_delay) CFGVFTPHREQUESTERENABLE = CFGVFTPHREQUESTERENABLE_delay;
  assign #(out_delay) CFGVFTPHSTMODE = CFGVFTPHSTMODE_delay;
  assign #(out_delay) CONFMCAPDESIGNSWITCH = CONFMCAPDESIGNSWITCH_delay;
  assign #(out_delay) CONFMCAPEOS = CONFMCAPEOS_delay;
  assign #(out_delay) CONFMCAPINUSEBYPCIE = CONFMCAPINUSEBYPCIE_delay;
  assign #(out_delay) CONFREQREADY = CONFREQREADY_delay;
  assign #(out_delay) CONFRESPRDATA = CONFRESPRDATA_delay;
  assign #(out_delay) CONFRESPVALID = CONFRESPVALID_delay;
  assign #(out_delay) DBGDATAOUT = DBGDATAOUT_delay;
  assign #(out_delay) DBGMCAPCSB = DBGMCAPCSB_delay;
  assign #(out_delay) DBGMCAPDATA = DBGMCAPDATA_delay;
  assign #(out_delay) DBGMCAPEOS = DBGMCAPEOS_delay;
  assign #(out_delay) DBGMCAPERROR = DBGMCAPERROR_delay;
  assign #(out_delay) DBGMCAPMODE = DBGMCAPMODE_delay;
  assign #(out_delay) DBGMCAPRDATAVALID = DBGMCAPRDATAVALID_delay;
  assign #(out_delay) DBGMCAPRDWRB = DBGMCAPRDWRB_delay;
  assign #(out_delay) DBGMCAPRESET = DBGMCAPRESET_delay;
  assign #(out_delay) DBGPLDATABLOCKRECEIVEDAFTEREDS = DBGPLDATABLOCKRECEIVEDAFTEREDS_delay;
  assign #(out_delay) DBGPLGEN3FRAMINGERRORDETECTED = DBGPLGEN3FRAMINGERRORDETECTED_delay;
  assign #(out_delay) DBGPLGEN3SYNCHEADERERRORDETECTED = DBGPLGEN3SYNCHEADERERRORDETECTED_delay;
  assign #(out_delay) DBGPLINFERREDRXELECTRICALIDLE = DBGPLINFERREDRXELECTRICALIDLE_delay;
  assign #(out_delay) DRPDO = DRPDO_delay;
  assign #(out_delay) DRPRDY = DRPRDY_delay;
  assign #(out_delay) LL2LMMASTERTLPSENT0 = LL2LMMASTERTLPSENT0_delay;
  assign #(out_delay) LL2LMMASTERTLPSENT1 = LL2LMMASTERTLPSENT1_delay;
  assign #(out_delay) LL2LMMASTERTLPSENTTLPID0 = LL2LMMASTERTLPSENTTLPID0_delay;
  assign #(out_delay) LL2LMMASTERTLPSENTTLPID1 = LL2LMMASTERTLPSENTTLPID1_delay;
  assign #(out_delay) LL2LMMAXISRXTDATA = LL2LMMAXISRXTDATA_delay;
  assign #(out_delay) LL2LMMAXISRXTUSER = LL2LMMAXISRXTUSER_delay;
  assign #(out_delay) LL2LMMAXISRXTVALID = LL2LMMAXISRXTVALID_delay;
  assign #(out_delay) LL2LMSAXISTXTREADY = LL2LMSAXISTXTREADY_delay;
  assign #(out_delay) MAXISCQTDATA = MAXISCQTDATA_delay;
  assign #(out_delay) MAXISCQTKEEP = MAXISCQTKEEP_delay;
  assign #(out_delay) MAXISCQTLAST = MAXISCQTLAST_delay;
  assign #(out_delay) MAXISCQTUSER = MAXISCQTUSER_delay;
  assign #(out_delay) MAXISCQTVALID = MAXISCQTVALID_delay;
  assign #(out_delay) MAXISRCTDATA = MAXISRCTDATA_delay;
  assign #(out_delay) MAXISRCTKEEP = MAXISRCTKEEP_delay;
  assign #(out_delay) MAXISRCTLAST = MAXISRCTLAST_delay;
  assign #(out_delay) MAXISRCTUSER = MAXISRCTUSER_delay;
  assign #(out_delay) MAXISRCTVALID = MAXISRCTVALID_delay;
  assign #(out_delay) MICOMPLETIONRAMREADADDRESSAL = MICOMPLETIONRAMREADADDRESSAL_delay;
  assign #(out_delay) MICOMPLETIONRAMREADADDRESSAU = MICOMPLETIONRAMREADADDRESSAU_delay;
  assign #(out_delay) MICOMPLETIONRAMREADADDRESSBL = MICOMPLETIONRAMREADADDRESSBL_delay;
  assign #(out_delay) MICOMPLETIONRAMREADADDRESSBU = MICOMPLETIONRAMREADADDRESSBU_delay;
  assign #(out_delay) MICOMPLETIONRAMREADENABLEL = MICOMPLETIONRAMREADENABLEL_delay;
  assign #(out_delay) MICOMPLETIONRAMREADENABLEU = MICOMPLETIONRAMREADENABLEU_delay;
  assign #(out_delay) MICOMPLETIONRAMWRITEADDRESSAL = MICOMPLETIONRAMWRITEADDRESSAL_delay;
  assign #(out_delay) MICOMPLETIONRAMWRITEADDRESSAU = MICOMPLETIONRAMWRITEADDRESSAU_delay;
  assign #(out_delay) MICOMPLETIONRAMWRITEADDRESSBL = MICOMPLETIONRAMWRITEADDRESSBL_delay;
  assign #(out_delay) MICOMPLETIONRAMWRITEADDRESSBU = MICOMPLETIONRAMWRITEADDRESSBU_delay;
  assign #(out_delay) MICOMPLETIONRAMWRITEDATAL = MICOMPLETIONRAMWRITEDATAL_delay;
  assign #(out_delay) MICOMPLETIONRAMWRITEDATAU = MICOMPLETIONRAMWRITEDATAU_delay;
  assign #(out_delay) MICOMPLETIONRAMWRITEENABLEL = MICOMPLETIONRAMWRITEENABLEL_delay;
  assign #(out_delay) MICOMPLETIONRAMWRITEENABLEU = MICOMPLETIONRAMWRITEENABLEU_delay;
  assign #(out_delay) MIREPLAYRAMADDRESS = MIREPLAYRAMADDRESS_delay;
  assign #(out_delay) MIREPLAYRAMREADENABLE = MIREPLAYRAMREADENABLE_delay;
  assign #(out_delay) MIREPLAYRAMWRITEDATA = MIREPLAYRAMWRITEDATA_delay;
  assign #(out_delay) MIREPLAYRAMWRITEENABLE = MIREPLAYRAMWRITEENABLE_delay;
  assign #(out_delay) MIREQUESTRAMREADADDRESSA = MIREQUESTRAMREADADDRESSA_delay;
  assign #(out_delay) MIREQUESTRAMREADADDRESSB = MIREQUESTRAMREADADDRESSB_delay;
  assign #(out_delay) MIREQUESTRAMREADENABLE = MIREQUESTRAMREADENABLE_delay;
  assign #(out_delay) MIREQUESTRAMWRITEADDRESSA = MIREQUESTRAMWRITEADDRESSA_delay;
  assign #(out_delay) MIREQUESTRAMWRITEADDRESSB = MIREQUESTRAMWRITEADDRESSB_delay;
  assign #(out_delay) MIREQUESTRAMWRITEDATA = MIREQUESTRAMWRITEDATA_delay;
  assign #(out_delay) MIREQUESTRAMWRITEENABLE = MIREQUESTRAMWRITEENABLE_delay;
  assign #(out_delay) PCIECQNPREQCOUNT = PCIECQNPREQCOUNT_delay;
  assign #(out_delay) PCIEPERST0B = PCIEPERST0B_delay;
  assign #(out_delay) PCIEPERST1B = PCIEPERST1B_delay;
  assign #(out_delay) PCIERQSEQNUM = PCIERQSEQNUM_delay;
  assign #(out_delay) PCIERQSEQNUMVLD = PCIERQSEQNUMVLD_delay;
  assign #(out_delay) PCIERQTAG = PCIERQTAG_delay;
  assign #(out_delay) PCIERQTAGAV = PCIERQTAGAV_delay;
  assign #(out_delay) PCIERQTAGVLD = PCIERQTAGVLD_delay;
  assign #(out_delay) PCIETFCNPDAV = PCIETFCNPDAV_delay;
  assign #(out_delay) PCIETFCNPHAV = PCIETFCNPHAV_delay;
  assign #(out_delay) PIPERX0EQCONTROL = PIPERX0EQCONTROL_delay;
  assign #(out_delay) PIPERX0EQLPLFFS = PIPERX0EQLPLFFS_delay;
  assign #(out_delay) PIPERX0EQLPTXPRESET = PIPERX0EQLPTXPRESET_delay;
  assign #(out_delay) PIPERX0EQPRESET = PIPERX0EQPRESET_delay;
  assign #(out_delay) PIPERX0POLARITY = PIPERX0POLARITY_delay;
  assign #(out_delay) PIPERX1EQCONTROL = PIPERX1EQCONTROL_delay;
  assign #(out_delay) PIPERX1EQLPLFFS = PIPERX1EQLPLFFS_delay;
  assign #(out_delay) PIPERX1EQLPTXPRESET = PIPERX1EQLPTXPRESET_delay;
  assign #(out_delay) PIPERX1EQPRESET = PIPERX1EQPRESET_delay;
  assign #(out_delay) PIPERX1POLARITY = PIPERX1POLARITY_delay;
  assign #(out_delay) PIPERX2EQCONTROL = PIPERX2EQCONTROL_delay;
  assign #(out_delay) PIPERX2EQLPLFFS = PIPERX2EQLPLFFS_delay;
  assign #(out_delay) PIPERX2EQLPTXPRESET = PIPERX2EQLPTXPRESET_delay;
  assign #(out_delay) PIPERX2EQPRESET = PIPERX2EQPRESET_delay;
  assign #(out_delay) PIPERX2POLARITY = PIPERX2POLARITY_delay;
  assign #(out_delay) PIPERX3EQCONTROL = PIPERX3EQCONTROL_delay;
  assign #(out_delay) PIPERX3EQLPLFFS = PIPERX3EQLPLFFS_delay;
  assign #(out_delay) PIPERX3EQLPTXPRESET = PIPERX3EQLPTXPRESET_delay;
  assign #(out_delay) PIPERX3EQPRESET = PIPERX3EQPRESET_delay;
  assign #(out_delay) PIPERX3POLARITY = PIPERX3POLARITY_delay;
  assign #(out_delay) PIPERX4EQCONTROL = PIPERX4EQCONTROL_delay;
  assign #(out_delay) PIPERX4EQLPLFFS = PIPERX4EQLPLFFS_delay;
  assign #(out_delay) PIPERX4EQLPTXPRESET = PIPERX4EQLPTXPRESET_delay;
  assign #(out_delay) PIPERX4EQPRESET = PIPERX4EQPRESET_delay;
  assign #(out_delay) PIPERX4POLARITY = PIPERX4POLARITY_delay;
  assign #(out_delay) PIPERX5EQCONTROL = PIPERX5EQCONTROL_delay;
  assign #(out_delay) PIPERX5EQLPLFFS = PIPERX5EQLPLFFS_delay;
  assign #(out_delay) PIPERX5EQLPTXPRESET = PIPERX5EQLPTXPRESET_delay;
  assign #(out_delay) PIPERX5EQPRESET = PIPERX5EQPRESET_delay;
  assign #(out_delay) PIPERX5POLARITY = PIPERX5POLARITY_delay;
  assign #(out_delay) PIPERX6EQCONTROL = PIPERX6EQCONTROL_delay;
  assign #(out_delay) PIPERX6EQLPLFFS = PIPERX6EQLPLFFS_delay;
  assign #(out_delay) PIPERX6EQLPTXPRESET = PIPERX6EQLPTXPRESET_delay;
  assign #(out_delay) PIPERX6EQPRESET = PIPERX6EQPRESET_delay;
  assign #(out_delay) PIPERX6POLARITY = PIPERX6POLARITY_delay;
  assign #(out_delay) PIPERX7EQCONTROL = PIPERX7EQCONTROL_delay;
  assign #(out_delay) PIPERX7EQLPLFFS = PIPERX7EQLPLFFS_delay;
  assign #(out_delay) PIPERX7EQLPTXPRESET = PIPERX7EQLPTXPRESET_delay;
  assign #(out_delay) PIPERX7EQPRESET = PIPERX7EQPRESET_delay;
  assign #(out_delay) PIPERX7POLARITY = PIPERX7POLARITY_delay;
  assign #(out_delay) PIPETX0CHARISK = PIPETX0CHARISK_delay;
  assign #(out_delay) PIPETX0COMPLIANCE = PIPETX0COMPLIANCE_delay;
  assign #(out_delay) PIPETX0DATA = PIPETX0DATA_delay;
  assign #(out_delay) PIPETX0DATAVALID = PIPETX0DATAVALID_delay;
  assign #(out_delay) PIPETX0DEEMPH = PIPETX0DEEMPH_delay;
  assign #(out_delay) PIPETX0ELECIDLE = PIPETX0ELECIDLE_delay;
  assign #(out_delay) PIPETX0EQCONTROL = PIPETX0EQCONTROL_delay;
  assign #(out_delay) PIPETX0EQDEEMPH = PIPETX0EQDEEMPH_delay;
  assign #(out_delay) PIPETX0EQPRESET = PIPETX0EQPRESET_delay;
  assign #(out_delay) PIPETX0MARGIN = PIPETX0MARGIN_delay;
  assign #(out_delay) PIPETX0POWERDOWN = PIPETX0POWERDOWN_delay;
  assign #(out_delay) PIPETX0RATE = PIPETX0RATE_delay;
  assign #(out_delay) PIPETX0RCVRDET = PIPETX0RCVRDET_delay;
  assign #(out_delay) PIPETX0RESET = PIPETX0RESET_delay;
  assign #(out_delay) PIPETX0STARTBLOCK = PIPETX0STARTBLOCK_delay;
  assign #(out_delay) PIPETX0SWING = PIPETX0SWING_delay;
  assign #(out_delay) PIPETX0SYNCHEADER = PIPETX0SYNCHEADER_delay;
  assign #(out_delay) PIPETX1CHARISK = PIPETX1CHARISK_delay;
  assign #(out_delay) PIPETX1COMPLIANCE = PIPETX1COMPLIANCE_delay;
  assign #(out_delay) PIPETX1DATA = PIPETX1DATA_delay;
  assign #(out_delay) PIPETX1DATAVALID = PIPETX1DATAVALID_delay;
  assign #(out_delay) PIPETX1DEEMPH = PIPETX1DEEMPH_delay;
  assign #(out_delay) PIPETX1ELECIDLE = PIPETX1ELECIDLE_delay;
  assign #(out_delay) PIPETX1EQCONTROL = PIPETX1EQCONTROL_delay;
  assign #(out_delay) PIPETX1EQDEEMPH = PIPETX1EQDEEMPH_delay;
  assign #(out_delay) PIPETX1EQPRESET = PIPETX1EQPRESET_delay;
  assign #(out_delay) PIPETX1MARGIN = PIPETX1MARGIN_delay;
  assign #(out_delay) PIPETX1POWERDOWN = PIPETX1POWERDOWN_delay;
  assign #(out_delay) PIPETX1RATE = PIPETX1RATE_delay;
  assign #(out_delay) PIPETX1RCVRDET = PIPETX1RCVRDET_delay;
  assign #(out_delay) PIPETX1RESET = PIPETX1RESET_delay;
  assign #(out_delay) PIPETX1STARTBLOCK = PIPETX1STARTBLOCK_delay;
  assign #(out_delay) PIPETX1SWING = PIPETX1SWING_delay;
  assign #(out_delay) PIPETX1SYNCHEADER = PIPETX1SYNCHEADER_delay;
  assign #(out_delay) PIPETX2CHARISK = PIPETX2CHARISK_delay;
  assign #(out_delay) PIPETX2COMPLIANCE = PIPETX2COMPLIANCE_delay;
  assign #(out_delay) PIPETX2DATA = PIPETX2DATA_delay;
  assign #(out_delay) PIPETX2DATAVALID = PIPETX2DATAVALID_delay;
  assign #(out_delay) PIPETX2DEEMPH = PIPETX2DEEMPH_delay;
  assign #(out_delay) PIPETX2ELECIDLE = PIPETX2ELECIDLE_delay;
  assign #(out_delay) PIPETX2EQCONTROL = PIPETX2EQCONTROL_delay;
  assign #(out_delay) PIPETX2EQDEEMPH = PIPETX2EQDEEMPH_delay;
  assign #(out_delay) PIPETX2EQPRESET = PIPETX2EQPRESET_delay;
  assign #(out_delay) PIPETX2MARGIN = PIPETX2MARGIN_delay;
  assign #(out_delay) PIPETX2POWERDOWN = PIPETX2POWERDOWN_delay;
  assign #(out_delay) PIPETX2RATE = PIPETX2RATE_delay;
  assign #(out_delay) PIPETX2RCVRDET = PIPETX2RCVRDET_delay;
  assign #(out_delay) PIPETX2RESET = PIPETX2RESET_delay;
  assign #(out_delay) PIPETX2STARTBLOCK = PIPETX2STARTBLOCK_delay;
  assign #(out_delay) PIPETX2SWING = PIPETX2SWING_delay;
  assign #(out_delay) PIPETX2SYNCHEADER = PIPETX2SYNCHEADER_delay;
  assign #(out_delay) PIPETX3CHARISK = PIPETX3CHARISK_delay;
  assign #(out_delay) PIPETX3COMPLIANCE = PIPETX3COMPLIANCE_delay;
  assign #(out_delay) PIPETX3DATA = PIPETX3DATA_delay;
  assign #(out_delay) PIPETX3DATAVALID = PIPETX3DATAVALID_delay;
  assign #(out_delay) PIPETX3DEEMPH = PIPETX3DEEMPH_delay;
  assign #(out_delay) PIPETX3ELECIDLE = PIPETX3ELECIDLE_delay;
  assign #(out_delay) PIPETX3EQCONTROL = PIPETX3EQCONTROL_delay;
  assign #(out_delay) PIPETX3EQDEEMPH = PIPETX3EQDEEMPH_delay;
  assign #(out_delay) PIPETX3EQPRESET = PIPETX3EQPRESET_delay;
  assign #(out_delay) PIPETX3MARGIN = PIPETX3MARGIN_delay;
  assign #(out_delay) PIPETX3POWERDOWN = PIPETX3POWERDOWN_delay;
  assign #(out_delay) PIPETX3RATE = PIPETX3RATE_delay;
  assign #(out_delay) PIPETX3RCVRDET = PIPETX3RCVRDET_delay;
  assign #(out_delay) PIPETX3RESET = PIPETX3RESET_delay;
  assign #(out_delay) PIPETX3STARTBLOCK = PIPETX3STARTBLOCK_delay;
  assign #(out_delay) PIPETX3SWING = PIPETX3SWING_delay;
  assign #(out_delay) PIPETX3SYNCHEADER = PIPETX3SYNCHEADER_delay;
  assign #(out_delay) PIPETX4CHARISK = PIPETX4CHARISK_delay;
  assign #(out_delay) PIPETX4COMPLIANCE = PIPETX4COMPLIANCE_delay;
  assign #(out_delay) PIPETX4DATA = PIPETX4DATA_delay;
  assign #(out_delay) PIPETX4DATAVALID = PIPETX4DATAVALID_delay;
  assign #(out_delay) PIPETX4DEEMPH = PIPETX4DEEMPH_delay;
  assign #(out_delay) PIPETX4ELECIDLE = PIPETX4ELECIDLE_delay;
  assign #(out_delay) PIPETX4EQCONTROL = PIPETX4EQCONTROL_delay;
  assign #(out_delay) PIPETX4EQDEEMPH = PIPETX4EQDEEMPH_delay;
  assign #(out_delay) PIPETX4EQPRESET = PIPETX4EQPRESET_delay;
  assign #(out_delay) PIPETX4MARGIN = PIPETX4MARGIN_delay;
  assign #(out_delay) PIPETX4POWERDOWN = PIPETX4POWERDOWN_delay;
  assign #(out_delay) PIPETX4RATE = PIPETX4RATE_delay;
  assign #(out_delay) PIPETX4RCVRDET = PIPETX4RCVRDET_delay;
  assign #(out_delay) PIPETX4RESET = PIPETX4RESET_delay;
  assign #(out_delay) PIPETX4STARTBLOCK = PIPETX4STARTBLOCK_delay;
  assign #(out_delay) PIPETX4SWING = PIPETX4SWING_delay;
  assign #(out_delay) PIPETX4SYNCHEADER = PIPETX4SYNCHEADER_delay;
  assign #(out_delay) PIPETX5CHARISK = PIPETX5CHARISK_delay;
  assign #(out_delay) PIPETX5COMPLIANCE = PIPETX5COMPLIANCE_delay;
  assign #(out_delay) PIPETX5DATA = PIPETX5DATA_delay;
  assign #(out_delay) PIPETX5DATAVALID = PIPETX5DATAVALID_delay;
  assign #(out_delay) PIPETX5DEEMPH = PIPETX5DEEMPH_delay;
  assign #(out_delay) PIPETX5ELECIDLE = PIPETX5ELECIDLE_delay;
  assign #(out_delay) PIPETX5EQCONTROL = PIPETX5EQCONTROL_delay;
  assign #(out_delay) PIPETX5EQDEEMPH = PIPETX5EQDEEMPH_delay;
  assign #(out_delay) PIPETX5EQPRESET = PIPETX5EQPRESET_delay;
  assign #(out_delay) PIPETX5MARGIN = PIPETX5MARGIN_delay;
  assign #(out_delay) PIPETX5POWERDOWN = PIPETX5POWERDOWN_delay;
  assign #(out_delay) PIPETX5RATE = PIPETX5RATE_delay;
  assign #(out_delay) PIPETX5RCVRDET = PIPETX5RCVRDET_delay;
  assign #(out_delay) PIPETX5RESET = PIPETX5RESET_delay;
  assign #(out_delay) PIPETX5STARTBLOCK = PIPETX5STARTBLOCK_delay;
  assign #(out_delay) PIPETX5SWING = PIPETX5SWING_delay;
  assign #(out_delay) PIPETX5SYNCHEADER = PIPETX5SYNCHEADER_delay;
  assign #(out_delay) PIPETX6CHARISK = PIPETX6CHARISK_delay;
  assign #(out_delay) PIPETX6COMPLIANCE = PIPETX6COMPLIANCE_delay;
  assign #(out_delay) PIPETX6DATA = PIPETX6DATA_delay;
  assign #(out_delay) PIPETX6DATAVALID = PIPETX6DATAVALID_delay;
  assign #(out_delay) PIPETX6DEEMPH = PIPETX6DEEMPH_delay;
  assign #(out_delay) PIPETX6ELECIDLE = PIPETX6ELECIDLE_delay;
  assign #(out_delay) PIPETX6EQCONTROL = PIPETX6EQCONTROL_delay;
  assign #(out_delay) PIPETX6EQDEEMPH = PIPETX6EQDEEMPH_delay;
  assign #(out_delay) PIPETX6EQPRESET = PIPETX6EQPRESET_delay;
  assign #(out_delay) PIPETX6MARGIN = PIPETX6MARGIN_delay;
  assign #(out_delay) PIPETX6POWERDOWN = PIPETX6POWERDOWN_delay;
  assign #(out_delay) PIPETX6RATE = PIPETX6RATE_delay;
  assign #(out_delay) PIPETX6RCVRDET = PIPETX6RCVRDET_delay;
  assign #(out_delay) PIPETX6RESET = PIPETX6RESET_delay;
  assign #(out_delay) PIPETX6STARTBLOCK = PIPETX6STARTBLOCK_delay;
  assign #(out_delay) PIPETX6SWING = PIPETX6SWING_delay;
  assign #(out_delay) PIPETX6SYNCHEADER = PIPETX6SYNCHEADER_delay;
  assign #(out_delay) PIPETX7CHARISK = PIPETX7CHARISK_delay;
  assign #(out_delay) PIPETX7COMPLIANCE = PIPETX7COMPLIANCE_delay;
  assign #(out_delay) PIPETX7DATA = PIPETX7DATA_delay;
  assign #(out_delay) PIPETX7DATAVALID = PIPETX7DATAVALID_delay;
  assign #(out_delay) PIPETX7DEEMPH = PIPETX7DEEMPH_delay;
  assign #(out_delay) PIPETX7ELECIDLE = PIPETX7ELECIDLE_delay;
  assign #(out_delay) PIPETX7EQCONTROL = PIPETX7EQCONTROL_delay;
  assign #(out_delay) PIPETX7EQDEEMPH = PIPETX7EQDEEMPH_delay;
  assign #(out_delay) PIPETX7EQPRESET = PIPETX7EQPRESET_delay;
  assign #(out_delay) PIPETX7MARGIN = PIPETX7MARGIN_delay;
  assign #(out_delay) PIPETX7POWERDOWN = PIPETX7POWERDOWN_delay;
  assign #(out_delay) PIPETX7RATE = PIPETX7RATE_delay;
  assign #(out_delay) PIPETX7RCVRDET = PIPETX7RCVRDET_delay;
  assign #(out_delay) PIPETX7RESET = PIPETX7RESET_delay;
  assign #(out_delay) PIPETX7STARTBLOCK = PIPETX7STARTBLOCK_delay;
  assign #(out_delay) PIPETX7SWING = PIPETX7SWING_delay;
  assign #(out_delay) PIPETX7SYNCHEADER = PIPETX7SYNCHEADER_delay;
  assign #(out_delay) PLEQINPROGRESS = PLEQINPROGRESS_delay;
  assign #(out_delay) PLEQPHASE = PLEQPHASE_delay;
  assign #(out_delay) SAXISCCTREADY = SAXISCCTREADY_delay;
  assign #(out_delay) SAXISRQTREADY = SAXISRQTREADY_delay;
  assign #(out_delay) SPAREOUT = SPAREOUT_delay;
  
`ifndef XIL_TIMING // inputs with timing checks
  assign #(inclk_delay) CORECLKMICOMPLETIONRAML_delay = CORECLKMICOMPLETIONRAML;
  assign #(inclk_delay) CORECLKMICOMPLETIONRAMU_delay = CORECLKMICOMPLETIONRAMU;
  assign #(inclk_delay) CORECLKMIREPLAYRAM_delay = CORECLKMIREPLAYRAM;
  assign #(inclk_delay) CORECLKMIREQUESTRAM_delay = CORECLKMIREQUESTRAM;
  assign #(inclk_delay) CORECLK_delay = CORECLK;
  assign #(inclk_delay) DRPCLK_delay = DRPCLK;
  assign #(inclk_delay) MCAPCLK_delay = MCAPCLK;
  assign #(inclk_delay) PIPECLK_delay = PIPECLK;
  assign #(inclk_delay) USERCLK_delay = USERCLK;

  assign #(in_delay) CFGCONFIGSPACEENABLE_delay = CFGCONFIGSPACEENABLE;
  assign #(in_delay) CFGERRCORIN_delay = CFGERRCORIN;
  assign #(in_delay) CFGERRUNCORIN_delay = CFGERRUNCORIN;
  assign #(in_delay) CFGEXTREADDATAVALID_delay = CFGEXTREADDATAVALID;
  assign #(in_delay) CFGHOTRESETIN_delay = CFGHOTRESETIN;
  assign #(in_delay) CFGINTERRUPTMSIPENDINGSTATUSDATAENABLE_delay = CFGINTERRUPTMSIPENDINGSTATUSDATAENABLE;
  assign #(in_delay) CFGINTERRUPTMSITPHPRESENT_delay = CFGINTERRUPTMSITPHPRESENT;
  assign #(in_delay) CFGINTERRUPTMSIXINT_delay = CFGINTERRUPTMSIXINT;
  assign #(in_delay) CFGLINKTRAININGENABLE_delay = CFGLINKTRAININGENABLE;
  assign #(in_delay) CFGMGMTREAD_delay = CFGMGMTREAD;
  assign #(in_delay) CFGMGMTTYPE1CFGREGACCESS_delay = CFGMGMTTYPE1CFGREGACCESS;
  assign #(in_delay) CFGMGMTWRITE_delay = CFGMGMTWRITE;
  assign #(in_delay) CFGMSGTRANSMIT_delay = CFGMSGTRANSMIT;
  assign #(in_delay) CFGPERFUNCTIONOUTPUTREQUEST_delay = CFGPERFUNCTIONOUTPUTREQUEST;
  assign #(in_delay) CFGPOWERSTATECHANGEACK_delay = CFGPOWERSTATECHANGEACK;
  assign #(in_delay) CFGREQPMTRANSITIONL23READY_delay = CFGREQPMTRANSITIONL23READY;
  assign #(in_delay) CFGTPHSTTREADDATAVALID_delay = CFGTPHSTTREADDATAVALID;
  assign #(in_delay) CONFMCAPREQUESTBYCONF_delay = CONFMCAPREQUESTBYCONF;
  assign #(in_delay) CONFREQVALID_delay = CONFREQVALID;
  assign #(in_delay) DBGCFGLOCALMGMTREGOVERRIDE_delay = DBGCFGLOCALMGMTREGOVERRIDE;
  assign #(in_delay) DRPEN_delay = DRPEN;
  assign #(in_delay) DRPWE_delay = DRPWE;
  assign #(in_delay) LL2LMSAXISTXTVALID_delay = LL2LMSAXISTXTVALID;
  assign #(in_delay) PCIECQNPREQ_delay = PCIECQNPREQ;
  assign #(in_delay) PIPERX0DATAVALID_delay = PIPERX0DATAVALID;
  assign #(in_delay) PIPERX0ELECIDLE_delay = PIPERX0ELECIDLE;
  assign #(in_delay) PIPERX0EQDONE_delay = PIPERX0EQDONE;
  assign #(in_delay) PIPERX0EQLPADAPTDONE_delay = PIPERX0EQLPADAPTDONE;
  assign #(in_delay) PIPERX0EQLPLFFSSEL_delay = PIPERX0EQLPLFFSSEL;
  assign #(in_delay) PIPERX0PHYSTATUS_delay = PIPERX0PHYSTATUS;
  assign #(in_delay) PIPERX0STARTBLOCK_delay = PIPERX0STARTBLOCK;
  assign #(in_delay) PIPERX0VALID_delay = PIPERX0VALID;
  assign #(in_delay) PIPERX1DATAVALID_delay = PIPERX1DATAVALID;
  assign #(in_delay) PIPERX1ELECIDLE_delay = PIPERX1ELECIDLE;
  assign #(in_delay) PIPERX1EQDONE_delay = PIPERX1EQDONE;
  assign #(in_delay) PIPERX1EQLPADAPTDONE_delay = PIPERX1EQLPADAPTDONE;
  assign #(in_delay) PIPERX1EQLPLFFSSEL_delay = PIPERX1EQLPLFFSSEL;
  assign #(in_delay) PIPERX1PHYSTATUS_delay = PIPERX1PHYSTATUS;
  assign #(in_delay) PIPERX1STARTBLOCK_delay = PIPERX1STARTBLOCK;
  assign #(in_delay) PIPERX1VALID_delay = PIPERX1VALID;
  assign #(in_delay) PIPERX2DATAVALID_delay = PIPERX2DATAVALID;
  assign #(in_delay) PIPERX2ELECIDLE_delay = PIPERX2ELECIDLE;
  assign #(in_delay) PIPERX2EQDONE_delay = PIPERX2EQDONE;
  assign #(in_delay) PIPERX2EQLPADAPTDONE_delay = PIPERX2EQLPADAPTDONE;
  assign #(in_delay) PIPERX2EQLPLFFSSEL_delay = PIPERX2EQLPLFFSSEL;
  assign #(in_delay) PIPERX2PHYSTATUS_delay = PIPERX2PHYSTATUS;
  assign #(in_delay) PIPERX2STARTBLOCK_delay = PIPERX2STARTBLOCK;
  assign #(in_delay) PIPERX2VALID_delay = PIPERX2VALID;
  assign #(in_delay) PIPERX3DATAVALID_delay = PIPERX3DATAVALID;
  assign #(in_delay) PIPERX3ELECIDLE_delay = PIPERX3ELECIDLE;
  assign #(in_delay) PIPERX3EQDONE_delay = PIPERX3EQDONE;
  assign #(in_delay) PIPERX3EQLPADAPTDONE_delay = PIPERX3EQLPADAPTDONE;
  assign #(in_delay) PIPERX3EQLPLFFSSEL_delay = PIPERX3EQLPLFFSSEL;
  assign #(in_delay) PIPERX3PHYSTATUS_delay = PIPERX3PHYSTATUS;
  assign #(in_delay) PIPERX3STARTBLOCK_delay = PIPERX3STARTBLOCK;
  assign #(in_delay) PIPERX3VALID_delay = PIPERX3VALID;
  assign #(in_delay) PIPERX4DATAVALID_delay = PIPERX4DATAVALID;
  assign #(in_delay) PIPERX4ELECIDLE_delay = PIPERX4ELECIDLE;
  assign #(in_delay) PIPERX4EQDONE_delay = PIPERX4EQDONE;
  assign #(in_delay) PIPERX4EQLPADAPTDONE_delay = PIPERX4EQLPADAPTDONE;
  assign #(in_delay) PIPERX4EQLPLFFSSEL_delay = PIPERX4EQLPLFFSSEL;
  assign #(in_delay) PIPERX4PHYSTATUS_delay = PIPERX4PHYSTATUS;
  assign #(in_delay) PIPERX4STARTBLOCK_delay = PIPERX4STARTBLOCK;
  assign #(in_delay) PIPERX4VALID_delay = PIPERX4VALID;
  assign #(in_delay) PIPERX5DATAVALID_delay = PIPERX5DATAVALID;
  assign #(in_delay) PIPERX5ELECIDLE_delay = PIPERX5ELECIDLE;
  assign #(in_delay) PIPERX5EQDONE_delay = PIPERX5EQDONE;
  assign #(in_delay) PIPERX5EQLPADAPTDONE_delay = PIPERX5EQLPADAPTDONE;
  assign #(in_delay) PIPERX5EQLPLFFSSEL_delay = PIPERX5EQLPLFFSSEL;
  assign #(in_delay) PIPERX5PHYSTATUS_delay = PIPERX5PHYSTATUS;
  assign #(in_delay) PIPERX5STARTBLOCK_delay = PIPERX5STARTBLOCK;
  assign #(in_delay) PIPERX5VALID_delay = PIPERX5VALID;
  assign #(in_delay) PIPERX6DATAVALID_delay = PIPERX6DATAVALID;
  assign #(in_delay) PIPERX6ELECIDLE_delay = PIPERX6ELECIDLE;
  assign #(in_delay) PIPERX6EQDONE_delay = PIPERX6EQDONE;
  assign #(in_delay) PIPERX6EQLPADAPTDONE_delay = PIPERX6EQLPADAPTDONE;
  assign #(in_delay) PIPERX6EQLPLFFSSEL_delay = PIPERX6EQLPLFFSSEL;
  assign #(in_delay) PIPERX6PHYSTATUS_delay = PIPERX6PHYSTATUS;
  assign #(in_delay) PIPERX6STARTBLOCK_delay = PIPERX6STARTBLOCK;
  assign #(in_delay) PIPERX6VALID_delay = PIPERX6VALID;
  assign #(in_delay) PIPERX7DATAVALID_delay = PIPERX7DATAVALID;
  assign #(in_delay) PIPERX7ELECIDLE_delay = PIPERX7ELECIDLE;
  assign #(in_delay) PIPERX7EQDONE_delay = PIPERX7EQDONE;
  assign #(in_delay) PIPERX7EQLPADAPTDONE_delay = PIPERX7EQLPADAPTDONE;
  assign #(in_delay) PIPERX7EQLPLFFSSEL_delay = PIPERX7EQLPLFFSSEL;
  assign #(in_delay) PIPERX7PHYSTATUS_delay = PIPERX7PHYSTATUS;
  assign #(in_delay) PIPERX7STARTBLOCK_delay = PIPERX7STARTBLOCK;
  assign #(in_delay) PIPERX7VALID_delay = PIPERX7VALID;
  assign #(in_delay) PIPETX0EQDONE_delay = PIPETX0EQDONE;
  assign #(in_delay) PIPETX1EQDONE_delay = PIPETX1EQDONE;
  assign #(in_delay) PIPETX2EQDONE_delay = PIPETX2EQDONE;
  assign #(in_delay) PIPETX3EQDONE_delay = PIPETX3EQDONE;
  assign #(in_delay) PIPETX4EQDONE_delay = PIPETX4EQDONE;
  assign #(in_delay) PIPETX5EQDONE_delay = PIPETX5EQDONE;
  assign #(in_delay) PIPETX6EQDONE_delay = PIPETX6EQDONE;
  assign #(in_delay) PIPETX7EQDONE_delay = PIPETX7EQDONE;
  assign #(in_delay) PLEQRESETEIEOSCOUNT_delay = PLEQRESETEIEOSCOUNT;
  assign #(in_delay) PLGEN2UPSTREAMPREFERDEEMPH_delay = PLGEN2UPSTREAMPREFERDEEMPH;
  assign #(in_delay) SAXISCCTLAST_delay = SAXISCCTLAST;
  assign #(in_delay) SAXISCCTVALID_delay = SAXISCCTVALID;
  assign #(in_delay) SAXISRQTLAST_delay = SAXISRQTLAST;
  assign #(in_delay) SAXISRQTVALID_delay = SAXISRQTVALID;
`endif //  `ifndef XIL_TIMING
// inputs with no timing checks

  assign #(in_delay) CFGDEVID_delay = CFGDEVID;
  assign #(in_delay) CFGDSBUSNUMBER_delay = CFGDSBUSNUMBER;
  assign #(in_delay) CFGDSDEVICENUMBER_delay = CFGDSDEVICENUMBER;
  assign #(in_delay) CFGDSFUNCTIONNUMBER_delay = CFGDSFUNCTIONNUMBER;
  assign #(in_delay) CFGDSN_delay = CFGDSN;
  assign #(in_delay) CFGDSPORTNUMBER_delay = CFGDSPORTNUMBER;
  assign #(in_delay) CFGEXTREADDATA_delay = CFGEXTREADDATA;
  assign #(in_delay) CFGFCSEL_delay = CFGFCSEL;
  assign #(in_delay) CFGFLRDONE_delay = CFGFLRDONE;
  assign #(in_delay) CFGINTERRUPTINT_delay = CFGINTERRUPTINT;
  assign #(in_delay) CFGINTERRUPTMSIATTR_delay = CFGINTERRUPTMSIATTR;
  assign #(in_delay) CFGINTERRUPTMSIFUNCTIONNUMBER_delay = CFGINTERRUPTMSIFUNCTIONNUMBER;
  assign #(in_delay) CFGINTERRUPTMSIINT_delay = CFGINTERRUPTMSIINT;
  assign #(in_delay) CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM_delay = CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM;
  assign #(in_delay) CFGINTERRUPTMSIPENDINGSTATUS_delay = CFGINTERRUPTMSIPENDINGSTATUS;
  assign #(in_delay) CFGINTERRUPTMSISELECT_delay = CFGINTERRUPTMSISELECT;
  assign #(in_delay) CFGINTERRUPTMSITPHSTTAG_delay = CFGINTERRUPTMSITPHSTTAG;
  assign #(in_delay) CFGINTERRUPTMSITPHTYPE_delay = CFGINTERRUPTMSITPHTYPE;
  assign #(in_delay) CFGINTERRUPTMSIXADDRESS_delay = CFGINTERRUPTMSIXADDRESS;
  assign #(in_delay) CFGINTERRUPTMSIXDATA_delay = CFGINTERRUPTMSIXDATA;
  assign #(in_delay) CFGINTERRUPTPENDING_delay = CFGINTERRUPTPENDING;
  assign #(in_delay) CFGMGMTADDR_delay = CFGMGMTADDR;
  assign #(in_delay) CFGMGMTBYTEENABLE_delay = CFGMGMTBYTEENABLE;
  assign #(in_delay) CFGMGMTWRITEDATA_delay = CFGMGMTWRITEDATA;
  assign #(in_delay) CFGMSGTRANSMITDATA_delay = CFGMSGTRANSMITDATA;
  assign #(in_delay) CFGMSGTRANSMITTYPE_delay = CFGMSGTRANSMITTYPE;
  assign #(in_delay) CFGPERFUNCSTATUSCONTROL_delay = CFGPERFUNCSTATUSCONTROL;
  assign #(in_delay) CFGPERFUNCTIONNUMBER_delay = CFGPERFUNCTIONNUMBER;
  assign #(in_delay) CFGREVID_delay = CFGREVID;
  assign #(in_delay) CFGSUBSYSID_delay = CFGSUBSYSID;
  assign #(in_delay) CFGSUBSYSVENDID_delay = CFGSUBSYSVENDID;
  assign #(in_delay) CFGTPHSTTREADDATA_delay = CFGTPHSTTREADDATA;
  assign #(in_delay) CFGVENDID_delay = CFGVENDID;
  assign #(in_delay) CFGVFFLRDONE_delay = CFGVFFLRDONE;
  assign #(in_delay) CONFREQDATA_delay = CONFREQDATA;
  assign #(in_delay) CONFREQREGNUM_delay = CONFREQREGNUM;
  assign #(in_delay) CONFREQTYPE_delay = CONFREQTYPE;
  assign #(in_delay) DBGDATASEL_delay = DBGDATASEL;
  assign #(in_delay) DRPADDR_delay = DRPADDR;
  assign #(in_delay) DRPDI_delay = DRPDI;
  assign #(in_delay) LL2LMSAXISTXTUSER_delay = LL2LMSAXISTXTUSER;
  assign #(in_delay) LL2LMTXTLPID0_delay = LL2LMTXTLPID0;
  assign #(in_delay) LL2LMTXTLPID1_delay = LL2LMTXTLPID1;
  assign #(in_delay) MAXISCQTREADY_delay = MAXISCQTREADY;
  assign #(in_delay) MAXISRCTREADY_delay = MAXISRCTREADY;
  assign #(in_delay) MCAPPERST0B_delay = MCAPPERST0B;
  assign #(in_delay) MCAPPERST1B_delay = MCAPPERST1B;
  assign #(in_delay) MGMTRESETN_delay = MGMTRESETN;
  assign #(in_delay) MGMTSTICKYRESETN_delay = MGMTSTICKYRESETN;
  assign #(in_delay) MICOMPLETIONRAMREADDATA_delay = MICOMPLETIONRAMREADDATA;
  assign #(in_delay) MIREPLAYRAMREADDATA_delay = MIREPLAYRAMREADDATA;
  assign #(in_delay) MIREQUESTRAMREADDATA_delay = MIREQUESTRAMREADDATA;
  assign #(in_delay) PIPEEQFS_delay = PIPEEQFS;
  assign #(in_delay) PIPEEQLF_delay = PIPEEQLF;
  assign #(in_delay) PIPERESETN_delay = PIPERESETN;
  assign #(in_delay) PIPERX0CHARISK_delay = PIPERX0CHARISK;
  assign #(in_delay) PIPERX0DATA_delay = PIPERX0DATA;
  assign #(in_delay) PIPERX0EQLPNEWTXCOEFFORPRESET_delay = PIPERX0EQLPNEWTXCOEFFORPRESET;
  assign #(in_delay) PIPERX0STATUS_delay = PIPERX0STATUS;
  assign #(in_delay) PIPERX0SYNCHEADER_delay = PIPERX0SYNCHEADER;
  assign #(in_delay) PIPERX1CHARISK_delay = PIPERX1CHARISK;
  assign #(in_delay) PIPERX1DATA_delay = PIPERX1DATA;
  assign #(in_delay) PIPERX1EQLPNEWTXCOEFFORPRESET_delay = PIPERX1EQLPNEWTXCOEFFORPRESET;
  assign #(in_delay) PIPERX1STATUS_delay = PIPERX1STATUS;
  assign #(in_delay) PIPERX1SYNCHEADER_delay = PIPERX1SYNCHEADER;
  assign #(in_delay) PIPERX2CHARISK_delay = PIPERX2CHARISK;
  assign #(in_delay) PIPERX2DATA_delay = PIPERX2DATA;
  assign #(in_delay) PIPERX2EQLPNEWTXCOEFFORPRESET_delay = PIPERX2EQLPNEWTXCOEFFORPRESET;
  assign #(in_delay) PIPERX2STATUS_delay = PIPERX2STATUS;
  assign #(in_delay) PIPERX2SYNCHEADER_delay = PIPERX2SYNCHEADER;
  assign #(in_delay) PIPERX3CHARISK_delay = PIPERX3CHARISK;
  assign #(in_delay) PIPERX3DATA_delay = PIPERX3DATA;
  assign #(in_delay) PIPERX3EQLPNEWTXCOEFFORPRESET_delay = PIPERX3EQLPNEWTXCOEFFORPRESET;
  assign #(in_delay) PIPERX3STATUS_delay = PIPERX3STATUS;
  assign #(in_delay) PIPERX3SYNCHEADER_delay = PIPERX3SYNCHEADER;
  assign #(in_delay) PIPERX4CHARISK_delay = PIPERX4CHARISK;
  assign #(in_delay) PIPERX4DATA_delay = PIPERX4DATA;
  assign #(in_delay) PIPERX4EQLPNEWTXCOEFFORPRESET_delay = PIPERX4EQLPNEWTXCOEFFORPRESET;
  assign #(in_delay) PIPERX4STATUS_delay = PIPERX4STATUS;
  assign #(in_delay) PIPERX4SYNCHEADER_delay = PIPERX4SYNCHEADER;
  assign #(in_delay) PIPERX5CHARISK_delay = PIPERX5CHARISK;
  assign #(in_delay) PIPERX5DATA_delay = PIPERX5DATA;
  assign #(in_delay) PIPERX5EQLPNEWTXCOEFFORPRESET_delay = PIPERX5EQLPNEWTXCOEFFORPRESET;
  assign #(in_delay) PIPERX5STATUS_delay = PIPERX5STATUS;
  assign #(in_delay) PIPERX5SYNCHEADER_delay = PIPERX5SYNCHEADER;
  assign #(in_delay) PIPERX6CHARISK_delay = PIPERX6CHARISK;
  assign #(in_delay) PIPERX6DATA_delay = PIPERX6DATA;
  assign #(in_delay) PIPERX6EQLPNEWTXCOEFFORPRESET_delay = PIPERX6EQLPNEWTXCOEFFORPRESET;
  assign #(in_delay) PIPERX6STATUS_delay = PIPERX6STATUS;
  assign #(in_delay) PIPERX6SYNCHEADER_delay = PIPERX6SYNCHEADER;
  assign #(in_delay) PIPERX7CHARISK_delay = PIPERX7CHARISK;
  assign #(in_delay) PIPERX7DATA_delay = PIPERX7DATA;
  assign #(in_delay) PIPERX7EQLPNEWTXCOEFFORPRESET_delay = PIPERX7EQLPNEWTXCOEFFORPRESET;
  assign #(in_delay) PIPERX7STATUS_delay = PIPERX7STATUS;
  assign #(in_delay) PIPERX7SYNCHEADER_delay = PIPERX7SYNCHEADER;
  assign #(in_delay) PIPETX0EQCOEFF_delay = PIPETX0EQCOEFF;
  assign #(in_delay) PIPETX1EQCOEFF_delay = PIPETX1EQCOEFF;
  assign #(in_delay) PIPETX2EQCOEFF_delay = PIPETX2EQCOEFF;
  assign #(in_delay) PIPETX3EQCOEFF_delay = PIPETX3EQCOEFF;
  assign #(in_delay) PIPETX4EQCOEFF_delay = PIPETX4EQCOEFF;
  assign #(in_delay) PIPETX5EQCOEFF_delay = PIPETX5EQCOEFF;
  assign #(in_delay) PIPETX6EQCOEFF_delay = PIPETX6EQCOEFF;
  assign #(in_delay) PIPETX7EQCOEFF_delay = PIPETX7EQCOEFF;
  assign #(in_delay) RESETN_delay = RESETN;
  assign #(in_delay) SAXISCCTDATA_delay = SAXISCCTDATA;
  assign #(in_delay) SAXISCCTKEEP_delay = SAXISCCTKEEP;
  assign #(in_delay) SAXISCCTUSER_delay = SAXISCCTUSER;
  assign #(in_delay) SAXISRQTDATA_delay = SAXISRQTDATA;
  assign #(in_delay) SAXISRQTKEEP_delay = SAXISRQTKEEP;
  assign #(in_delay) SAXISRQTUSER_delay = SAXISRQTUSER;
  assign #(in_delay) SPAREIN_delay = SPAREIN;

  assign CFGCURRENTSPEED_delay = CFGCURRENTSPEED_out;
  assign CFGDPASUBSTATECHANGE_delay = CFGDPASUBSTATECHANGE_out;
  assign CFGERRCOROUT_delay = CFGERRCOROUT_out;
  assign CFGERRFATALOUT_delay = CFGERRFATALOUT_out;
  assign CFGERRNONFATALOUT_delay = CFGERRNONFATALOUT_out;
  assign CFGEXTFUNCTIONNUMBER_delay = CFGEXTFUNCTIONNUMBER_out;
  assign CFGEXTREADRECEIVED_delay = CFGEXTREADRECEIVED_out;
  assign CFGEXTREGISTERNUMBER_delay = CFGEXTREGISTERNUMBER_out;
  assign CFGEXTWRITEBYTEENABLE_delay = CFGEXTWRITEBYTEENABLE_out;
  assign CFGEXTWRITEDATA_delay = CFGEXTWRITEDATA_out;
  assign CFGEXTWRITERECEIVED_delay = CFGEXTWRITERECEIVED_out;
  assign CFGFCCPLD_delay = CFGFCCPLD_out;
  assign CFGFCCPLH_delay = CFGFCCPLH_out;
  assign CFGFCNPD_delay = CFGFCNPD_out;
  assign CFGFCNPH_delay = CFGFCNPH_out;
  assign CFGFCPD_delay = CFGFCPD_out;
  assign CFGFCPH_delay = CFGFCPH_out;
  assign CFGFLRINPROCESS_delay = CFGFLRINPROCESS_out;
  assign CFGFUNCTIONPOWERSTATE_delay = CFGFUNCTIONPOWERSTATE_out;
  assign CFGFUNCTIONSTATUS_delay = CFGFUNCTIONSTATUS_out;
  assign CFGHOTRESETOUT_delay = CFGHOTRESETOUT_out;
  assign CFGINTERRUPTMSIDATA_delay = CFGINTERRUPTMSIDATA_out;
  assign CFGINTERRUPTMSIENABLE_delay = CFGINTERRUPTMSIENABLE_out;
  assign CFGINTERRUPTMSIFAIL_delay = CFGINTERRUPTMSIFAIL_out;
  assign CFGINTERRUPTMSIMASKUPDATE_delay = CFGINTERRUPTMSIMASKUPDATE_out;
  assign CFGINTERRUPTMSIMMENABLE_delay = CFGINTERRUPTMSIMMENABLE_out;
  assign CFGINTERRUPTMSISENT_delay = CFGINTERRUPTMSISENT_out;
  assign CFGINTERRUPTMSIVFENABLE_delay = CFGINTERRUPTMSIVFENABLE_out;
  assign CFGINTERRUPTMSIXENABLE_delay = CFGINTERRUPTMSIXENABLE_out;
  assign CFGINTERRUPTMSIXFAIL_delay = CFGINTERRUPTMSIXFAIL_out;
  assign CFGINTERRUPTMSIXMASK_delay = CFGINTERRUPTMSIXMASK_out;
  assign CFGINTERRUPTMSIXSENT_delay = CFGINTERRUPTMSIXSENT_out;
  assign CFGINTERRUPTMSIXVFENABLE_delay = CFGINTERRUPTMSIXVFENABLE_out;
  assign CFGINTERRUPTMSIXVFMASK_delay = CFGINTERRUPTMSIXVFMASK_out;
  assign CFGINTERRUPTSENT_delay = CFGINTERRUPTSENT_out;
  assign CFGLINKPOWERSTATE_delay = CFGLINKPOWERSTATE_out;
  assign CFGLOCALERROR_delay = CFGLOCALERROR_out;
  assign CFGLTRENABLE_delay = CFGLTRENABLE_out;
  assign CFGLTSSMSTATE_delay = CFGLTSSMSTATE_out;
  assign CFGMAXPAYLOAD_delay = CFGMAXPAYLOAD_out;
  assign CFGMAXREADREQ_delay = CFGMAXREADREQ_out;
  assign CFGMGMTREADDATA_delay = CFGMGMTREADDATA_out;
  assign CFGMGMTREADWRITEDONE_delay = CFGMGMTREADWRITEDONE_out;
  assign CFGMSGRECEIVEDDATA_delay = CFGMSGRECEIVEDDATA_out;
  assign CFGMSGRECEIVEDTYPE_delay = CFGMSGRECEIVEDTYPE_out;
  assign CFGMSGRECEIVED_delay = CFGMSGRECEIVED_out;
  assign CFGMSGTRANSMITDONE_delay = CFGMSGTRANSMITDONE_out;
  assign CFGNEGOTIATEDWIDTH_delay = CFGNEGOTIATEDWIDTH_out;
  assign CFGOBFFENABLE_delay = CFGOBFFENABLE_out;
  assign CFGPERFUNCSTATUSDATA_delay = CFGPERFUNCSTATUSDATA_out;
  assign CFGPERFUNCTIONUPDATEDONE_delay = CFGPERFUNCTIONUPDATEDONE_out;
  assign CFGPHYLINKDOWN_delay = CFGPHYLINKDOWN_out;
  assign CFGPHYLINKSTATUS_delay = CFGPHYLINKSTATUS_out;
  assign CFGPLSTATUSCHANGE_delay = CFGPLSTATUSCHANGE_out;
  assign CFGPOWERSTATECHANGEINTERRUPT_delay = CFGPOWERSTATECHANGEINTERRUPT_out;
  assign CFGRCBSTATUS_delay = CFGRCBSTATUS_out;
  assign CFGTPHFUNCTIONNUM_delay = CFGTPHFUNCTIONNUM_out;
  assign CFGTPHREQUESTERENABLE_delay = CFGTPHREQUESTERENABLE_out;
  assign CFGTPHSTMODE_delay = CFGTPHSTMODE_out;
  assign CFGTPHSTTADDRESS_delay = CFGTPHSTTADDRESS_out;
  assign CFGTPHSTTREADENABLE_delay = CFGTPHSTTREADENABLE_out;
  assign CFGTPHSTTWRITEBYTEVALID_delay = CFGTPHSTTWRITEBYTEVALID_out;
  assign CFGTPHSTTWRITEDATA_delay = CFGTPHSTTWRITEDATA_out;
  assign CFGTPHSTTWRITEENABLE_delay = CFGTPHSTTWRITEENABLE_out;
  assign CFGVFFLRINPROCESS_delay = CFGVFFLRINPROCESS_out;
  assign CFGVFPOWERSTATE_delay = CFGVFPOWERSTATE_out;
  assign CFGVFSTATUS_delay = CFGVFSTATUS_out;
  assign CFGVFTPHREQUESTERENABLE_delay = CFGVFTPHREQUESTERENABLE_out;
  assign CFGVFTPHSTMODE_delay = CFGVFTPHSTMODE_out;
  assign CONFMCAPDESIGNSWITCH_delay = CONFMCAPDESIGNSWITCH_out;
  assign CONFMCAPEOS_delay = CONFMCAPEOS_out;
  assign CONFMCAPINUSEBYPCIE_delay = CONFMCAPINUSEBYPCIE_out;
  assign CONFREQREADY_delay = CONFREQREADY_out;
  assign CONFRESPRDATA_delay = CONFRESPRDATA_out;
  assign CONFRESPVALID_delay = CONFRESPVALID_out;
  assign DBGDATAOUT_delay = DBGDATAOUT_out;
  assign DBGMCAPCSB_delay = DBGMCAPCSB_out;
  assign DBGMCAPDATA_delay = DBGMCAPDATA_out;
  assign DBGMCAPEOS_delay = DBGMCAPEOS_out;
  assign DBGMCAPERROR_delay = DBGMCAPERROR_out;
  assign DBGMCAPMODE_delay = DBGMCAPMODE_out;
  assign DBGMCAPRDATAVALID_delay = DBGMCAPRDATAVALID_out;
  assign DBGMCAPRDWRB_delay = DBGMCAPRDWRB_out;
  assign DBGMCAPRESET_delay = DBGMCAPRESET_out;
  assign DBGPLDATABLOCKRECEIVEDAFTEREDS_delay = DBGPLDATABLOCKRECEIVEDAFTEREDS_out;
  assign DBGPLGEN3FRAMINGERRORDETECTED_delay = DBGPLGEN3FRAMINGERRORDETECTED_out;
  assign DBGPLGEN3SYNCHEADERERRORDETECTED_delay = DBGPLGEN3SYNCHEADERERRORDETECTED_out;
  assign DBGPLINFERREDRXELECTRICALIDLE_delay = DBGPLINFERREDRXELECTRICALIDLE_out;
  assign DRPDO_delay = DRPDO_out;
  assign DRPRDY_delay = DRPRDY_out;
  assign LL2LMMASTERTLPSENT0_delay = LL2LMMASTERTLPSENT0_out;
  assign LL2LMMASTERTLPSENT1_delay = LL2LMMASTERTLPSENT1_out;
  assign LL2LMMASTERTLPSENTTLPID0_delay = LL2LMMASTERTLPSENTTLPID0_out;
  assign LL2LMMASTERTLPSENTTLPID1_delay = LL2LMMASTERTLPSENTTLPID1_out;
  assign LL2LMMAXISRXTDATA_delay = LL2LMMAXISRXTDATA_out;
  assign LL2LMMAXISRXTUSER_delay = LL2LMMAXISRXTUSER_out;
  assign LL2LMMAXISRXTVALID_delay = LL2LMMAXISRXTVALID_out;
  assign LL2LMSAXISTXTREADY_delay = LL2LMSAXISTXTREADY_out;
  assign MAXISCQTDATA_delay = MAXISCQTDATA_out;
  assign MAXISCQTKEEP_delay = MAXISCQTKEEP_out;
  assign MAXISCQTLAST_delay = MAXISCQTLAST_out;
  assign MAXISCQTUSER_delay = MAXISCQTUSER_out;
  assign MAXISCQTVALID_delay = MAXISCQTVALID_out;
  assign MAXISRCTDATA_delay = MAXISRCTDATA_out;
  assign MAXISRCTKEEP_delay = MAXISRCTKEEP_out;
  assign MAXISRCTLAST_delay = MAXISRCTLAST_out;
  assign MAXISRCTUSER_delay = MAXISRCTUSER_out;
  assign MAXISRCTVALID_delay = MAXISRCTVALID_out;
  assign MICOMPLETIONRAMREADADDRESSAL_delay = MICOMPLETIONRAMREADADDRESSAL_out;
  assign MICOMPLETIONRAMREADADDRESSAU_delay = MICOMPLETIONRAMREADADDRESSAU_out;
  assign MICOMPLETIONRAMREADADDRESSBL_delay = MICOMPLETIONRAMREADADDRESSBL_out;
  assign MICOMPLETIONRAMREADADDRESSBU_delay = MICOMPLETIONRAMREADADDRESSBU_out;
  assign MICOMPLETIONRAMREADENABLEL_delay = MICOMPLETIONRAMREADENABLEL_out;
  assign MICOMPLETIONRAMREADENABLEU_delay = MICOMPLETIONRAMREADENABLEU_out;
  assign MICOMPLETIONRAMWRITEADDRESSAL_delay = MICOMPLETIONRAMWRITEADDRESSAL_out;
  assign MICOMPLETIONRAMWRITEADDRESSAU_delay = MICOMPLETIONRAMWRITEADDRESSAU_out;
  assign MICOMPLETIONRAMWRITEADDRESSBL_delay = MICOMPLETIONRAMWRITEADDRESSBL_out;
  assign MICOMPLETIONRAMWRITEADDRESSBU_delay = MICOMPLETIONRAMWRITEADDRESSBU_out;
  assign MICOMPLETIONRAMWRITEDATAL_delay = MICOMPLETIONRAMWRITEDATAL_out;
  assign MICOMPLETIONRAMWRITEDATAU_delay = MICOMPLETIONRAMWRITEDATAU_out;
  assign MICOMPLETIONRAMWRITEENABLEL_delay = MICOMPLETIONRAMWRITEENABLEL_out;
  assign MICOMPLETIONRAMWRITEENABLEU_delay = MICOMPLETIONRAMWRITEENABLEU_out;
  assign MIREPLAYRAMADDRESS_delay = MIREPLAYRAMADDRESS_out;
  assign MIREPLAYRAMREADENABLE_delay = MIREPLAYRAMREADENABLE_out;
  assign MIREPLAYRAMWRITEDATA_delay = MIREPLAYRAMWRITEDATA_out;
  assign MIREPLAYRAMWRITEENABLE_delay = MIREPLAYRAMWRITEENABLE_out;
  assign MIREQUESTRAMREADADDRESSA_delay = MIREQUESTRAMREADADDRESSA_out;
  assign MIREQUESTRAMREADADDRESSB_delay = MIREQUESTRAMREADADDRESSB_out;
  assign MIREQUESTRAMREADENABLE_delay = MIREQUESTRAMREADENABLE_out;
  assign MIREQUESTRAMWRITEADDRESSA_delay = MIREQUESTRAMWRITEADDRESSA_out;
  assign MIREQUESTRAMWRITEADDRESSB_delay = MIREQUESTRAMWRITEADDRESSB_out;
  assign MIREQUESTRAMWRITEDATA_delay = MIREQUESTRAMWRITEDATA_out;
  assign MIREQUESTRAMWRITEENABLE_delay = MIREQUESTRAMWRITEENABLE_out;
  assign PCIECQNPREQCOUNT_delay = PCIECQNPREQCOUNT_out;
  assign PCIEPERST0B_delay = PCIEPERST0B_out;
  assign PCIEPERST1B_delay = PCIEPERST1B_out;
  assign PCIERQSEQNUMVLD_delay = PCIERQSEQNUMVLD_out;
  assign PCIERQSEQNUM_delay = PCIERQSEQNUM_out;
  assign PCIERQTAGAV_delay = PCIERQTAGAV_out;
  assign PCIERQTAGVLD_delay = PCIERQTAGVLD_out;
  assign PCIERQTAG_delay = PCIERQTAG_out;
  assign PCIETFCNPDAV_delay = PCIETFCNPDAV_out;
  assign PCIETFCNPHAV_delay = PCIETFCNPHAV_out;
  assign PIPERX0EQCONTROL_delay = PIPERX0EQCONTROL_out;
  assign PIPERX0EQLPLFFS_delay = PIPERX0EQLPLFFS_out;
  assign PIPERX0EQLPTXPRESET_delay = PIPERX0EQLPTXPRESET_out;
  assign PIPERX0EQPRESET_delay = PIPERX0EQPRESET_out;
  assign PIPERX0POLARITY_delay = PIPERX0POLARITY_out;
  assign PIPERX1EQCONTROL_delay = PIPERX1EQCONTROL_out;
  assign PIPERX1EQLPLFFS_delay = PIPERX1EQLPLFFS_out;
  assign PIPERX1EQLPTXPRESET_delay = PIPERX1EQLPTXPRESET_out;
  assign PIPERX1EQPRESET_delay = PIPERX1EQPRESET_out;
  assign PIPERX1POLARITY_delay = PIPERX1POLARITY_out;
  assign PIPERX2EQCONTROL_delay = PIPERX2EQCONTROL_out;
  assign PIPERX2EQLPLFFS_delay = PIPERX2EQLPLFFS_out;
  assign PIPERX2EQLPTXPRESET_delay = PIPERX2EQLPTXPRESET_out;
  assign PIPERX2EQPRESET_delay = PIPERX2EQPRESET_out;
  assign PIPERX2POLARITY_delay = PIPERX2POLARITY_out;
  assign PIPERX3EQCONTROL_delay = PIPERX3EQCONTROL_out;
  assign PIPERX3EQLPLFFS_delay = PIPERX3EQLPLFFS_out;
  assign PIPERX3EQLPTXPRESET_delay = PIPERX3EQLPTXPRESET_out;
  assign PIPERX3EQPRESET_delay = PIPERX3EQPRESET_out;
  assign PIPERX3POLARITY_delay = PIPERX3POLARITY_out;
  assign PIPERX4EQCONTROL_delay = PIPERX4EQCONTROL_out;
  assign PIPERX4EQLPLFFS_delay = PIPERX4EQLPLFFS_out;
  assign PIPERX4EQLPTXPRESET_delay = PIPERX4EQLPTXPRESET_out;
  assign PIPERX4EQPRESET_delay = PIPERX4EQPRESET_out;
  assign PIPERX4POLARITY_delay = PIPERX4POLARITY_out;
  assign PIPERX5EQCONTROL_delay = PIPERX5EQCONTROL_out;
  assign PIPERX5EQLPLFFS_delay = PIPERX5EQLPLFFS_out;
  assign PIPERX5EQLPTXPRESET_delay = PIPERX5EQLPTXPRESET_out;
  assign PIPERX5EQPRESET_delay = PIPERX5EQPRESET_out;
  assign PIPERX5POLARITY_delay = PIPERX5POLARITY_out;
  assign PIPERX6EQCONTROL_delay = PIPERX6EQCONTROL_out;
  assign PIPERX6EQLPLFFS_delay = PIPERX6EQLPLFFS_out;
  assign PIPERX6EQLPTXPRESET_delay = PIPERX6EQLPTXPRESET_out;
  assign PIPERX6EQPRESET_delay = PIPERX6EQPRESET_out;
  assign PIPERX6POLARITY_delay = PIPERX6POLARITY_out;
  assign PIPERX7EQCONTROL_delay = PIPERX7EQCONTROL_out;
  assign PIPERX7EQLPLFFS_delay = PIPERX7EQLPLFFS_out;
  assign PIPERX7EQLPTXPRESET_delay = PIPERX7EQLPTXPRESET_out;
  assign PIPERX7EQPRESET_delay = PIPERX7EQPRESET_out;
  assign PIPERX7POLARITY_delay = PIPERX7POLARITY_out;
  assign PIPETX0CHARISK_delay = PIPETX0CHARISK_out;
  assign PIPETX0COMPLIANCE_delay = PIPETX0COMPLIANCE_out;
  assign PIPETX0DATAVALID_delay = PIPETX0DATAVALID_out;
  assign PIPETX0DATA_delay = PIPETX0DATA_out;
  assign PIPETX0DEEMPH_delay = PIPETX0DEEMPH_out;
  assign PIPETX0ELECIDLE_delay = PIPETX0ELECIDLE_out;
  assign PIPETX0EQCONTROL_delay = PIPETX0EQCONTROL_out;
  assign PIPETX0EQDEEMPH_delay = PIPETX0EQDEEMPH_out;
  assign PIPETX0EQPRESET_delay = PIPETX0EQPRESET_out;
  assign PIPETX0MARGIN_delay = PIPETX0MARGIN_out;
  assign PIPETX0POWERDOWN_delay = PIPETX0POWERDOWN_out;
  assign PIPETX0RATE_delay = PIPETX0RATE_out;
  assign PIPETX0RCVRDET_delay = PIPETX0RCVRDET_out;
  assign PIPETX0RESET_delay = PIPETX0RESET_out;
  assign PIPETX0STARTBLOCK_delay = PIPETX0STARTBLOCK_out;
  assign PIPETX0SWING_delay = PIPETX0SWING_out;
  assign PIPETX0SYNCHEADER_delay = PIPETX0SYNCHEADER_out;
  assign PIPETX1CHARISK_delay = PIPETX1CHARISK_out;
  assign PIPETX1COMPLIANCE_delay = PIPETX1COMPLIANCE_out;
  assign PIPETX1DATAVALID_delay = PIPETX1DATAVALID_out;
  assign PIPETX1DATA_delay = PIPETX1DATA_out;
  assign PIPETX1DEEMPH_delay = PIPETX1DEEMPH_out;
  assign PIPETX1ELECIDLE_delay = PIPETX1ELECIDLE_out;
  assign PIPETX1EQCONTROL_delay = PIPETX1EQCONTROL_out;
  assign PIPETX1EQDEEMPH_delay = PIPETX1EQDEEMPH_out;
  assign PIPETX1EQPRESET_delay = PIPETX1EQPRESET_out;
  assign PIPETX1MARGIN_delay = PIPETX1MARGIN_out;
  assign PIPETX1POWERDOWN_delay = PIPETX1POWERDOWN_out;
  assign PIPETX1RATE_delay = PIPETX1RATE_out;
  assign PIPETX1RCVRDET_delay = PIPETX1RCVRDET_out;
  assign PIPETX1RESET_delay = PIPETX1RESET_out;
  assign PIPETX1STARTBLOCK_delay = PIPETX1STARTBLOCK_out;
  assign PIPETX1SWING_delay = PIPETX1SWING_out;
  assign PIPETX1SYNCHEADER_delay = PIPETX1SYNCHEADER_out;
  assign PIPETX2CHARISK_delay = PIPETX2CHARISK_out;
  assign PIPETX2COMPLIANCE_delay = PIPETX2COMPLIANCE_out;
  assign PIPETX2DATAVALID_delay = PIPETX2DATAVALID_out;
  assign PIPETX2DATA_delay = PIPETX2DATA_out;
  assign PIPETX2DEEMPH_delay = PIPETX2DEEMPH_out;
  assign PIPETX2ELECIDLE_delay = PIPETX2ELECIDLE_out;
  assign PIPETX2EQCONTROL_delay = PIPETX2EQCONTROL_out;
  assign PIPETX2EQDEEMPH_delay = PIPETX2EQDEEMPH_out;
  assign PIPETX2EQPRESET_delay = PIPETX2EQPRESET_out;
  assign PIPETX2MARGIN_delay = PIPETX2MARGIN_out;
  assign PIPETX2POWERDOWN_delay = PIPETX2POWERDOWN_out;
  assign PIPETX2RATE_delay = PIPETX2RATE_out;
  assign PIPETX2RCVRDET_delay = PIPETX2RCVRDET_out;
  assign PIPETX2RESET_delay = PIPETX2RESET_out;
  assign PIPETX2STARTBLOCK_delay = PIPETX2STARTBLOCK_out;
  assign PIPETX2SWING_delay = PIPETX2SWING_out;
  assign PIPETX2SYNCHEADER_delay = PIPETX2SYNCHEADER_out;
  assign PIPETX3CHARISK_delay = PIPETX3CHARISK_out;
  assign PIPETX3COMPLIANCE_delay = PIPETX3COMPLIANCE_out;
  assign PIPETX3DATAVALID_delay = PIPETX3DATAVALID_out;
  assign PIPETX3DATA_delay = PIPETX3DATA_out;
  assign PIPETX3DEEMPH_delay = PIPETX3DEEMPH_out;
  assign PIPETX3ELECIDLE_delay = PIPETX3ELECIDLE_out;
  assign PIPETX3EQCONTROL_delay = PIPETX3EQCONTROL_out;
  assign PIPETX3EQDEEMPH_delay = PIPETX3EQDEEMPH_out;
  assign PIPETX3EQPRESET_delay = PIPETX3EQPRESET_out;
  assign PIPETX3MARGIN_delay = PIPETX3MARGIN_out;
  assign PIPETX3POWERDOWN_delay = PIPETX3POWERDOWN_out;
  assign PIPETX3RATE_delay = PIPETX3RATE_out;
  assign PIPETX3RCVRDET_delay = PIPETX3RCVRDET_out;
  assign PIPETX3RESET_delay = PIPETX3RESET_out;
  assign PIPETX3STARTBLOCK_delay = PIPETX3STARTBLOCK_out;
  assign PIPETX3SWING_delay = PIPETX3SWING_out;
  assign PIPETX3SYNCHEADER_delay = PIPETX3SYNCHEADER_out;
  assign PIPETX4CHARISK_delay = PIPETX4CHARISK_out;
  assign PIPETX4COMPLIANCE_delay = PIPETX4COMPLIANCE_out;
  assign PIPETX4DATAVALID_delay = PIPETX4DATAVALID_out;
  assign PIPETX4DATA_delay = PIPETX4DATA_out;
  assign PIPETX4DEEMPH_delay = PIPETX4DEEMPH_out;
  assign PIPETX4ELECIDLE_delay = PIPETX4ELECIDLE_out;
  assign PIPETX4EQCONTROL_delay = PIPETX4EQCONTROL_out;
  assign PIPETX4EQDEEMPH_delay = PIPETX4EQDEEMPH_out;
  assign PIPETX4EQPRESET_delay = PIPETX4EQPRESET_out;
  assign PIPETX4MARGIN_delay = PIPETX4MARGIN_out;
  assign PIPETX4POWERDOWN_delay = PIPETX4POWERDOWN_out;
  assign PIPETX4RATE_delay = PIPETX4RATE_out;
  assign PIPETX4RCVRDET_delay = PIPETX4RCVRDET_out;
  assign PIPETX4RESET_delay = PIPETX4RESET_out;
  assign PIPETX4STARTBLOCK_delay = PIPETX4STARTBLOCK_out;
  assign PIPETX4SWING_delay = PIPETX4SWING_out;
  assign PIPETX4SYNCHEADER_delay = PIPETX4SYNCHEADER_out;
  assign PIPETX5CHARISK_delay = PIPETX5CHARISK_out;
  assign PIPETX5COMPLIANCE_delay = PIPETX5COMPLIANCE_out;
  assign PIPETX5DATAVALID_delay = PIPETX5DATAVALID_out;
  assign PIPETX5DATA_delay = PIPETX5DATA_out;
  assign PIPETX5DEEMPH_delay = PIPETX5DEEMPH_out;
  assign PIPETX5ELECIDLE_delay = PIPETX5ELECIDLE_out;
  assign PIPETX5EQCONTROL_delay = PIPETX5EQCONTROL_out;
  assign PIPETX5EQDEEMPH_delay = PIPETX5EQDEEMPH_out;
  assign PIPETX5EQPRESET_delay = PIPETX5EQPRESET_out;
  assign PIPETX5MARGIN_delay = PIPETX5MARGIN_out;
  assign PIPETX5POWERDOWN_delay = PIPETX5POWERDOWN_out;
  assign PIPETX5RATE_delay = PIPETX5RATE_out;
  assign PIPETX5RCVRDET_delay = PIPETX5RCVRDET_out;
  assign PIPETX5RESET_delay = PIPETX5RESET_out;
  assign PIPETX5STARTBLOCK_delay = PIPETX5STARTBLOCK_out;
  assign PIPETX5SWING_delay = PIPETX5SWING_out;
  assign PIPETX5SYNCHEADER_delay = PIPETX5SYNCHEADER_out;
  assign PIPETX6CHARISK_delay = PIPETX6CHARISK_out;
  assign PIPETX6COMPLIANCE_delay = PIPETX6COMPLIANCE_out;
  assign PIPETX6DATAVALID_delay = PIPETX6DATAVALID_out;
  assign PIPETX6DATA_delay = PIPETX6DATA_out;
  assign PIPETX6DEEMPH_delay = PIPETX6DEEMPH_out;
  assign PIPETX6ELECIDLE_delay = PIPETX6ELECIDLE_out;
  assign PIPETX6EQCONTROL_delay = PIPETX6EQCONTROL_out;
  assign PIPETX6EQDEEMPH_delay = PIPETX6EQDEEMPH_out;
  assign PIPETX6EQPRESET_delay = PIPETX6EQPRESET_out;
  assign PIPETX6MARGIN_delay = PIPETX6MARGIN_out;
  assign PIPETX6POWERDOWN_delay = PIPETX6POWERDOWN_out;
  assign PIPETX6RATE_delay = PIPETX6RATE_out;
  assign PIPETX6RCVRDET_delay = PIPETX6RCVRDET_out;
  assign PIPETX6RESET_delay = PIPETX6RESET_out;
  assign PIPETX6STARTBLOCK_delay = PIPETX6STARTBLOCK_out;
  assign PIPETX6SWING_delay = PIPETX6SWING_out;
  assign PIPETX6SYNCHEADER_delay = PIPETX6SYNCHEADER_out;
  assign PIPETX7CHARISK_delay = PIPETX7CHARISK_out;
  assign PIPETX7COMPLIANCE_delay = PIPETX7COMPLIANCE_out;
  assign PIPETX7DATAVALID_delay = PIPETX7DATAVALID_out;
  assign PIPETX7DATA_delay = PIPETX7DATA_out;
  assign PIPETX7DEEMPH_delay = PIPETX7DEEMPH_out;
  assign PIPETX7ELECIDLE_delay = PIPETX7ELECIDLE_out;
  assign PIPETX7EQCONTROL_delay = PIPETX7EQCONTROL_out;
  assign PIPETX7EQDEEMPH_delay = PIPETX7EQDEEMPH_out;
  assign PIPETX7EQPRESET_delay = PIPETX7EQPRESET_out;
  assign PIPETX7MARGIN_delay = PIPETX7MARGIN_out;
  assign PIPETX7POWERDOWN_delay = PIPETX7POWERDOWN_out;
  assign PIPETX7RATE_delay = PIPETX7RATE_out;
  assign PIPETX7RCVRDET_delay = PIPETX7RCVRDET_out;
  assign PIPETX7RESET_delay = PIPETX7RESET_out;
  assign PIPETX7STARTBLOCK_delay = PIPETX7STARTBLOCK_out;
  assign PIPETX7SWING_delay = PIPETX7SWING_out;
  assign PIPETX7SYNCHEADER_delay = PIPETX7SYNCHEADER_out;
  assign PLEQINPROGRESS_delay = PLEQINPROGRESS_out;
  assign PLEQPHASE_delay = PLEQPHASE_out;
  assign SAXISCCTREADY_delay = SAXISCCTREADY_out;
  assign SAXISRQTREADY_delay = SAXISRQTREADY_out;
  assign SPAREOUT_delay = SPAREOUT_out;

  assign CFGCONFIGSPACEENABLE_in = (CFGCONFIGSPACEENABLE === 1'bz) || CFGCONFIGSPACEENABLE_delay; // rv 1
  assign CFGDEVID_in[0] = (CFGDEVID[0] !== 1'bz) && CFGDEVID_delay[0]; // rv 0
  assign CFGDEVID_in[10] = (CFGDEVID[10] !== 1'bz) && CFGDEVID_delay[10]; // rv 0
  assign CFGDEVID_in[11] = (CFGDEVID[11] !== 1'bz) && CFGDEVID_delay[11]; // rv 0
  assign CFGDEVID_in[12] = (CFGDEVID[12] !== 1'bz) && CFGDEVID_delay[12]; // rv 0
  assign CFGDEVID_in[13] = (CFGDEVID[13] !== 1'bz) && CFGDEVID_delay[13]; // rv 0
  assign CFGDEVID_in[14] = (CFGDEVID[14] !== 1'bz) && CFGDEVID_delay[14]; // rv 0
  assign CFGDEVID_in[15] = (CFGDEVID[15] !== 1'bz) && CFGDEVID_delay[15]; // rv 0
  assign CFGDEVID_in[1] = (CFGDEVID[1] !== 1'bz) && CFGDEVID_delay[1]; // rv 0
  assign CFGDEVID_in[2] = (CFGDEVID[2] !== 1'bz) && CFGDEVID_delay[2]; // rv 0
  assign CFGDEVID_in[3] = (CFGDEVID[3] !== 1'bz) && CFGDEVID_delay[3]; // rv 0
  assign CFGDEVID_in[4] = (CFGDEVID[4] !== 1'bz) && CFGDEVID_delay[4]; // rv 0
  assign CFGDEVID_in[5] = (CFGDEVID[5] !== 1'bz) && CFGDEVID_delay[5]; // rv 0
  assign CFGDEVID_in[6] = (CFGDEVID[6] !== 1'bz) && CFGDEVID_delay[6]; // rv 0
  assign CFGDEVID_in[7] = (CFGDEVID[7] !== 1'bz) && CFGDEVID_delay[7]; // rv 0
  assign CFGDEVID_in[8] = (CFGDEVID[8] !== 1'bz) && CFGDEVID_delay[8]; // rv 0
  assign CFGDEVID_in[9] = (CFGDEVID[9] !== 1'bz) && CFGDEVID_delay[9]; // rv 0
  assign CFGDSBUSNUMBER_in[0] = (CFGDSBUSNUMBER[0] !== 1'bz) && CFGDSBUSNUMBER_delay[0]; // rv 0
  assign CFGDSBUSNUMBER_in[1] = (CFGDSBUSNUMBER[1] !== 1'bz) && CFGDSBUSNUMBER_delay[1]; // rv 0
  assign CFGDSBUSNUMBER_in[2] = (CFGDSBUSNUMBER[2] !== 1'bz) && CFGDSBUSNUMBER_delay[2]; // rv 0
  assign CFGDSBUSNUMBER_in[3] = (CFGDSBUSNUMBER[3] !== 1'bz) && CFGDSBUSNUMBER_delay[3]; // rv 0
  assign CFGDSBUSNUMBER_in[4] = (CFGDSBUSNUMBER[4] !== 1'bz) && CFGDSBUSNUMBER_delay[4]; // rv 0
  assign CFGDSBUSNUMBER_in[5] = (CFGDSBUSNUMBER[5] !== 1'bz) && CFGDSBUSNUMBER_delay[5]; // rv 0
  assign CFGDSBUSNUMBER_in[6] = (CFGDSBUSNUMBER[6] !== 1'bz) && CFGDSBUSNUMBER_delay[6]; // rv 0
  assign CFGDSBUSNUMBER_in[7] = (CFGDSBUSNUMBER[7] !== 1'bz) && CFGDSBUSNUMBER_delay[7]; // rv 0
  assign CFGDSDEVICENUMBER_in[0] = (CFGDSDEVICENUMBER[0] !== 1'bz) && CFGDSDEVICENUMBER_delay[0]; // rv 0
  assign CFGDSDEVICENUMBER_in[1] = (CFGDSDEVICENUMBER[1] !== 1'bz) && CFGDSDEVICENUMBER_delay[1]; // rv 0
  assign CFGDSDEVICENUMBER_in[2] = (CFGDSDEVICENUMBER[2] !== 1'bz) && CFGDSDEVICENUMBER_delay[2]; // rv 0
  assign CFGDSDEVICENUMBER_in[3] = (CFGDSDEVICENUMBER[3] !== 1'bz) && CFGDSDEVICENUMBER_delay[3]; // rv 0
  assign CFGDSDEVICENUMBER_in[4] = (CFGDSDEVICENUMBER[4] !== 1'bz) && CFGDSDEVICENUMBER_delay[4]; // rv 0
  assign CFGDSFUNCTIONNUMBER_in[0] = (CFGDSFUNCTIONNUMBER[0] !== 1'bz) && CFGDSFUNCTIONNUMBER_delay[0]; // rv 0
  assign CFGDSFUNCTIONNUMBER_in[1] = (CFGDSFUNCTIONNUMBER[1] !== 1'bz) && CFGDSFUNCTIONNUMBER_delay[1]; // rv 0
  assign CFGDSFUNCTIONNUMBER_in[2] = (CFGDSFUNCTIONNUMBER[2] !== 1'bz) && CFGDSFUNCTIONNUMBER_delay[2]; // rv 0
  assign CFGDSN_in[0] = (CFGDSN[0] !== 1'bz) && CFGDSN_delay[0]; // rv 0
  assign CFGDSN_in[10] = (CFGDSN[10] !== 1'bz) && CFGDSN_delay[10]; // rv 0
  assign CFGDSN_in[11] = (CFGDSN[11] !== 1'bz) && CFGDSN_delay[11]; // rv 0
  assign CFGDSN_in[12] = (CFGDSN[12] !== 1'bz) && CFGDSN_delay[12]; // rv 0
  assign CFGDSN_in[13] = (CFGDSN[13] !== 1'bz) && CFGDSN_delay[13]; // rv 0
  assign CFGDSN_in[14] = (CFGDSN[14] !== 1'bz) && CFGDSN_delay[14]; // rv 0
  assign CFGDSN_in[15] = (CFGDSN[15] !== 1'bz) && CFGDSN_delay[15]; // rv 0
  assign CFGDSN_in[16] = (CFGDSN[16] !== 1'bz) && CFGDSN_delay[16]; // rv 0
  assign CFGDSN_in[17] = (CFGDSN[17] !== 1'bz) && CFGDSN_delay[17]; // rv 0
  assign CFGDSN_in[18] = (CFGDSN[18] !== 1'bz) && CFGDSN_delay[18]; // rv 0
  assign CFGDSN_in[19] = (CFGDSN[19] !== 1'bz) && CFGDSN_delay[19]; // rv 0
  assign CFGDSN_in[1] = (CFGDSN[1] !== 1'bz) && CFGDSN_delay[1]; // rv 0
  assign CFGDSN_in[20] = (CFGDSN[20] !== 1'bz) && CFGDSN_delay[20]; // rv 0
  assign CFGDSN_in[21] = (CFGDSN[21] !== 1'bz) && CFGDSN_delay[21]; // rv 0
  assign CFGDSN_in[22] = (CFGDSN[22] !== 1'bz) && CFGDSN_delay[22]; // rv 0
  assign CFGDSN_in[23] = (CFGDSN[23] !== 1'bz) && CFGDSN_delay[23]; // rv 0
  assign CFGDSN_in[24] = (CFGDSN[24] !== 1'bz) && CFGDSN_delay[24]; // rv 0
  assign CFGDSN_in[25] = (CFGDSN[25] !== 1'bz) && CFGDSN_delay[25]; // rv 0
  assign CFGDSN_in[26] = (CFGDSN[26] !== 1'bz) && CFGDSN_delay[26]; // rv 0
  assign CFGDSN_in[27] = (CFGDSN[27] !== 1'bz) && CFGDSN_delay[27]; // rv 0
  assign CFGDSN_in[28] = (CFGDSN[28] !== 1'bz) && CFGDSN_delay[28]; // rv 0
  assign CFGDSN_in[29] = (CFGDSN[29] !== 1'bz) && CFGDSN_delay[29]; // rv 0
  assign CFGDSN_in[2] = (CFGDSN[2] !== 1'bz) && CFGDSN_delay[2]; // rv 0
  assign CFGDSN_in[30] = (CFGDSN[30] !== 1'bz) && CFGDSN_delay[30]; // rv 0
  assign CFGDSN_in[31] = (CFGDSN[31] !== 1'bz) && CFGDSN_delay[31]; // rv 0
  assign CFGDSN_in[32] = (CFGDSN[32] !== 1'bz) && CFGDSN_delay[32]; // rv 0
  assign CFGDSN_in[33] = (CFGDSN[33] !== 1'bz) && CFGDSN_delay[33]; // rv 0
  assign CFGDSN_in[34] = (CFGDSN[34] !== 1'bz) && CFGDSN_delay[34]; // rv 0
  assign CFGDSN_in[35] = (CFGDSN[35] !== 1'bz) && CFGDSN_delay[35]; // rv 0
  assign CFGDSN_in[36] = (CFGDSN[36] !== 1'bz) && CFGDSN_delay[36]; // rv 0
  assign CFGDSN_in[37] = (CFGDSN[37] !== 1'bz) && CFGDSN_delay[37]; // rv 0
  assign CFGDSN_in[38] = (CFGDSN[38] !== 1'bz) && CFGDSN_delay[38]; // rv 0
  assign CFGDSN_in[39] = (CFGDSN[39] !== 1'bz) && CFGDSN_delay[39]; // rv 0
  assign CFGDSN_in[3] = (CFGDSN[3] !== 1'bz) && CFGDSN_delay[3]; // rv 0
  assign CFGDSN_in[40] = (CFGDSN[40] !== 1'bz) && CFGDSN_delay[40]; // rv 0
  assign CFGDSN_in[41] = (CFGDSN[41] !== 1'bz) && CFGDSN_delay[41]; // rv 0
  assign CFGDSN_in[42] = (CFGDSN[42] !== 1'bz) && CFGDSN_delay[42]; // rv 0
  assign CFGDSN_in[43] = (CFGDSN[43] !== 1'bz) && CFGDSN_delay[43]; // rv 0
  assign CFGDSN_in[44] = (CFGDSN[44] !== 1'bz) && CFGDSN_delay[44]; // rv 0
  assign CFGDSN_in[45] = (CFGDSN[45] !== 1'bz) && CFGDSN_delay[45]; // rv 0
  assign CFGDSN_in[46] = (CFGDSN[46] !== 1'bz) && CFGDSN_delay[46]; // rv 0
  assign CFGDSN_in[47] = (CFGDSN[47] !== 1'bz) && CFGDSN_delay[47]; // rv 0
  assign CFGDSN_in[48] = (CFGDSN[48] !== 1'bz) && CFGDSN_delay[48]; // rv 0
  assign CFGDSN_in[49] = (CFGDSN[49] !== 1'bz) && CFGDSN_delay[49]; // rv 0
  assign CFGDSN_in[4] = (CFGDSN[4] !== 1'bz) && CFGDSN_delay[4]; // rv 0
  assign CFGDSN_in[50] = (CFGDSN[50] !== 1'bz) && CFGDSN_delay[50]; // rv 0
  assign CFGDSN_in[51] = (CFGDSN[51] !== 1'bz) && CFGDSN_delay[51]; // rv 0
  assign CFGDSN_in[52] = (CFGDSN[52] !== 1'bz) && CFGDSN_delay[52]; // rv 0
  assign CFGDSN_in[53] = (CFGDSN[53] !== 1'bz) && CFGDSN_delay[53]; // rv 0
  assign CFGDSN_in[54] = (CFGDSN[54] !== 1'bz) && CFGDSN_delay[54]; // rv 0
  assign CFGDSN_in[55] = (CFGDSN[55] !== 1'bz) && CFGDSN_delay[55]; // rv 0
  assign CFGDSN_in[56] = (CFGDSN[56] !== 1'bz) && CFGDSN_delay[56]; // rv 0
  assign CFGDSN_in[57] = (CFGDSN[57] !== 1'bz) && CFGDSN_delay[57]; // rv 0
  assign CFGDSN_in[58] = (CFGDSN[58] !== 1'bz) && CFGDSN_delay[58]; // rv 0
  assign CFGDSN_in[59] = (CFGDSN[59] !== 1'bz) && CFGDSN_delay[59]; // rv 0
  assign CFGDSN_in[5] = (CFGDSN[5] !== 1'bz) && CFGDSN_delay[5]; // rv 0
  assign CFGDSN_in[60] = (CFGDSN[60] !== 1'bz) && CFGDSN_delay[60]; // rv 0
  assign CFGDSN_in[61] = (CFGDSN[61] !== 1'bz) && CFGDSN_delay[61]; // rv 0
  assign CFGDSN_in[62] = (CFGDSN[62] !== 1'bz) && CFGDSN_delay[62]; // rv 0
  assign CFGDSN_in[63] = (CFGDSN[63] !== 1'bz) && CFGDSN_delay[63]; // rv 0
  assign CFGDSN_in[6] = (CFGDSN[6] !== 1'bz) && CFGDSN_delay[6]; // rv 0
  assign CFGDSN_in[7] = (CFGDSN[7] !== 1'bz) && CFGDSN_delay[7]; // rv 0
  assign CFGDSN_in[8] = (CFGDSN[8] !== 1'bz) && CFGDSN_delay[8]; // rv 0
  assign CFGDSN_in[9] = (CFGDSN[9] !== 1'bz) && CFGDSN_delay[9]; // rv 0
  assign CFGDSPORTNUMBER_in[0] = (CFGDSPORTNUMBER[0] !== 1'bz) && CFGDSPORTNUMBER_delay[0]; // rv 0
  assign CFGDSPORTNUMBER_in[1] = (CFGDSPORTNUMBER[1] !== 1'bz) && CFGDSPORTNUMBER_delay[1]; // rv 0
  assign CFGDSPORTNUMBER_in[2] = (CFGDSPORTNUMBER[2] !== 1'bz) && CFGDSPORTNUMBER_delay[2]; // rv 0
  assign CFGDSPORTNUMBER_in[3] = (CFGDSPORTNUMBER[3] !== 1'bz) && CFGDSPORTNUMBER_delay[3]; // rv 0
  assign CFGDSPORTNUMBER_in[4] = (CFGDSPORTNUMBER[4] !== 1'bz) && CFGDSPORTNUMBER_delay[4]; // rv 0
  assign CFGDSPORTNUMBER_in[5] = (CFGDSPORTNUMBER[5] !== 1'bz) && CFGDSPORTNUMBER_delay[5]; // rv 0
  assign CFGDSPORTNUMBER_in[6] = (CFGDSPORTNUMBER[6] !== 1'bz) && CFGDSPORTNUMBER_delay[6]; // rv 0
  assign CFGDSPORTNUMBER_in[7] = (CFGDSPORTNUMBER[7] !== 1'bz) && CFGDSPORTNUMBER_delay[7]; // rv 0
  assign CFGERRCORIN_in = (CFGERRCORIN !== 1'bz) && CFGERRCORIN_delay; // rv 0
  assign CFGERRUNCORIN_in = (CFGERRUNCORIN !== 1'bz) && CFGERRUNCORIN_delay; // rv 0
  assign CFGEXTREADDATAVALID_in = (CFGEXTREADDATAVALID !== 1'bz) && CFGEXTREADDATAVALID_delay; // rv 0
  assign CFGEXTREADDATA_in[0] = (CFGEXTREADDATA[0] !== 1'bz) && CFGEXTREADDATA_delay[0]; // rv 0
  assign CFGEXTREADDATA_in[10] = (CFGEXTREADDATA[10] !== 1'bz) && CFGEXTREADDATA_delay[10]; // rv 0
  assign CFGEXTREADDATA_in[11] = (CFGEXTREADDATA[11] !== 1'bz) && CFGEXTREADDATA_delay[11]; // rv 0
  assign CFGEXTREADDATA_in[12] = (CFGEXTREADDATA[12] !== 1'bz) && CFGEXTREADDATA_delay[12]; // rv 0
  assign CFGEXTREADDATA_in[13] = (CFGEXTREADDATA[13] !== 1'bz) && CFGEXTREADDATA_delay[13]; // rv 0
  assign CFGEXTREADDATA_in[14] = (CFGEXTREADDATA[14] !== 1'bz) && CFGEXTREADDATA_delay[14]; // rv 0
  assign CFGEXTREADDATA_in[15] = (CFGEXTREADDATA[15] !== 1'bz) && CFGEXTREADDATA_delay[15]; // rv 0
  assign CFGEXTREADDATA_in[16] = (CFGEXTREADDATA[16] !== 1'bz) && CFGEXTREADDATA_delay[16]; // rv 0
  assign CFGEXTREADDATA_in[17] = (CFGEXTREADDATA[17] !== 1'bz) && CFGEXTREADDATA_delay[17]; // rv 0
  assign CFGEXTREADDATA_in[18] = (CFGEXTREADDATA[18] !== 1'bz) && CFGEXTREADDATA_delay[18]; // rv 0
  assign CFGEXTREADDATA_in[19] = (CFGEXTREADDATA[19] !== 1'bz) && CFGEXTREADDATA_delay[19]; // rv 0
  assign CFGEXTREADDATA_in[1] = (CFGEXTREADDATA[1] !== 1'bz) && CFGEXTREADDATA_delay[1]; // rv 0
  assign CFGEXTREADDATA_in[20] = (CFGEXTREADDATA[20] !== 1'bz) && CFGEXTREADDATA_delay[20]; // rv 0
  assign CFGEXTREADDATA_in[21] = (CFGEXTREADDATA[21] !== 1'bz) && CFGEXTREADDATA_delay[21]; // rv 0
  assign CFGEXTREADDATA_in[22] = (CFGEXTREADDATA[22] !== 1'bz) && CFGEXTREADDATA_delay[22]; // rv 0
  assign CFGEXTREADDATA_in[23] = (CFGEXTREADDATA[23] !== 1'bz) && CFGEXTREADDATA_delay[23]; // rv 0
  assign CFGEXTREADDATA_in[24] = (CFGEXTREADDATA[24] !== 1'bz) && CFGEXTREADDATA_delay[24]; // rv 0
  assign CFGEXTREADDATA_in[25] = (CFGEXTREADDATA[25] !== 1'bz) && CFGEXTREADDATA_delay[25]; // rv 0
  assign CFGEXTREADDATA_in[26] = (CFGEXTREADDATA[26] !== 1'bz) && CFGEXTREADDATA_delay[26]; // rv 0
  assign CFGEXTREADDATA_in[27] = (CFGEXTREADDATA[27] !== 1'bz) && CFGEXTREADDATA_delay[27]; // rv 0
  assign CFGEXTREADDATA_in[28] = (CFGEXTREADDATA[28] !== 1'bz) && CFGEXTREADDATA_delay[28]; // rv 0
  assign CFGEXTREADDATA_in[29] = (CFGEXTREADDATA[29] !== 1'bz) && CFGEXTREADDATA_delay[29]; // rv 0
  assign CFGEXTREADDATA_in[2] = (CFGEXTREADDATA[2] !== 1'bz) && CFGEXTREADDATA_delay[2]; // rv 0
  assign CFGEXTREADDATA_in[30] = (CFGEXTREADDATA[30] !== 1'bz) && CFGEXTREADDATA_delay[30]; // rv 0
  assign CFGEXTREADDATA_in[31] = (CFGEXTREADDATA[31] !== 1'bz) && CFGEXTREADDATA_delay[31]; // rv 0
  assign CFGEXTREADDATA_in[3] = (CFGEXTREADDATA[3] !== 1'bz) && CFGEXTREADDATA_delay[3]; // rv 0
  assign CFGEXTREADDATA_in[4] = (CFGEXTREADDATA[4] !== 1'bz) && CFGEXTREADDATA_delay[4]; // rv 0
  assign CFGEXTREADDATA_in[5] = (CFGEXTREADDATA[5] !== 1'bz) && CFGEXTREADDATA_delay[5]; // rv 0
  assign CFGEXTREADDATA_in[6] = (CFGEXTREADDATA[6] !== 1'bz) && CFGEXTREADDATA_delay[6]; // rv 0
  assign CFGEXTREADDATA_in[7] = (CFGEXTREADDATA[7] !== 1'bz) && CFGEXTREADDATA_delay[7]; // rv 0
  assign CFGEXTREADDATA_in[8] = (CFGEXTREADDATA[8] !== 1'bz) && CFGEXTREADDATA_delay[8]; // rv 0
  assign CFGEXTREADDATA_in[9] = (CFGEXTREADDATA[9] !== 1'bz) && CFGEXTREADDATA_delay[9]; // rv 0
  assign CFGFCSEL_in[0] = (CFGFCSEL[0] !== 1'bz) && CFGFCSEL_delay[0]; // rv 0
  assign CFGFCSEL_in[1] = (CFGFCSEL[1] !== 1'bz) && CFGFCSEL_delay[1]; // rv 0
  assign CFGFCSEL_in[2] = (CFGFCSEL[2] !== 1'bz) && CFGFCSEL_delay[2]; // rv 0
  assign CFGFLRDONE_in[0] = (CFGFLRDONE[0] !== 1'bz) && CFGFLRDONE_delay[0]; // rv 0
  assign CFGFLRDONE_in[1] = (CFGFLRDONE[1] !== 1'bz) && CFGFLRDONE_delay[1]; // rv 0
  assign CFGFLRDONE_in[2] = (CFGFLRDONE[2] !== 1'bz) && CFGFLRDONE_delay[2]; // rv 0
  assign CFGFLRDONE_in[3] = (CFGFLRDONE[3] !== 1'bz) && CFGFLRDONE_delay[3]; // rv 0
  assign CFGHOTRESETIN_in = (CFGHOTRESETIN !== 1'bz) && CFGHOTRESETIN_delay; // rv 0
  assign CFGINTERRUPTINT_in[0] = (CFGINTERRUPTINT[0] !== 1'bz) && CFGINTERRUPTINT_delay[0]; // rv 0
  assign CFGINTERRUPTINT_in[1] = (CFGINTERRUPTINT[1] !== 1'bz) && CFGINTERRUPTINT_delay[1]; // rv 0
  assign CFGINTERRUPTINT_in[2] = (CFGINTERRUPTINT[2] !== 1'bz) && CFGINTERRUPTINT_delay[2]; // rv 0
  assign CFGINTERRUPTINT_in[3] = (CFGINTERRUPTINT[3] !== 1'bz) && CFGINTERRUPTINT_delay[3]; // rv 0
  assign CFGINTERRUPTMSIATTR_in[0] = (CFGINTERRUPTMSIATTR[0] !== 1'bz) && CFGINTERRUPTMSIATTR_delay[0]; // rv 0
  assign CFGINTERRUPTMSIATTR_in[1] = (CFGINTERRUPTMSIATTR[1] !== 1'bz) && CFGINTERRUPTMSIATTR_delay[1]; // rv 0
  assign CFGINTERRUPTMSIATTR_in[2] = (CFGINTERRUPTMSIATTR[2] !== 1'bz) && CFGINTERRUPTMSIATTR_delay[2]; // rv 0
  assign CFGINTERRUPTMSIFUNCTIONNUMBER_in[0] = (CFGINTERRUPTMSIFUNCTIONNUMBER[0] !== 1'bz) && CFGINTERRUPTMSIFUNCTIONNUMBER_delay[0]; // rv 0
  assign CFGINTERRUPTMSIFUNCTIONNUMBER_in[1] = (CFGINTERRUPTMSIFUNCTIONNUMBER[1] !== 1'bz) && CFGINTERRUPTMSIFUNCTIONNUMBER_delay[1]; // rv 0
  assign CFGINTERRUPTMSIFUNCTIONNUMBER_in[2] = (CFGINTERRUPTMSIFUNCTIONNUMBER[2] !== 1'bz) && CFGINTERRUPTMSIFUNCTIONNUMBER_delay[2]; // rv 0
  assign CFGINTERRUPTMSIFUNCTIONNUMBER_in[3] = (CFGINTERRUPTMSIFUNCTIONNUMBER[3] !== 1'bz) && CFGINTERRUPTMSIFUNCTIONNUMBER_delay[3]; // rv 0
  assign CFGINTERRUPTMSIINT_in[0] = (CFGINTERRUPTMSIINT[0] !== 1'bz) && CFGINTERRUPTMSIINT_delay[0]; // rv 0
  assign CFGINTERRUPTMSIINT_in[10] = (CFGINTERRUPTMSIINT[10] !== 1'bz) && CFGINTERRUPTMSIINT_delay[10]; // rv 0
  assign CFGINTERRUPTMSIINT_in[11] = (CFGINTERRUPTMSIINT[11] !== 1'bz) && CFGINTERRUPTMSIINT_delay[11]; // rv 0
  assign CFGINTERRUPTMSIINT_in[12] = (CFGINTERRUPTMSIINT[12] !== 1'bz) && CFGINTERRUPTMSIINT_delay[12]; // rv 0
  assign CFGINTERRUPTMSIINT_in[13] = (CFGINTERRUPTMSIINT[13] !== 1'bz) && CFGINTERRUPTMSIINT_delay[13]; // rv 0
  assign CFGINTERRUPTMSIINT_in[14] = (CFGINTERRUPTMSIINT[14] !== 1'bz) && CFGINTERRUPTMSIINT_delay[14]; // rv 0
  assign CFGINTERRUPTMSIINT_in[15] = (CFGINTERRUPTMSIINT[15] !== 1'bz) && CFGINTERRUPTMSIINT_delay[15]; // rv 0
  assign CFGINTERRUPTMSIINT_in[16] = (CFGINTERRUPTMSIINT[16] !== 1'bz) && CFGINTERRUPTMSIINT_delay[16]; // rv 0
  assign CFGINTERRUPTMSIINT_in[17] = (CFGINTERRUPTMSIINT[17] !== 1'bz) && CFGINTERRUPTMSIINT_delay[17]; // rv 0
  assign CFGINTERRUPTMSIINT_in[18] = (CFGINTERRUPTMSIINT[18] !== 1'bz) && CFGINTERRUPTMSIINT_delay[18]; // rv 0
  assign CFGINTERRUPTMSIINT_in[19] = (CFGINTERRUPTMSIINT[19] !== 1'bz) && CFGINTERRUPTMSIINT_delay[19]; // rv 0
  assign CFGINTERRUPTMSIINT_in[1] = (CFGINTERRUPTMSIINT[1] !== 1'bz) && CFGINTERRUPTMSIINT_delay[1]; // rv 0
  assign CFGINTERRUPTMSIINT_in[20] = (CFGINTERRUPTMSIINT[20] !== 1'bz) && CFGINTERRUPTMSIINT_delay[20]; // rv 0
  assign CFGINTERRUPTMSIINT_in[21] = (CFGINTERRUPTMSIINT[21] !== 1'bz) && CFGINTERRUPTMSIINT_delay[21]; // rv 0
  assign CFGINTERRUPTMSIINT_in[22] = (CFGINTERRUPTMSIINT[22] !== 1'bz) && CFGINTERRUPTMSIINT_delay[22]; // rv 0
  assign CFGINTERRUPTMSIINT_in[23] = (CFGINTERRUPTMSIINT[23] !== 1'bz) && CFGINTERRUPTMSIINT_delay[23]; // rv 0
  assign CFGINTERRUPTMSIINT_in[24] = (CFGINTERRUPTMSIINT[24] !== 1'bz) && CFGINTERRUPTMSIINT_delay[24]; // rv 0
  assign CFGINTERRUPTMSIINT_in[25] = (CFGINTERRUPTMSIINT[25] !== 1'bz) && CFGINTERRUPTMSIINT_delay[25]; // rv 0
  assign CFGINTERRUPTMSIINT_in[26] = (CFGINTERRUPTMSIINT[26] !== 1'bz) && CFGINTERRUPTMSIINT_delay[26]; // rv 0
  assign CFGINTERRUPTMSIINT_in[27] = (CFGINTERRUPTMSIINT[27] !== 1'bz) && CFGINTERRUPTMSIINT_delay[27]; // rv 0
  assign CFGINTERRUPTMSIINT_in[28] = (CFGINTERRUPTMSIINT[28] !== 1'bz) && CFGINTERRUPTMSIINT_delay[28]; // rv 0
  assign CFGINTERRUPTMSIINT_in[29] = (CFGINTERRUPTMSIINT[29] !== 1'bz) && CFGINTERRUPTMSIINT_delay[29]; // rv 0
  assign CFGINTERRUPTMSIINT_in[2] = (CFGINTERRUPTMSIINT[2] !== 1'bz) && CFGINTERRUPTMSIINT_delay[2]; // rv 0
  assign CFGINTERRUPTMSIINT_in[30] = (CFGINTERRUPTMSIINT[30] !== 1'bz) && CFGINTERRUPTMSIINT_delay[30]; // rv 0
  assign CFGINTERRUPTMSIINT_in[31] = (CFGINTERRUPTMSIINT[31] !== 1'bz) && CFGINTERRUPTMSIINT_delay[31]; // rv 0
  assign CFGINTERRUPTMSIINT_in[3] = (CFGINTERRUPTMSIINT[3] !== 1'bz) && CFGINTERRUPTMSIINT_delay[3]; // rv 0
  assign CFGINTERRUPTMSIINT_in[4] = (CFGINTERRUPTMSIINT[4] !== 1'bz) && CFGINTERRUPTMSIINT_delay[4]; // rv 0
  assign CFGINTERRUPTMSIINT_in[5] = (CFGINTERRUPTMSIINT[5] !== 1'bz) && CFGINTERRUPTMSIINT_delay[5]; // rv 0
  assign CFGINTERRUPTMSIINT_in[6] = (CFGINTERRUPTMSIINT[6] !== 1'bz) && CFGINTERRUPTMSIINT_delay[6]; // rv 0
  assign CFGINTERRUPTMSIINT_in[7] = (CFGINTERRUPTMSIINT[7] !== 1'bz) && CFGINTERRUPTMSIINT_delay[7]; // rv 0
  assign CFGINTERRUPTMSIINT_in[8] = (CFGINTERRUPTMSIINT[8] !== 1'bz) && CFGINTERRUPTMSIINT_delay[8]; // rv 0
  assign CFGINTERRUPTMSIINT_in[9] = (CFGINTERRUPTMSIINT[9] !== 1'bz) && CFGINTERRUPTMSIINT_delay[9]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUSDATAENABLE_in = (CFGINTERRUPTMSIPENDINGSTATUSDATAENABLE !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUSDATAENABLE_delay; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM_in[0] = (CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM[0] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM_delay[0]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM_in[1] = (CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM[1] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM_delay[1]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM_in[2] = (CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM[2] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM_delay[2]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM_in[3] = (CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM[3] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM_delay[3]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[0] = (CFGINTERRUPTMSIPENDINGSTATUS[0] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[0]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[10] = (CFGINTERRUPTMSIPENDINGSTATUS[10] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[10]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[11] = (CFGINTERRUPTMSIPENDINGSTATUS[11] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[11]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[12] = (CFGINTERRUPTMSIPENDINGSTATUS[12] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[12]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[13] = (CFGINTERRUPTMSIPENDINGSTATUS[13] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[13]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[14] = (CFGINTERRUPTMSIPENDINGSTATUS[14] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[14]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[15] = (CFGINTERRUPTMSIPENDINGSTATUS[15] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[15]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[16] = (CFGINTERRUPTMSIPENDINGSTATUS[16] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[16]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[17] = (CFGINTERRUPTMSIPENDINGSTATUS[17] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[17]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[18] = (CFGINTERRUPTMSIPENDINGSTATUS[18] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[18]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[19] = (CFGINTERRUPTMSIPENDINGSTATUS[19] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[19]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[1] = (CFGINTERRUPTMSIPENDINGSTATUS[1] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[1]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[20] = (CFGINTERRUPTMSIPENDINGSTATUS[20] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[20]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[21] = (CFGINTERRUPTMSIPENDINGSTATUS[21] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[21]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[22] = (CFGINTERRUPTMSIPENDINGSTATUS[22] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[22]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[23] = (CFGINTERRUPTMSIPENDINGSTATUS[23] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[23]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[24] = (CFGINTERRUPTMSIPENDINGSTATUS[24] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[24]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[25] = (CFGINTERRUPTMSIPENDINGSTATUS[25] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[25]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[26] = (CFGINTERRUPTMSIPENDINGSTATUS[26] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[26]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[27] = (CFGINTERRUPTMSIPENDINGSTATUS[27] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[27]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[28] = (CFGINTERRUPTMSIPENDINGSTATUS[28] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[28]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[29] = (CFGINTERRUPTMSIPENDINGSTATUS[29] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[29]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[2] = (CFGINTERRUPTMSIPENDINGSTATUS[2] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[2]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[30] = (CFGINTERRUPTMSIPENDINGSTATUS[30] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[30]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[31] = (CFGINTERRUPTMSIPENDINGSTATUS[31] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[31]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[3] = (CFGINTERRUPTMSIPENDINGSTATUS[3] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[3]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[4] = (CFGINTERRUPTMSIPENDINGSTATUS[4] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[4]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[5] = (CFGINTERRUPTMSIPENDINGSTATUS[5] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[5]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[6] = (CFGINTERRUPTMSIPENDINGSTATUS[6] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[6]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[7] = (CFGINTERRUPTMSIPENDINGSTATUS[7] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[7]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[8] = (CFGINTERRUPTMSIPENDINGSTATUS[8] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[8]; // rv 0
  assign CFGINTERRUPTMSIPENDINGSTATUS_in[9] = (CFGINTERRUPTMSIPENDINGSTATUS[9] !== 1'bz) && CFGINTERRUPTMSIPENDINGSTATUS_delay[9]; // rv 0
  assign CFGINTERRUPTMSISELECT_in[0] = (CFGINTERRUPTMSISELECT[0] !== 1'bz) && CFGINTERRUPTMSISELECT_delay[0]; // rv 0
  assign CFGINTERRUPTMSISELECT_in[1] = (CFGINTERRUPTMSISELECT[1] !== 1'bz) && CFGINTERRUPTMSISELECT_delay[1]; // rv 0
  assign CFGINTERRUPTMSISELECT_in[2] = (CFGINTERRUPTMSISELECT[2] !== 1'bz) && CFGINTERRUPTMSISELECT_delay[2]; // rv 0
  assign CFGINTERRUPTMSISELECT_in[3] = (CFGINTERRUPTMSISELECT[3] !== 1'bz) && CFGINTERRUPTMSISELECT_delay[3]; // rv 0
  assign CFGINTERRUPTMSITPHPRESENT_in = (CFGINTERRUPTMSITPHPRESENT !== 1'bz) && CFGINTERRUPTMSITPHPRESENT_delay; // rv 0
  assign CFGINTERRUPTMSITPHSTTAG_in[0] = (CFGINTERRUPTMSITPHSTTAG[0] !== 1'bz) && CFGINTERRUPTMSITPHSTTAG_delay[0]; // rv 0
  assign CFGINTERRUPTMSITPHSTTAG_in[1] = (CFGINTERRUPTMSITPHSTTAG[1] !== 1'bz) && CFGINTERRUPTMSITPHSTTAG_delay[1]; // rv 0
  assign CFGINTERRUPTMSITPHSTTAG_in[2] = (CFGINTERRUPTMSITPHSTTAG[2] !== 1'bz) && CFGINTERRUPTMSITPHSTTAG_delay[2]; // rv 0
  assign CFGINTERRUPTMSITPHSTTAG_in[3] = (CFGINTERRUPTMSITPHSTTAG[3] !== 1'bz) && CFGINTERRUPTMSITPHSTTAG_delay[3]; // rv 0
  assign CFGINTERRUPTMSITPHSTTAG_in[4] = (CFGINTERRUPTMSITPHSTTAG[4] !== 1'bz) && CFGINTERRUPTMSITPHSTTAG_delay[4]; // rv 0
  assign CFGINTERRUPTMSITPHSTTAG_in[5] = (CFGINTERRUPTMSITPHSTTAG[5] !== 1'bz) && CFGINTERRUPTMSITPHSTTAG_delay[5]; // rv 0
  assign CFGINTERRUPTMSITPHSTTAG_in[6] = (CFGINTERRUPTMSITPHSTTAG[6] !== 1'bz) && CFGINTERRUPTMSITPHSTTAG_delay[6]; // rv 0
  assign CFGINTERRUPTMSITPHSTTAG_in[7] = (CFGINTERRUPTMSITPHSTTAG[7] !== 1'bz) && CFGINTERRUPTMSITPHSTTAG_delay[7]; // rv 0
  assign CFGINTERRUPTMSITPHSTTAG_in[8] = (CFGINTERRUPTMSITPHSTTAG[8] !== 1'bz) && CFGINTERRUPTMSITPHSTTAG_delay[8]; // rv 0
  assign CFGINTERRUPTMSITPHTYPE_in[0] = (CFGINTERRUPTMSITPHTYPE[0] !== 1'bz) && CFGINTERRUPTMSITPHTYPE_delay[0]; // rv 0
  assign CFGINTERRUPTMSITPHTYPE_in[1] = (CFGINTERRUPTMSITPHTYPE[1] !== 1'bz) && CFGINTERRUPTMSITPHTYPE_delay[1]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[0] = (CFGINTERRUPTMSIXADDRESS[0] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[0]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[10] = (CFGINTERRUPTMSIXADDRESS[10] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[10]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[11] = (CFGINTERRUPTMSIXADDRESS[11] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[11]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[12] = (CFGINTERRUPTMSIXADDRESS[12] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[12]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[13] = (CFGINTERRUPTMSIXADDRESS[13] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[13]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[14] = (CFGINTERRUPTMSIXADDRESS[14] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[14]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[15] = (CFGINTERRUPTMSIXADDRESS[15] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[15]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[16] = (CFGINTERRUPTMSIXADDRESS[16] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[16]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[17] = (CFGINTERRUPTMSIXADDRESS[17] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[17]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[18] = (CFGINTERRUPTMSIXADDRESS[18] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[18]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[19] = (CFGINTERRUPTMSIXADDRESS[19] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[19]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[1] = (CFGINTERRUPTMSIXADDRESS[1] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[1]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[20] = (CFGINTERRUPTMSIXADDRESS[20] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[20]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[21] = (CFGINTERRUPTMSIXADDRESS[21] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[21]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[22] = (CFGINTERRUPTMSIXADDRESS[22] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[22]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[23] = (CFGINTERRUPTMSIXADDRESS[23] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[23]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[24] = (CFGINTERRUPTMSIXADDRESS[24] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[24]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[25] = (CFGINTERRUPTMSIXADDRESS[25] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[25]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[26] = (CFGINTERRUPTMSIXADDRESS[26] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[26]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[27] = (CFGINTERRUPTMSIXADDRESS[27] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[27]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[28] = (CFGINTERRUPTMSIXADDRESS[28] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[28]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[29] = (CFGINTERRUPTMSIXADDRESS[29] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[29]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[2] = (CFGINTERRUPTMSIXADDRESS[2] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[2]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[30] = (CFGINTERRUPTMSIXADDRESS[30] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[30]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[31] = (CFGINTERRUPTMSIXADDRESS[31] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[31]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[32] = (CFGINTERRUPTMSIXADDRESS[32] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[32]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[33] = (CFGINTERRUPTMSIXADDRESS[33] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[33]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[34] = (CFGINTERRUPTMSIXADDRESS[34] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[34]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[35] = (CFGINTERRUPTMSIXADDRESS[35] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[35]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[36] = (CFGINTERRUPTMSIXADDRESS[36] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[36]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[37] = (CFGINTERRUPTMSIXADDRESS[37] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[37]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[38] = (CFGINTERRUPTMSIXADDRESS[38] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[38]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[39] = (CFGINTERRUPTMSIXADDRESS[39] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[39]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[3] = (CFGINTERRUPTMSIXADDRESS[3] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[3]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[40] = (CFGINTERRUPTMSIXADDRESS[40] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[40]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[41] = (CFGINTERRUPTMSIXADDRESS[41] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[41]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[42] = (CFGINTERRUPTMSIXADDRESS[42] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[42]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[43] = (CFGINTERRUPTMSIXADDRESS[43] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[43]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[44] = (CFGINTERRUPTMSIXADDRESS[44] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[44]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[45] = (CFGINTERRUPTMSIXADDRESS[45] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[45]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[46] = (CFGINTERRUPTMSIXADDRESS[46] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[46]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[47] = (CFGINTERRUPTMSIXADDRESS[47] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[47]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[48] = (CFGINTERRUPTMSIXADDRESS[48] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[48]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[49] = (CFGINTERRUPTMSIXADDRESS[49] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[49]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[4] = (CFGINTERRUPTMSIXADDRESS[4] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[4]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[50] = (CFGINTERRUPTMSIXADDRESS[50] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[50]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[51] = (CFGINTERRUPTMSIXADDRESS[51] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[51]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[52] = (CFGINTERRUPTMSIXADDRESS[52] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[52]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[53] = (CFGINTERRUPTMSIXADDRESS[53] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[53]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[54] = (CFGINTERRUPTMSIXADDRESS[54] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[54]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[55] = (CFGINTERRUPTMSIXADDRESS[55] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[55]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[56] = (CFGINTERRUPTMSIXADDRESS[56] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[56]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[57] = (CFGINTERRUPTMSIXADDRESS[57] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[57]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[58] = (CFGINTERRUPTMSIXADDRESS[58] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[58]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[59] = (CFGINTERRUPTMSIXADDRESS[59] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[59]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[5] = (CFGINTERRUPTMSIXADDRESS[5] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[5]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[60] = (CFGINTERRUPTMSIXADDRESS[60] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[60]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[61] = (CFGINTERRUPTMSIXADDRESS[61] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[61]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[62] = (CFGINTERRUPTMSIXADDRESS[62] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[62]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[63] = (CFGINTERRUPTMSIXADDRESS[63] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[63]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[6] = (CFGINTERRUPTMSIXADDRESS[6] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[6]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[7] = (CFGINTERRUPTMSIXADDRESS[7] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[7]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[8] = (CFGINTERRUPTMSIXADDRESS[8] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[8]; // rv 0
  assign CFGINTERRUPTMSIXADDRESS_in[9] = (CFGINTERRUPTMSIXADDRESS[9] !== 1'bz) && CFGINTERRUPTMSIXADDRESS_delay[9]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[0] = (CFGINTERRUPTMSIXDATA[0] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[0]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[10] = (CFGINTERRUPTMSIXDATA[10] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[10]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[11] = (CFGINTERRUPTMSIXDATA[11] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[11]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[12] = (CFGINTERRUPTMSIXDATA[12] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[12]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[13] = (CFGINTERRUPTMSIXDATA[13] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[13]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[14] = (CFGINTERRUPTMSIXDATA[14] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[14]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[15] = (CFGINTERRUPTMSIXDATA[15] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[15]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[16] = (CFGINTERRUPTMSIXDATA[16] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[16]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[17] = (CFGINTERRUPTMSIXDATA[17] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[17]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[18] = (CFGINTERRUPTMSIXDATA[18] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[18]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[19] = (CFGINTERRUPTMSIXDATA[19] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[19]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[1] = (CFGINTERRUPTMSIXDATA[1] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[1]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[20] = (CFGINTERRUPTMSIXDATA[20] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[20]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[21] = (CFGINTERRUPTMSIXDATA[21] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[21]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[22] = (CFGINTERRUPTMSIXDATA[22] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[22]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[23] = (CFGINTERRUPTMSIXDATA[23] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[23]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[24] = (CFGINTERRUPTMSIXDATA[24] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[24]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[25] = (CFGINTERRUPTMSIXDATA[25] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[25]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[26] = (CFGINTERRUPTMSIXDATA[26] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[26]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[27] = (CFGINTERRUPTMSIXDATA[27] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[27]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[28] = (CFGINTERRUPTMSIXDATA[28] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[28]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[29] = (CFGINTERRUPTMSIXDATA[29] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[29]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[2] = (CFGINTERRUPTMSIXDATA[2] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[2]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[30] = (CFGINTERRUPTMSIXDATA[30] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[30]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[31] = (CFGINTERRUPTMSIXDATA[31] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[31]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[3] = (CFGINTERRUPTMSIXDATA[3] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[3]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[4] = (CFGINTERRUPTMSIXDATA[4] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[4]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[5] = (CFGINTERRUPTMSIXDATA[5] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[5]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[6] = (CFGINTERRUPTMSIXDATA[6] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[6]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[7] = (CFGINTERRUPTMSIXDATA[7] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[7]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[8] = (CFGINTERRUPTMSIXDATA[8] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[8]; // rv 0
  assign CFGINTERRUPTMSIXDATA_in[9] = (CFGINTERRUPTMSIXDATA[9] !== 1'bz) && CFGINTERRUPTMSIXDATA_delay[9]; // rv 0
  assign CFGINTERRUPTMSIXINT_in = (CFGINTERRUPTMSIXINT !== 1'bz) && CFGINTERRUPTMSIXINT_delay; // rv 0
  assign CFGINTERRUPTPENDING_in[0] = (CFGINTERRUPTPENDING[0] !== 1'bz) && CFGINTERRUPTPENDING_delay[0]; // rv 0
  assign CFGINTERRUPTPENDING_in[1] = (CFGINTERRUPTPENDING[1] !== 1'bz) && CFGINTERRUPTPENDING_delay[1]; // rv 0
  assign CFGINTERRUPTPENDING_in[2] = (CFGINTERRUPTPENDING[2] !== 1'bz) && CFGINTERRUPTPENDING_delay[2]; // rv 0
  assign CFGINTERRUPTPENDING_in[3] = (CFGINTERRUPTPENDING[3] !== 1'bz) && CFGINTERRUPTPENDING_delay[3]; // rv 0
  assign CFGLINKTRAININGENABLE_in = (CFGLINKTRAININGENABLE === 1'bz) || CFGLINKTRAININGENABLE_delay; // rv 1
  assign CFGMGMTADDR_in[0] = (CFGMGMTADDR[0] !== 1'bz) && CFGMGMTADDR_delay[0]; // rv 0
  assign CFGMGMTADDR_in[10] = (CFGMGMTADDR[10] !== 1'bz) && CFGMGMTADDR_delay[10]; // rv 0
  assign CFGMGMTADDR_in[11] = (CFGMGMTADDR[11] !== 1'bz) && CFGMGMTADDR_delay[11]; // rv 0
  assign CFGMGMTADDR_in[12] = (CFGMGMTADDR[12] !== 1'bz) && CFGMGMTADDR_delay[12]; // rv 0
  assign CFGMGMTADDR_in[13] = (CFGMGMTADDR[13] !== 1'bz) && CFGMGMTADDR_delay[13]; // rv 0
  assign CFGMGMTADDR_in[14] = (CFGMGMTADDR[14] !== 1'bz) && CFGMGMTADDR_delay[14]; // rv 0
  assign CFGMGMTADDR_in[15] = (CFGMGMTADDR[15] !== 1'bz) && CFGMGMTADDR_delay[15]; // rv 0
  assign CFGMGMTADDR_in[16] = (CFGMGMTADDR[16] !== 1'bz) && CFGMGMTADDR_delay[16]; // rv 0
  assign CFGMGMTADDR_in[17] = (CFGMGMTADDR[17] !== 1'bz) && CFGMGMTADDR_delay[17]; // rv 0
  assign CFGMGMTADDR_in[18] = (CFGMGMTADDR[18] !== 1'bz) && CFGMGMTADDR_delay[18]; // rv 0
  assign CFGMGMTADDR_in[1] = (CFGMGMTADDR[1] !== 1'bz) && CFGMGMTADDR_delay[1]; // rv 0
  assign CFGMGMTADDR_in[2] = (CFGMGMTADDR[2] !== 1'bz) && CFGMGMTADDR_delay[2]; // rv 0
  assign CFGMGMTADDR_in[3] = (CFGMGMTADDR[3] !== 1'bz) && CFGMGMTADDR_delay[3]; // rv 0
  assign CFGMGMTADDR_in[4] = (CFGMGMTADDR[4] !== 1'bz) && CFGMGMTADDR_delay[4]; // rv 0
  assign CFGMGMTADDR_in[5] = (CFGMGMTADDR[5] !== 1'bz) && CFGMGMTADDR_delay[5]; // rv 0
  assign CFGMGMTADDR_in[6] = (CFGMGMTADDR[6] !== 1'bz) && CFGMGMTADDR_delay[6]; // rv 0
  assign CFGMGMTADDR_in[7] = (CFGMGMTADDR[7] !== 1'bz) && CFGMGMTADDR_delay[7]; // rv 0
  assign CFGMGMTADDR_in[8] = (CFGMGMTADDR[8] !== 1'bz) && CFGMGMTADDR_delay[8]; // rv 0
  assign CFGMGMTADDR_in[9] = (CFGMGMTADDR[9] !== 1'bz) && CFGMGMTADDR_delay[9]; // rv 0
  assign CFGMGMTBYTEENABLE_in[0] = (CFGMGMTBYTEENABLE[0] !== 1'bz) && CFGMGMTBYTEENABLE_delay[0]; // rv 0
  assign CFGMGMTBYTEENABLE_in[1] = (CFGMGMTBYTEENABLE[1] !== 1'bz) && CFGMGMTBYTEENABLE_delay[1]; // rv 0
  assign CFGMGMTBYTEENABLE_in[2] = (CFGMGMTBYTEENABLE[2] !== 1'bz) && CFGMGMTBYTEENABLE_delay[2]; // rv 0
  assign CFGMGMTBYTEENABLE_in[3] = (CFGMGMTBYTEENABLE[3] !== 1'bz) && CFGMGMTBYTEENABLE_delay[3]; // rv 0
  assign CFGMGMTREAD_in = (CFGMGMTREAD !== 1'bz) && CFGMGMTREAD_delay; // rv 0
  assign CFGMGMTTYPE1CFGREGACCESS_in = (CFGMGMTTYPE1CFGREGACCESS !== 1'bz) && CFGMGMTTYPE1CFGREGACCESS_delay; // rv 0
  assign CFGMGMTWRITEDATA_in[0] = (CFGMGMTWRITEDATA[0] !== 1'bz) && CFGMGMTWRITEDATA_delay[0]; // rv 0
  assign CFGMGMTWRITEDATA_in[10] = (CFGMGMTWRITEDATA[10] !== 1'bz) && CFGMGMTWRITEDATA_delay[10]; // rv 0
  assign CFGMGMTWRITEDATA_in[11] = (CFGMGMTWRITEDATA[11] !== 1'bz) && CFGMGMTWRITEDATA_delay[11]; // rv 0
  assign CFGMGMTWRITEDATA_in[12] = (CFGMGMTWRITEDATA[12] !== 1'bz) && CFGMGMTWRITEDATA_delay[12]; // rv 0
  assign CFGMGMTWRITEDATA_in[13] = (CFGMGMTWRITEDATA[13] !== 1'bz) && CFGMGMTWRITEDATA_delay[13]; // rv 0
  assign CFGMGMTWRITEDATA_in[14] = (CFGMGMTWRITEDATA[14] !== 1'bz) && CFGMGMTWRITEDATA_delay[14]; // rv 0
  assign CFGMGMTWRITEDATA_in[15] = (CFGMGMTWRITEDATA[15] !== 1'bz) && CFGMGMTWRITEDATA_delay[15]; // rv 0
  assign CFGMGMTWRITEDATA_in[16] = (CFGMGMTWRITEDATA[16] !== 1'bz) && CFGMGMTWRITEDATA_delay[16]; // rv 0
  assign CFGMGMTWRITEDATA_in[17] = (CFGMGMTWRITEDATA[17] !== 1'bz) && CFGMGMTWRITEDATA_delay[17]; // rv 0
  assign CFGMGMTWRITEDATA_in[18] = (CFGMGMTWRITEDATA[18] !== 1'bz) && CFGMGMTWRITEDATA_delay[18]; // rv 0
  assign CFGMGMTWRITEDATA_in[19] = (CFGMGMTWRITEDATA[19] !== 1'bz) && CFGMGMTWRITEDATA_delay[19]; // rv 0
  assign CFGMGMTWRITEDATA_in[1] = (CFGMGMTWRITEDATA[1] !== 1'bz) && CFGMGMTWRITEDATA_delay[1]; // rv 0
  assign CFGMGMTWRITEDATA_in[20] = (CFGMGMTWRITEDATA[20] !== 1'bz) && CFGMGMTWRITEDATA_delay[20]; // rv 0
  assign CFGMGMTWRITEDATA_in[21] = (CFGMGMTWRITEDATA[21] !== 1'bz) && CFGMGMTWRITEDATA_delay[21]; // rv 0
  assign CFGMGMTWRITEDATA_in[22] = (CFGMGMTWRITEDATA[22] !== 1'bz) && CFGMGMTWRITEDATA_delay[22]; // rv 0
  assign CFGMGMTWRITEDATA_in[23] = (CFGMGMTWRITEDATA[23] !== 1'bz) && CFGMGMTWRITEDATA_delay[23]; // rv 0
  assign CFGMGMTWRITEDATA_in[24] = (CFGMGMTWRITEDATA[24] !== 1'bz) && CFGMGMTWRITEDATA_delay[24]; // rv 0
  assign CFGMGMTWRITEDATA_in[25] = (CFGMGMTWRITEDATA[25] !== 1'bz) && CFGMGMTWRITEDATA_delay[25]; // rv 0
  assign CFGMGMTWRITEDATA_in[26] = (CFGMGMTWRITEDATA[26] !== 1'bz) && CFGMGMTWRITEDATA_delay[26]; // rv 0
  assign CFGMGMTWRITEDATA_in[27] = (CFGMGMTWRITEDATA[27] !== 1'bz) && CFGMGMTWRITEDATA_delay[27]; // rv 0
  assign CFGMGMTWRITEDATA_in[28] = (CFGMGMTWRITEDATA[28] !== 1'bz) && CFGMGMTWRITEDATA_delay[28]; // rv 0
  assign CFGMGMTWRITEDATA_in[29] = (CFGMGMTWRITEDATA[29] !== 1'bz) && CFGMGMTWRITEDATA_delay[29]; // rv 0
  assign CFGMGMTWRITEDATA_in[2] = (CFGMGMTWRITEDATA[2] !== 1'bz) && CFGMGMTWRITEDATA_delay[2]; // rv 0
  assign CFGMGMTWRITEDATA_in[30] = (CFGMGMTWRITEDATA[30] !== 1'bz) && CFGMGMTWRITEDATA_delay[30]; // rv 0
  assign CFGMGMTWRITEDATA_in[31] = (CFGMGMTWRITEDATA[31] !== 1'bz) && CFGMGMTWRITEDATA_delay[31]; // rv 0
  assign CFGMGMTWRITEDATA_in[3] = (CFGMGMTWRITEDATA[3] !== 1'bz) && CFGMGMTWRITEDATA_delay[3]; // rv 0
  assign CFGMGMTWRITEDATA_in[4] = (CFGMGMTWRITEDATA[4] !== 1'bz) && CFGMGMTWRITEDATA_delay[4]; // rv 0
  assign CFGMGMTWRITEDATA_in[5] = (CFGMGMTWRITEDATA[5] !== 1'bz) && CFGMGMTWRITEDATA_delay[5]; // rv 0
  assign CFGMGMTWRITEDATA_in[6] = (CFGMGMTWRITEDATA[6] !== 1'bz) && CFGMGMTWRITEDATA_delay[6]; // rv 0
  assign CFGMGMTWRITEDATA_in[7] = (CFGMGMTWRITEDATA[7] !== 1'bz) && CFGMGMTWRITEDATA_delay[7]; // rv 0
  assign CFGMGMTWRITEDATA_in[8] = (CFGMGMTWRITEDATA[8] !== 1'bz) && CFGMGMTWRITEDATA_delay[8]; // rv 0
  assign CFGMGMTWRITEDATA_in[9] = (CFGMGMTWRITEDATA[9] !== 1'bz) && CFGMGMTWRITEDATA_delay[9]; // rv 0
  assign CFGMGMTWRITE_in = (CFGMGMTWRITE !== 1'bz) && CFGMGMTWRITE_delay; // rv 0
  assign CFGMSGTRANSMITDATA_in[0] = (CFGMSGTRANSMITDATA[0] !== 1'bz) && CFGMSGTRANSMITDATA_delay[0]; // rv 0
  assign CFGMSGTRANSMITDATA_in[10] = (CFGMSGTRANSMITDATA[10] !== 1'bz) && CFGMSGTRANSMITDATA_delay[10]; // rv 0
  assign CFGMSGTRANSMITDATA_in[11] = (CFGMSGTRANSMITDATA[11] !== 1'bz) && CFGMSGTRANSMITDATA_delay[11]; // rv 0
  assign CFGMSGTRANSMITDATA_in[12] = (CFGMSGTRANSMITDATA[12] !== 1'bz) && CFGMSGTRANSMITDATA_delay[12]; // rv 0
  assign CFGMSGTRANSMITDATA_in[13] = (CFGMSGTRANSMITDATA[13] !== 1'bz) && CFGMSGTRANSMITDATA_delay[13]; // rv 0
  assign CFGMSGTRANSMITDATA_in[14] = (CFGMSGTRANSMITDATA[14] !== 1'bz) && CFGMSGTRANSMITDATA_delay[14]; // rv 0
  assign CFGMSGTRANSMITDATA_in[15] = (CFGMSGTRANSMITDATA[15] !== 1'bz) && CFGMSGTRANSMITDATA_delay[15]; // rv 0
  assign CFGMSGTRANSMITDATA_in[16] = (CFGMSGTRANSMITDATA[16] !== 1'bz) && CFGMSGTRANSMITDATA_delay[16]; // rv 0
  assign CFGMSGTRANSMITDATA_in[17] = (CFGMSGTRANSMITDATA[17] !== 1'bz) && CFGMSGTRANSMITDATA_delay[17]; // rv 0
  assign CFGMSGTRANSMITDATA_in[18] = (CFGMSGTRANSMITDATA[18] !== 1'bz) && CFGMSGTRANSMITDATA_delay[18]; // rv 0
  assign CFGMSGTRANSMITDATA_in[19] = (CFGMSGTRANSMITDATA[19] !== 1'bz) && CFGMSGTRANSMITDATA_delay[19]; // rv 0
  assign CFGMSGTRANSMITDATA_in[1] = (CFGMSGTRANSMITDATA[1] !== 1'bz) && CFGMSGTRANSMITDATA_delay[1]; // rv 0
  assign CFGMSGTRANSMITDATA_in[20] = (CFGMSGTRANSMITDATA[20] !== 1'bz) && CFGMSGTRANSMITDATA_delay[20]; // rv 0
  assign CFGMSGTRANSMITDATA_in[21] = (CFGMSGTRANSMITDATA[21] !== 1'bz) && CFGMSGTRANSMITDATA_delay[21]; // rv 0
  assign CFGMSGTRANSMITDATA_in[22] = (CFGMSGTRANSMITDATA[22] !== 1'bz) && CFGMSGTRANSMITDATA_delay[22]; // rv 0
  assign CFGMSGTRANSMITDATA_in[23] = (CFGMSGTRANSMITDATA[23] !== 1'bz) && CFGMSGTRANSMITDATA_delay[23]; // rv 0
  assign CFGMSGTRANSMITDATA_in[24] = (CFGMSGTRANSMITDATA[24] !== 1'bz) && CFGMSGTRANSMITDATA_delay[24]; // rv 0
  assign CFGMSGTRANSMITDATA_in[25] = (CFGMSGTRANSMITDATA[25] !== 1'bz) && CFGMSGTRANSMITDATA_delay[25]; // rv 0
  assign CFGMSGTRANSMITDATA_in[26] = (CFGMSGTRANSMITDATA[26] !== 1'bz) && CFGMSGTRANSMITDATA_delay[26]; // rv 0
  assign CFGMSGTRANSMITDATA_in[27] = (CFGMSGTRANSMITDATA[27] !== 1'bz) && CFGMSGTRANSMITDATA_delay[27]; // rv 0
  assign CFGMSGTRANSMITDATA_in[28] = (CFGMSGTRANSMITDATA[28] !== 1'bz) && CFGMSGTRANSMITDATA_delay[28]; // rv 0
  assign CFGMSGTRANSMITDATA_in[29] = (CFGMSGTRANSMITDATA[29] !== 1'bz) && CFGMSGTRANSMITDATA_delay[29]; // rv 0
  assign CFGMSGTRANSMITDATA_in[2] = (CFGMSGTRANSMITDATA[2] !== 1'bz) && CFGMSGTRANSMITDATA_delay[2]; // rv 0
  assign CFGMSGTRANSMITDATA_in[30] = (CFGMSGTRANSMITDATA[30] !== 1'bz) && CFGMSGTRANSMITDATA_delay[30]; // rv 0
  assign CFGMSGTRANSMITDATA_in[31] = (CFGMSGTRANSMITDATA[31] !== 1'bz) && CFGMSGTRANSMITDATA_delay[31]; // rv 0
  assign CFGMSGTRANSMITDATA_in[3] = (CFGMSGTRANSMITDATA[3] !== 1'bz) && CFGMSGTRANSMITDATA_delay[3]; // rv 0
  assign CFGMSGTRANSMITDATA_in[4] = (CFGMSGTRANSMITDATA[4] !== 1'bz) && CFGMSGTRANSMITDATA_delay[4]; // rv 0
  assign CFGMSGTRANSMITDATA_in[5] = (CFGMSGTRANSMITDATA[5] !== 1'bz) && CFGMSGTRANSMITDATA_delay[5]; // rv 0
  assign CFGMSGTRANSMITDATA_in[6] = (CFGMSGTRANSMITDATA[6] !== 1'bz) && CFGMSGTRANSMITDATA_delay[6]; // rv 0
  assign CFGMSGTRANSMITDATA_in[7] = (CFGMSGTRANSMITDATA[7] !== 1'bz) && CFGMSGTRANSMITDATA_delay[7]; // rv 0
  assign CFGMSGTRANSMITDATA_in[8] = (CFGMSGTRANSMITDATA[8] !== 1'bz) && CFGMSGTRANSMITDATA_delay[8]; // rv 0
  assign CFGMSGTRANSMITDATA_in[9] = (CFGMSGTRANSMITDATA[9] !== 1'bz) && CFGMSGTRANSMITDATA_delay[9]; // rv 0
  assign CFGMSGTRANSMITTYPE_in[0] = (CFGMSGTRANSMITTYPE[0] !== 1'bz) && CFGMSGTRANSMITTYPE_delay[0]; // rv 0
  assign CFGMSGTRANSMITTYPE_in[1] = (CFGMSGTRANSMITTYPE[1] !== 1'bz) && CFGMSGTRANSMITTYPE_delay[1]; // rv 0
  assign CFGMSGTRANSMITTYPE_in[2] = (CFGMSGTRANSMITTYPE[2] !== 1'bz) && CFGMSGTRANSMITTYPE_delay[2]; // rv 0
  assign CFGMSGTRANSMIT_in = (CFGMSGTRANSMIT !== 1'bz) && CFGMSGTRANSMIT_delay; // rv 0
  assign CFGPERFUNCSTATUSCONTROL_in[0] = (CFGPERFUNCSTATUSCONTROL[0] !== 1'bz) && CFGPERFUNCSTATUSCONTROL_delay[0]; // rv 0
  assign CFGPERFUNCSTATUSCONTROL_in[1] = (CFGPERFUNCSTATUSCONTROL[1] !== 1'bz) && CFGPERFUNCSTATUSCONTROL_delay[1]; // rv 0
  assign CFGPERFUNCSTATUSCONTROL_in[2] = (CFGPERFUNCSTATUSCONTROL[2] !== 1'bz) && CFGPERFUNCSTATUSCONTROL_delay[2]; // rv 0
  assign CFGPERFUNCTIONNUMBER_in[0] = (CFGPERFUNCTIONNUMBER[0] !== 1'bz) && CFGPERFUNCTIONNUMBER_delay[0]; // rv 0
  assign CFGPERFUNCTIONNUMBER_in[1] = (CFGPERFUNCTIONNUMBER[1] !== 1'bz) && CFGPERFUNCTIONNUMBER_delay[1]; // rv 0
  assign CFGPERFUNCTIONNUMBER_in[2] = (CFGPERFUNCTIONNUMBER[2] !== 1'bz) && CFGPERFUNCTIONNUMBER_delay[2]; // rv 0
  assign CFGPERFUNCTIONNUMBER_in[3] = (CFGPERFUNCTIONNUMBER[3] !== 1'bz) && CFGPERFUNCTIONNUMBER_delay[3]; // rv 0
  assign CFGPERFUNCTIONOUTPUTREQUEST_in = (CFGPERFUNCTIONOUTPUTREQUEST !== 1'bz) && CFGPERFUNCTIONOUTPUTREQUEST_delay; // rv 0
  assign CFGPOWERSTATECHANGEACK_in = (CFGPOWERSTATECHANGEACK === 1'bz) || CFGPOWERSTATECHANGEACK_delay; // rv 1
  assign CFGREQPMTRANSITIONL23READY_in = (CFGREQPMTRANSITIONL23READY !== 1'bz) && CFGREQPMTRANSITIONL23READY_delay; // rv 0
  assign CFGREVID_in[0] = (CFGREVID[0] !== 1'bz) && CFGREVID_delay[0]; // rv 0
  assign CFGREVID_in[1] = (CFGREVID[1] !== 1'bz) && CFGREVID_delay[1]; // rv 0
  assign CFGREVID_in[2] = (CFGREVID[2] !== 1'bz) && CFGREVID_delay[2]; // rv 0
  assign CFGREVID_in[3] = (CFGREVID[3] !== 1'bz) && CFGREVID_delay[3]; // rv 0
  assign CFGREVID_in[4] = (CFGREVID[4] !== 1'bz) && CFGREVID_delay[4]; // rv 0
  assign CFGREVID_in[5] = (CFGREVID[5] !== 1'bz) && CFGREVID_delay[5]; // rv 0
  assign CFGREVID_in[6] = (CFGREVID[6] !== 1'bz) && CFGREVID_delay[6]; // rv 0
  assign CFGREVID_in[7] = (CFGREVID[7] !== 1'bz) && CFGREVID_delay[7]; // rv 0
  assign CFGSUBSYSID_in[0] = (CFGSUBSYSID[0] !== 1'bz) && CFGSUBSYSID_delay[0]; // rv 0
  assign CFGSUBSYSID_in[10] = (CFGSUBSYSID[10] !== 1'bz) && CFGSUBSYSID_delay[10]; // rv 0
  assign CFGSUBSYSID_in[11] = (CFGSUBSYSID[11] !== 1'bz) && CFGSUBSYSID_delay[11]; // rv 0
  assign CFGSUBSYSID_in[12] = (CFGSUBSYSID[12] !== 1'bz) && CFGSUBSYSID_delay[12]; // rv 0
  assign CFGSUBSYSID_in[13] = (CFGSUBSYSID[13] !== 1'bz) && CFGSUBSYSID_delay[13]; // rv 0
  assign CFGSUBSYSID_in[14] = (CFGSUBSYSID[14] !== 1'bz) && CFGSUBSYSID_delay[14]; // rv 0
  assign CFGSUBSYSID_in[15] = (CFGSUBSYSID[15] !== 1'bz) && CFGSUBSYSID_delay[15]; // rv 0
  assign CFGSUBSYSID_in[1] = (CFGSUBSYSID[1] !== 1'bz) && CFGSUBSYSID_delay[1]; // rv 0
  assign CFGSUBSYSID_in[2] = (CFGSUBSYSID[2] !== 1'bz) && CFGSUBSYSID_delay[2]; // rv 0
  assign CFGSUBSYSID_in[3] = (CFGSUBSYSID[3] !== 1'bz) && CFGSUBSYSID_delay[3]; // rv 0
  assign CFGSUBSYSID_in[4] = (CFGSUBSYSID[4] !== 1'bz) && CFGSUBSYSID_delay[4]; // rv 0
  assign CFGSUBSYSID_in[5] = (CFGSUBSYSID[5] !== 1'bz) && CFGSUBSYSID_delay[5]; // rv 0
  assign CFGSUBSYSID_in[6] = (CFGSUBSYSID[6] !== 1'bz) && CFGSUBSYSID_delay[6]; // rv 0
  assign CFGSUBSYSID_in[7] = (CFGSUBSYSID[7] !== 1'bz) && CFGSUBSYSID_delay[7]; // rv 0
  assign CFGSUBSYSID_in[8] = (CFGSUBSYSID[8] !== 1'bz) && CFGSUBSYSID_delay[8]; // rv 0
  assign CFGSUBSYSID_in[9] = (CFGSUBSYSID[9] !== 1'bz) && CFGSUBSYSID_delay[9]; // rv 0
  assign CFGSUBSYSVENDID_in[0] = (CFGSUBSYSVENDID[0] !== 1'bz) && CFGSUBSYSVENDID_delay[0]; // rv 0
  assign CFGSUBSYSVENDID_in[10] = (CFGSUBSYSVENDID[10] !== 1'bz) && CFGSUBSYSVENDID_delay[10]; // rv 0
  assign CFGSUBSYSVENDID_in[11] = (CFGSUBSYSVENDID[11] !== 1'bz) && CFGSUBSYSVENDID_delay[11]; // rv 0
  assign CFGSUBSYSVENDID_in[12] = (CFGSUBSYSVENDID[12] !== 1'bz) && CFGSUBSYSVENDID_delay[12]; // rv 0
  assign CFGSUBSYSVENDID_in[13] = (CFGSUBSYSVENDID[13] !== 1'bz) && CFGSUBSYSVENDID_delay[13]; // rv 0
  assign CFGSUBSYSVENDID_in[14] = (CFGSUBSYSVENDID[14] !== 1'bz) && CFGSUBSYSVENDID_delay[14]; // rv 0
  assign CFGSUBSYSVENDID_in[15] = (CFGSUBSYSVENDID[15] !== 1'bz) && CFGSUBSYSVENDID_delay[15]; // rv 0
  assign CFGSUBSYSVENDID_in[1] = (CFGSUBSYSVENDID[1] !== 1'bz) && CFGSUBSYSVENDID_delay[1]; // rv 0
  assign CFGSUBSYSVENDID_in[2] = (CFGSUBSYSVENDID[2] !== 1'bz) && CFGSUBSYSVENDID_delay[2]; // rv 0
  assign CFGSUBSYSVENDID_in[3] = (CFGSUBSYSVENDID[3] !== 1'bz) && CFGSUBSYSVENDID_delay[3]; // rv 0
  assign CFGSUBSYSVENDID_in[4] = (CFGSUBSYSVENDID[4] !== 1'bz) && CFGSUBSYSVENDID_delay[4]; // rv 0
  assign CFGSUBSYSVENDID_in[5] = (CFGSUBSYSVENDID[5] !== 1'bz) && CFGSUBSYSVENDID_delay[5]; // rv 0
  assign CFGSUBSYSVENDID_in[6] = (CFGSUBSYSVENDID[6] !== 1'bz) && CFGSUBSYSVENDID_delay[6]; // rv 0
  assign CFGSUBSYSVENDID_in[7] = (CFGSUBSYSVENDID[7] !== 1'bz) && CFGSUBSYSVENDID_delay[7]; // rv 0
  assign CFGSUBSYSVENDID_in[8] = (CFGSUBSYSVENDID[8] !== 1'bz) && CFGSUBSYSVENDID_delay[8]; // rv 0
  assign CFGSUBSYSVENDID_in[9] = (CFGSUBSYSVENDID[9] !== 1'bz) && CFGSUBSYSVENDID_delay[9]; // rv 0
  assign CFGTPHSTTREADDATAVALID_in = (CFGTPHSTTREADDATAVALID !== 1'bz) && CFGTPHSTTREADDATAVALID_delay; // rv 0
  assign CFGTPHSTTREADDATA_in[0] = (CFGTPHSTTREADDATA[0] !== 1'bz) && CFGTPHSTTREADDATA_delay[0]; // rv 0
  assign CFGTPHSTTREADDATA_in[10] = (CFGTPHSTTREADDATA[10] !== 1'bz) && CFGTPHSTTREADDATA_delay[10]; // rv 0
  assign CFGTPHSTTREADDATA_in[11] = (CFGTPHSTTREADDATA[11] !== 1'bz) && CFGTPHSTTREADDATA_delay[11]; // rv 0
  assign CFGTPHSTTREADDATA_in[12] = (CFGTPHSTTREADDATA[12] !== 1'bz) && CFGTPHSTTREADDATA_delay[12]; // rv 0
  assign CFGTPHSTTREADDATA_in[13] = (CFGTPHSTTREADDATA[13] !== 1'bz) && CFGTPHSTTREADDATA_delay[13]; // rv 0
  assign CFGTPHSTTREADDATA_in[14] = (CFGTPHSTTREADDATA[14] !== 1'bz) && CFGTPHSTTREADDATA_delay[14]; // rv 0
  assign CFGTPHSTTREADDATA_in[15] = (CFGTPHSTTREADDATA[15] !== 1'bz) && CFGTPHSTTREADDATA_delay[15]; // rv 0
  assign CFGTPHSTTREADDATA_in[16] = (CFGTPHSTTREADDATA[16] !== 1'bz) && CFGTPHSTTREADDATA_delay[16]; // rv 0
  assign CFGTPHSTTREADDATA_in[17] = (CFGTPHSTTREADDATA[17] !== 1'bz) && CFGTPHSTTREADDATA_delay[17]; // rv 0
  assign CFGTPHSTTREADDATA_in[18] = (CFGTPHSTTREADDATA[18] !== 1'bz) && CFGTPHSTTREADDATA_delay[18]; // rv 0
  assign CFGTPHSTTREADDATA_in[19] = (CFGTPHSTTREADDATA[19] !== 1'bz) && CFGTPHSTTREADDATA_delay[19]; // rv 0
  assign CFGTPHSTTREADDATA_in[1] = (CFGTPHSTTREADDATA[1] !== 1'bz) && CFGTPHSTTREADDATA_delay[1]; // rv 0
  assign CFGTPHSTTREADDATA_in[20] = (CFGTPHSTTREADDATA[20] !== 1'bz) && CFGTPHSTTREADDATA_delay[20]; // rv 0
  assign CFGTPHSTTREADDATA_in[21] = (CFGTPHSTTREADDATA[21] !== 1'bz) && CFGTPHSTTREADDATA_delay[21]; // rv 0
  assign CFGTPHSTTREADDATA_in[22] = (CFGTPHSTTREADDATA[22] !== 1'bz) && CFGTPHSTTREADDATA_delay[22]; // rv 0
  assign CFGTPHSTTREADDATA_in[23] = (CFGTPHSTTREADDATA[23] !== 1'bz) && CFGTPHSTTREADDATA_delay[23]; // rv 0
  assign CFGTPHSTTREADDATA_in[24] = (CFGTPHSTTREADDATA[24] !== 1'bz) && CFGTPHSTTREADDATA_delay[24]; // rv 0
  assign CFGTPHSTTREADDATA_in[25] = (CFGTPHSTTREADDATA[25] !== 1'bz) && CFGTPHSTTREADDATA_delay[25]; // rv 0
  assign CFGTPHSTTREADDATA_in[26] = (CFGTPHSTTREADDATA[26] !== 1'bz) && CFGTPHSTTREADDATA_delay[26]; // rv 0
  assign CFGTPHSTTREADDATA_in[27] = (CFGTPHSTTREADDATA[27] !== 1'bz) && CFGTPHSTTREADDATA_delay[27]; // rv 0
  assign CFGTPHSTTREADDATA_in[28] = (CFGTPHSTTREADDATA[28] !== 1'bz) && CFGTPHSTTREADDATA_delay[28]; // rv 0
  assign CFGTPHSTTREADDATA_in[29] = (CFGTPHSTTREADDATA[29] !== 1'bz) && CFGTPHSTTREADDATA_delay[29]; // rv 0
  assign CFGTPHSTTREADDATA_in[2] = (CFGTPHSTTREADDATA[2] !== 1'bz) && CFGTPHSTTREADDATA_delay[2]; // rv 0
  assign CFGTPHSTTREADDATA_in[30] = (CFGTPHSTTREADDATA[30] !== 1'bz) && CFGTPHSTTREADDATA_delay[30]; // rv 0
  assign CFGTPHSTTREADDATA_in[31] = (CFGTPHSTTREADDATA[31] !== 1'bz) && CFGTPHSTTREADDATA_delay[31]; // rv 0
  assign CFGTPHSTTREADDATA_in[3] = (CFGTPHSTTREADDATA[3] !== 1'bz) && CFGTPHSTTREADDATA_delay[3]; // rv 0
  assign CFGTPHSTTREADDATA_in[4] = (CFGTPHSTTREADDATA[4] !== 1'bz) && CFGTPHSTTREADDATA_delay[4]; // rv 0
  assign CFGTPHSTTREADDATA_in[5] = (CFGTPHSTTREADDATA[5] !== 1'bz) && CFGTPHSTTREADDATA_delay[5]; // rv 0
  assign CFGTPHSTTREADDATA_in[6] = (CFGTPHSTTREADDATA[6] !== 1'bz) && CFGTPHSTTREADDATA_delay[6]; // rv 0
  assign CFGTPHSTTREADDATA_in[7] = (CFGTPHSTTREADDATA[7] !== 1'bz) && CFGTPHSTTREADDATA_delay[7]; // rv 0
  assign CFGTPHSTTREADDATA_in[8] = (CFGTPHSTTREADDATA[8] !== 1'bz) && CFGTPHSTTREADDATA_delay[8]; // rv 0
  assign CFGTPHSTTREADDATA_in[9] = (CFGTPHSTTREADDATA[9] !== 1'bz) && CFGTPHSTTREADDATA_delay[9]; // rv 0
  assign CFGVENDID_in[0] = (CFGVENDID[0] !== 1'bz) && CFGVENDID_delay[0]; // rv 0
  assign CFGVENDID_in[10] = (CFGVENDID[10] !== 1'bz) && CFGVENDID_delay[10]; // rv 0
  assign CFGVENDID_in[11] = (CFGVENDID[11] !== 1'bz) && CFGVENDID_delay[11]; // rv 0
  assign CFGVENDID_in[12] = (CFGVENDID[12] !== 1'bz) && CFGVENDID_delay[12]; // rv 0
  assign CFGVENDID_in[13] = (CFGVENDID[13] !== 1'bz) && CFGVENDID_delay[13]; // rv 0
  assign CFGVENDID_in[14] = (CFGVENDID[14] !== 1'bz) && CFGVENDID_delay[14]; // rv 0
  assign CFGVENDID_in[15] = (CFGVENDID[15] !== 1'bz) && CFGVENDID_delay[15]; // rv 0
  assign CFGVENDID_in[1] = (CFGVENDID[1] !== 1'bz) && CFGVENDID_delay[1]; // rv 0
  assign CFGVENDID_in[2] = (CFGVENDID[2] !== 1'bz) && CFGVENDID_delay[2]; // rv 0
  assign CFGVENDID_in[3] = (CFGVENDID[3] !== 1'bz) && CFGVENDID_delay[3]; // rv 0
  assign CFGVENDID_in[4] = (CFGVENDID[4] !== 1'bz) && CFGVENDID_delay[4]; // rv 0
  assign CFGVENDID_in[5] = (CFGVENDID[5] !== 1'bz) && CFGVENDID_delay[5]; // rv 0
  assign CFGVENDID_in[6] = (CFGVENDID[6] !== 1'bz) && CFGVENDID_delay[6]; // rv 0
  assign CFGVENDID_in[7] = (CFGVENDID[7] !== 1'bz) && CFGVENDID_delay[7]; // rv 0
  assign CFGVENDID_in[8] = (CFGVENDID[8] !== 1'bz) && CFGVENDID_delay[8]; // rv 0
  assign CFGVENDID_in[9] = (CFGVENDID[9] !== 1'bz) && CFGVENDID_delay[9]; // rv 0
  assign CFGVFFLRDONE_in[0] = (CFGVFFLRDONE[0] !== 1'bz) && CFGVFFLRDONE_delay[0]; // rv 0
  assign CFGVFFLRDONE_in[1] = (CFGVFFLRDONE[1] !== 1'bz) && CFGVFFLRDONE_delay[1]; // rv 0
  assign CFGVFFLRDONE_in[2] = (CFGVFFLRDONE[2] !== 1'bz) && CFGVFFLRDONE_delay[2]; // rv 0
  assign CFGVFFLRDONE_in[3] = (CFGVFFLRDONE[3] !== 1'bz) && CFGVFFLRDONE_delay[3]; // rv 0
  assign CFGVFFLRDONE_in[4] = (CFGVFFLRDONE[4] !== 1'bz) && CFGVFFLRDONE_delay[4]; // rv 0
  assign CFGVFFLRDONE_in[5] = (CFGVFFLRDONE[5] !== 1'bz) && CFGVFFLRDONE_delay[5]; // rv 0
  assign CFGVFFLRDONE_in[6] = (CFGVFFLRDONE[6] !== 1'bz) && CFGVFFLRDONE_delay[6]; // rv 0
  assign CFGVFFLRDONE_in[7] = (CFGVFFLRDONE[7] !== 1'bz) && CFGVFFLRDONE_delay[7]; // rv 0
  assign CONFMCAPREQUESTBYCONF_in = (CONFMCAPREQUESTBYCONF !== 1'bz) && CONFMCAPREQUESTBYCONF_delay; // rv 0
  assign CONFREQDATA_in[0] = (CONFREQDATA[0] !== 1'bz) && CONFREQDATA_delay[0]; // rv 0
  assign CONFREQDATA_in[10] = (CONFREQDATA[10] !== 1'bz) && CONFREQDATA_delay[10]; // rv 0
  assign CONFREQDATA_in[11] = (CONFREQDATA[11] !== 1'bz) && CONFREQDATA_delay[11]; // rv 0
  assign CONFREQDATA_in[12] = (CONFREQDATA[12] !== 1'bz) && CONFREQDATA_delay[12]; // rv 0
  assign CONFREQDATA_in[13] = (CONFREQDATA[13] !== 1'bz) && CONFREQDATA_delay[13]; // rv 0
  assign CONFREQDATA_in[14] = (CONFREQDATA[14] !== 1'bz) && CONFREQDATA_delay[14]; // rv 0
  assign CONFREQDATA_in[15] = (CONFREQDATA[15] !== 1'bz) && CONFREQDATA_delay[15]; // rv 0
  assign CONFREQDATA_in[16] = (CONFREQDATA[16] !== 1'bz) && CONFREQDATA_delay[16]; // rv 0
  assign CONFREQDATA_in[17] = (CONFREQDATA[17] !== 1'bz) && CONFREQDATA_delay[17]; // rv 0
  assign CONFREQDATA_in[18] = (CONFREQDATA[18] !== 1'bz) && CONFREQDATA_delay[18]; // rv 0
  assign CONFREQDATA_in[19] = (CONFREQDATA[19] !== 1'bz) && CONFREQDATA_delay[19]; // rv 0
  assign CONFREQDATA_in[1] = (CONFREQDATA[1] !== 1'bz) && CONFREQDATA_delay[1]; // rv 0
  assign CONFREQDATA_in[20] = (CONFREQDATA[20] !== 1'bz) && CONFREQDATA_delay[20]; // rv 0
  assign CONFREQDATA_in[21] = (CONFREQDATA[21] !== 1'bz) && CONFREQDATA_delay[21]; // rv 0
  assign CONFREQDATA_in[22] = (CONFREQDATA[22] !== 1'bz) && CONFREQDATA_delay[22]; // rv 0
  assign CONFREQDATA_in[23] = (CONFREQDATA[23] !== 1'bz) && CONFREQDATA_delay[23]; // rv 0
  assign CONFREQDATA_in[24] = (CONFREQDATA[24] !== 1'bz) && CONFREQDATA_delay[24]; // rv 0
  assign CONFREQDATA_in[25] = (CONFREQDATA[25] !== 1'bz) && CONFREQDATA_delay[25]; // rv 0
  assign CONFREQDATA_in[26] = (CONFREQDATA[26] !== 1'bz) && CONFREQDATA_delay[26]; // rv 0
  assign CONFREQDATA_in[27] = (CONFREQDATA[27] !== 1'bz) && CONFREQDATA_delay[27]; // rv 0
  assign CONFREQDATA_in[28] = (CONFREQDATA[28] !== 1'bz) && CONFREQDATA_delay[28]; // rv 0
  assign CONFREQDATA_in[29] = (CONFREQDATA[29] !== 1'bz) && CONFREQDATA_delay[29]; // rv 0
  assign CONFREQDATA_in[2] = (CONFREQDATA[2] !== 1'bz) && CONFREQDATA_delay[2]; // rv 0
  assign CONFREQDATA_in[30] = (CONFREQDATA[30] !== 1'bz) && CONFREQDATA_delay[30]; // rv 0
  assign CONFREQDATA_in[31] = (CONFREQDATA[31] !== 1'bz) && CONFREQDATA_delay[31]; // rv 0
  assign CONFREQDATA_in[3] = (CONFREQDATA[3] !== 1'bz) && CONFREQDATA_delay[3]; // rv 0
  assign CONFREQDATA_in[4] = (CONFREQDATA[4] !== 1'bz) && CONFREQDATA_delay[4]; // rv 0
  assign CONFREQDATA_in[5] = (CONFREQDATA[5] !== 1'bz) && CONFREQDATA_delay[5]; // rv 0
  assign CONFREQDATA_in[6] = (CONFREQDATA[6] !== 1'bz) && CONFREQDATA_delay[6]; // rv 0
  assign CONFREQDATA_in[7] = (CONFREQDATA[7] !== 1'bz) && CONFREQDATA_delay[7]; // rv 0
  assign CONFREQDATA_in[8] = (CONFREQDATA[8] !== 1'bz) && CONFREQDATA_delay[8]; // rv 0
  assign CONFREQDATA_in[9] = (CONFREQDATA[9] !== 1'bz) && CONFREQDATA_delay[9]; // rv 0
  assign CONFREQREGNUM_in[0] = (CONFREQREGNUM[0] !== 1'bz) && CONFREQREGNUM_delay[0]; // rv 0
  assign CONFREQREGNUM_in[1] = (CONFREQREGNUM[1] !== 1'bz) && CONFREQREGNUM_delay[1]; // rv 0
  assign CONFREQREGNUM_in[2] = (CONFREQREGNUM[2] !== 1'bz) && CONFREQREGNUM_delay[2]; // rv 0
  assign CONFREQREGNUM_in[3] = (CONFREQREGNUM[3] !== 1'bz) && CONFREQREGNUM_delay[3]; // rv 0
  assign CONFREQTYPE_in[0] = (CONFREQTYPE[0] !== 1'bz) && CONFREQTYPE_delay[0]; // rv 0
  assign CONFREQTYPE_in[1] = (CONFREQTYPE[1] !== 1'bz) && CONFREQTYPE_delay[1]; // rv 0
  assign CONFREQVALID_in = (CONFREQVALID !== 1'bz) && CONFREQVALID_delay; // rv 0
  assign CORECLKMICOMPLETIONRAML_in = (CORECLKMICOMPLETIONRAML !== 1'bz) && CORECLKMICOMPLETIONRAML_delay; // rv 0
  assign CORECLKMICOMPLETIONRAMU_in = (CORECLKMICOMPLETIONRAMU !== 1'bz) && CORECLKMICOMPLETIONRAMU_delay; // rv 0
  assign CORECLKMIREPLAYRAM_in = (CORECLKMIREPLAYRAM !== 1'bz) && CORECLKMIREPLAYRAM_delay; // rv 0
  assign CORECLKMIREQUESTRAM_in = (CORECLKMIREQUESTRAM !== 1'bz) && CORECLKMIREQUESTRAM_delay; // rv 0
  assign CORECLK_in = (CORECLK !== 1'bz) && CORECLK_delay; // rv 0
  assign DBGCFGLOCALMGMTREGOVERRIDE_in = (DBGCFGLOCALMGMTREGOVERRIDE !== 1'bz) && DBGCFGLOCALMGMTREGOVERRIDE_delay; // rv 0
  assign DBGDATASEL_in[0] = (DBGDATASEL[0] !== 1'bz) && DBGDATASEL_delay[0]; // rv 0
  assign DBGDATASEL_in[1] = (DBGDATASEL[1] !== 1'bz) && DBGDATASEL_delay[1]; // rv 0
  assign DBGDATASEL_in[2] = (DBGDATASEL[2] !== 1'bz) && DBGDATASEL_delay[2]; // rv 0
  assign DBGDATASEL_in[3] = (DBGDATASEL[3] !== 1'bz) && DBGDATASEL_delay[3]; // rv 0
  assign DRPADDR_in[0] = (DRPADDR[0] !== 1'bz) && DRPADDR_delay[0]; // rv 0
  assign DRPADDR_in[1] = (DRPADDR[1] !== 1'bz) && DRPADDR_delay[1]; // rv 0
  assign DRPADDR_in[2] = (DRPADDR[2] !== 1'bz) && DRPADDR_delay[2]; // rv 0
  assign DRPADDR_in[3] = (DRPADDR[3] !== 1'bz) && DRPADDR_delay[3]; // rv 0
  assign DRPADDR_in[4] = (DRPADDR[4] !== 1'bz) && DRPADDR_delay[4]; // rv 0
  assign DRPADDR_in[5] = (DRPADDR[5] !== 1'bz) && DRPADDR_delay[5]; // rv 0
  assign DRPADDR_in[6] = (DRPADDR[6] !== 1'bz) && DRPADDR_delay[6]; // rv 0
  assign DRPADDR_in[7] = (DRPADDR[7] !== 1'bz) && DRPADDR_delay[7]; // rv 0
  assign DRPADDR_in[8] = (DRPADDR[8] !== 1'bz) && DRPADDR_delay[8]; // rv 0
  assign DRPADDR_in[9] = (DRPADDR[9] !== 1'bz) && DRPADDR_delay[9]; // rv 0
  assign DRPCLK_in = (DRPCLK !== 1'bz) && DRPCLK_delay; // rv 0
  assign DRPDI_in[0] = (DRPDI[0] !== 1'bz) && DRPDI_delay[0]; // rv 0
  assign DRPDI_in[10] = (DRPDI[10] !== 1'bz) && DRPDI_delay[10]; // rv 0
  assign DRPDI_in[11] = (DRPDI[11] !== 1'bz) && DRPDI_delay[11]; // rv 0
  assign DRPDI_in[12] = (DRPDI[12] !== 1'bz) && DRPDI_delay[12]; // rv 0
  assign DRPDI_in[13] = (DRPDI[13] !== 1'bz) && DRPDI_delay[13]; // rv 0
  assign DRPDI_in[14] = (DRPDI[14] !== 1'bz) && DRPDI_delay[14]; // rv 0
  assign DRPDI_in[15] = (DRPDI[15] !== 1'bz) && DRPDI_delay[15]; // rv 0
  assign DRPDI_in[1] = (DRPDI[1] !== 1'bz) && DRPDI_delay[1]; // rv 0
  assign DRPDI_in[2] = (DRPDI[2] !== 1'bz) && DRPDI_delay[2]; // rv 0
  assign DRPDI_in[3] = (DRPDI[3] !== 1'bz) && DRPDI_delay[3]; // rv 0
  assign DRPDI_in[4] = (DRPDI[4] !== 1'bz) && DRPDI_delay[4]; // rv 0
  assign DRPDI_in[5] = (DRPDI[5] !== 1'bz) && DRPDI_delay[5]; // rv 0
  assign DRPDI_in[6] = (DRPDI[6] !== 1'bz) && DRPDI_delay[6]; // rv 0
  assign DRPDI_in[7] = (DRPDI[7] !== 1'bz) && DRPDI_delay[7]; // rv 0
  assign DRPDI_in[8] = (DRPDI[8] !== 1'bz) && DRPDI_delay[8]; // rv 0
  assign DRPDI_in[9] = (DRPDI[9] !== 1'bz) && DRPDI_delay[9]; // rv 0
  assign DRPEN_in = (DRPEN !== 1'bz) && DRPEN_delay; // rv 0
  assign DRPWE_in = (DRPWE !== 1'bz) && DRPWE_delay; // rv 0
  assign LL2LMSAXISTXTUSER_in[0] = (LL2LMSAXISTXTUSER[0] !== 1'bz) && LL2LMSAXISTXTUSER_delay[0]; // rv 0
  assign LL2LMSAXISTXTUSER_in[10] = (LL2LMSAXISTXTUSER[10] !== 1'bz) && LL2LMSAXISTXTUSER_delay[10]; // rv 0
  assign LL2LMSAXISTXTUSER_in[11] = (LL2LMSAXISTXTUSER[11] !== 1'bz) && LL2LMSAXISTXTUSER_delay[11]; // rv 0
  assign LL2LMSAXISTXTUSER_in[12] = (LL2LMSAXISTXTUSER[12] !== 1'bz) && LL2LMSAXISTXTUSER_delay[12]; // rv 0
  assign LL2LMSAXISTXTUSER_in[13] = (LL2LMSAXISTXTUSER[13] !== 1'bz) && LL2LMSAXISTXTUSER_delay[13]; // rv 0
  assign LL2LMSAXISTXTUSER_in[1] = (LL2LMSAXISTXTUSER[1] !== 1'bz) && LL2LMSAXISTXTUSER_delay[1]; // rv 0
  assign LL2LMSAXISTXTUSER_in[2] = (LL2LMSAXISTXTUSER[2] !== 1'bz) && LL2LMSAXISTXTUSER_delay[2]; // rv 0
  assign LL2LMSAXISTXTUSER_in[3] = (LL2LMSAXISTXTUSER[3] !== 1'bz) && LL2LMSAXISTXTUSER_delay[3]; // rv 0
  assign LL2LMSAXISTXTUSER_in[4] = (LL2LMSAXISTXTUSER[4] !== 1'bz) && LL2LMSAXISTXTUSER_delay[4]; // rv 0
  assign LL2LMSAXISTXTUSER_in[5] = (LL2LMSAXISTXTUSER[5] !== 1'bz) && LL2LMSAXISTXTUSER_delay[5]; // rv 0
  assign LL2LMSAXISTXTUSER_in[6] = (LL2LMSAXISTXTUSER[6] !== 1'bz) && LL2LMSAXISTXTUSER_delay[6]; // rv 0
  assign LL2LMSAXISTXTUSER_in[7] = (LL2LMSAXISTXTUSER[7] !== 1'bz) && LL2LMSAXISTXTUSER_delay[7]; // rv 0
  assign LL2LMSAXISTXTUSER_in[8] = (LL2LMSAXISTXTUSER[8] !== 1'bz) && LL2LMSAXISTXTUSER_delay[8]; // rv 0
  assign LL2LMSAXISTXTUSER_in[9] = (LL2LMSAXISTXTUSER[9] !== 1'bz) && LL2LMSAXISTXTUSER_delay[9]; // rv 0
  assign LL2LMSAXISTXTVALID_in = (LL2LMSAXISTXTVALID !== 1'bz) && LL2LMSAXISTXTVALID_delay; // rv 0
  assign LL2LMTXTLPID0_in[0] = (LL2LMTXTLPID0[0] !== 1'bz) && LL2LMTXTLPID0_delay[0]; // rv 0
  assign LL2LMTXTLPID0_in[1] = (LL2LMTXTLPID0[1] !== 1'bz) && LL2LMTXTLPID0_delay[1]; // rv 0
  assign LL2LMTXTLPID0_in[2] = (LL2LMTXTLPID0[2] !== 1'bz) && LL2LMTXTLPID0_delay[2]; // rv 0
  assign LL2LMTXTLPID0_in[3] = (LL2LMTXTLPID0[3] !== 1'bz) && LL2LMTXTLPID0_delay[3]; // rv 0
  assign LL2LMTXTLPID1_in[0] = (LL2LMTXTLPID1[0] !== 1'bz) && LL2LMTXTLPID1_delay[0]; // rv 0
  assign LL2LMTXTLPID1_in[1] = (LL2LMTXTLPID1[1] !== 1'bz) && LL2LMTXTLPID1_delay[1]; // rv 0
  assign LL2LMTXTLPID1_in[2] = (LL2LMTXTLPID1[2] !== 1'bz) && LL2LMTXTLPID1_delay[2]; // rv 0
  assign LL2LMTXTLPID1_in[3] = (LL2LMTXTLPID1[3] !== 1'bz) && LL2LMTXTLPID1_delay[3]; // rv 0
  assign MAXISCQTREADY_in[0] = (MAXISCQTREADY[0] !== 1'bz) && MAXISCQTREADY_delay[0]; // rv 0
  assign MAXISCQTREADY_in[10] = (MAXISCQTREADY[10] !== 1'bz) && MAXISCQTREADY_delay[10]; // rv 0
  assign MAXISCQTREADY_in[11] = (MAXISCQTREADY[11] !== 1'bz) && MAXISCQTREADY_delay[11]; // rv 0
  assign MAXISCQTREADY_in[12] = (MAXISCQTREADY[12] !== 1'bz) && MAXISCQTREADY_delay[12]; // rv 0
  assign MAXISCQTREADY_in[13] = (MAXISCQTREADY[13] !== 1'bz) && MAXISCQTREADY_delay[13]; // rv 0
  assign MAXISCQTREADY_in[14] = (MAXISCQTREADY[14] !== 1'bz) && MAXISCQTREADY_delay[14]; // rv 0
  assign MAXISCQTREADY_in[15] = (MAXISCQTREADY[15] !== 1'bz) && MAXISCQTREADY_delay[15]; // rv 0
  assign MAXISCQTREADY_in[16] = (MAXISCQTREADY[16] !== 1'bz) && MAXISCQTREADY_delay[16]; // rv 0
  assign MAXISCQTREADY_in[17] = (MAXISCQTREADY[17] !== 1'bz) && MAXISCQTREADY_delay[17]; // rv 0
  assign MAXISCQTREADY_in[18] = (MAXISCQTREADY[18] !== 1'bz) && MAXISCQTREADY_delay[18]; // rv 0
  assign MAXISCQTREADY_in[19] = (MAXISCQTREADY[19] !== 1'bz) && MAXISCQTREADY_delay[19]; // rv 0
  assign MAXISCQTREADY_in[1] = (MAXISCQTREADY[1] !== 1'bz) && MAXISCQTREADY_delay[1]; // rv 0
  assign MAXISCQTREADY_in[20] = (MAXISCQTREADY[20] !== 1'bz) && MAXISCQTREADY_delay[20]; // rv 0
  assign MAXISCQTREADY_in[21] = (MAXISCQTREADY[21] !== 1'bz) && MAXISCQTREADY_delay[21]; // rv 0
  assign MAXISCQTREADY_in[2] = (MAXISCQTREADY[2] !== 1'bz) && MAXISCQTREADY_delay[2]; // rv 0
  assign MAXISCQTREADY_in[3] = (MAXISCQTREADY[3] !== 1'bz) && MAXISCQTREADY_delay[3]; // rv 0
  assign MAXISCQTREADY_in[4] = (MAXISCQTREADY[4] !== 1'bz) && MAXISCQTREADY_delay[4]; // rv 0
  assign MAXISCQTREADY_in[5] = (MAXISCQTREADY[5] !== 1'bz) && MAXISCQTREADY_delay[5]; // rv 0
  assign MAXISCQTREADY_in[6] = (MAXISCQTREADY[6] !== 1'bz) && MAXISCQTREADY_delay[6]; // rv 0
  assign MAXISCQTREADY_in[7] = (MAXISCQTREADY[7] !== 1'bz) && MAXISCQTREADY_delay[7]; // rv 0
  assign MAXISCQTREADY_in[8] = (MAXISCQTREADY[8] !== 1'bz) && MAXISCQTREADY_delay[8]; // rv 0
  assign MAXISCQTREADY_in[9] = (MAXISCQTREADY[9] !== 1'bz) && MAXISCQTREADY_delay[9]; // rv 0
  assign MAXISRCTREADY_in[0] = (MAXISRCTREADY[0] !== 1'bz) && MAXISRCTREADY_delay[0]; // rv 0
  assign MAXISRCTREADY_in[10] = (MAXISRCTREADY[10] !== 1'bz) && MAXISRCTREADY_delay[10]; // rv 0
  assign MAXISRCTREADY_in[11] = (MAXISRCTREADY[11] !== 1'bz) && MAXISRCTREADY_delay[11]; // rv 0
  assign MAXISRCTREADY_in[12] = (MAXISRCTREADY[12] !== 1'bz) && MAXISRCTREADY_delay[12]; // rv 0
  assign MAXISRCTREADY_in[13] = (MAXISRCTREADY[13] !== 1'bz) && MAXISRCTREADY_delay[13]; // rv 0
  assign MAXISRCTREADY_in[14] = (MAXISRCTREADY[14] !== 1'bz) && MAXISRCTREADY_delay[14]; // rv 0
  assign MAXISRCTREADY_in[15] = (MAXISRCTREADY[15] !== 1'bz) && MAXISRCTREADY_delay[15]; // rv 0
  assign MAXISRCTREADY_in[16] = (MAXISRCTREADY[16] !== 1'bz) && MAXISRCTREADY_delay[16]; // rv 0
  assign MAXISRCTREADY_in[17] = (MAXISRCTREADY[17] !== 1'bz) && MAXISRCTREADY_delay[17]; // rv 0
  assign MAXISRCTREADY_in[18] = (MAXISRCTREADY[18] !== 1'bz) && MAXISRCTREADY_delay[18]; // rv 0
  assign MAXISRCTREADY_in[19] = (MAXISRCTREADY[19] !== 1'bz) && MAXISRCTREADY_delay[19]; // rv 0
  assign MAXISRCTREADY_in[1] = (MAXISRCTREADY[1] !== 1'bz) && MAXISRCTREADY_delay[1]; // rv 0
  assign MAXISRCTREADY_in[20] = (MAXISRCTREADY[20] !== 1'bz) && MAXISRCTREADY_delay[20]; // rv 0
  assign MAXISRCTREADY_in[21] = (MAXISRCTREADY[21] !== 1'bz) && MAXISRCTREADY_delay[21]; // rv 0
  assign MAXISRCTREADY_in[2] = (MAXISRCTREADY[2] !== 1'bz) && MAXISRCTREADY_delay[2]; // rv 0
  assign MAXISRCTREADY_in[3] = (MAXISRCTREADY[3] !== 1'bz) && MAXISRCTREADY_delay[3]; // rv 0
  assign MAXISRCTREADY_in[4] = (MAXISRCTREADY[4] !== 1'bz) && MAXISRCTREADY_delay[4]; // rv 0
  assign MAXISRCTREADY_in[5] = (MAXISRCTREADY[5] !== 1'bz) && MAXISRCTREADY_delay[5]; // rv 0
  assign MAXISRCTREADY_in[6] = (MAXISRCTREADY[6] !== 1'bz) && MAXISRCTREADY_delay[6]; // rv 0
  assign MAXISRCTREADY_in[7] = (MAXISRCTREADY[7] !== 1'bz) && MAXISRCTREADY_delay[7]; // rv 0
  assign MAXISRCTREADY_in[8] = (MAXISRCTREADY[8] !== 1'bz) && MAXISRCTREADY_delay[8]; // rv 0
  assign MAXISRCTREADY_in[9] = (MAXISRCTREADY[9] !== 1'bz) && MAXISRCTREADY_delay[9]; // rv 0
  assign MCAPCLK_in = (MCAPCLK !== 1'bz) && MCAPCLK_delay; // rv 0
  assign MCAPPERST0B_in = (MCAPPERST0B === 1'bz) || MCAPPERST0B_delay; // rv 1
  assign MCAPPERST1B_in = (MCAPPERST1B === 1'bz) || MCAPPERST1B_delay; // rv 1
  assign MGMTRESETN_in = (MGMTRESETN !== 1'bz) && MGMTRESETN_delay; // rv 0
  assign MGMTSTICKYRESETN_in = (MGMTSTICKYRESETN !== 1'bz) && MGMTSTICKYRESETN_delay; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[0] = (MICOMPLETIONRAMREADDATA[0] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[0]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[100] = (MICOMPLETIONRAMREADDATA[100] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[100]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[101] = (MICOMPLETIONRAMREADDATA[101] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[101]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[102] = (MICOMPLETIONRAMREADDATA[102] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[102]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[103] = (MICOMPLETIONRAMREADDATA[103] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[103]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[104] = (MICOMPLETIONRAMREADDATA[104] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[104]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[105] = (MICOMPLETIONRAMREADDATA[105] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[105]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[106] = (MICOMPLETIONRAMREADDATA[106] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[106]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[107] = (MICOMPLETIONRAMREADDATA[107] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[107]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[108] = (MICOMPLETIONRAMREADDATA[108] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[108]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[109] = (MICOMPLETIONRAMREADDATA[109] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[109]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[10] = (MICOMPLETIONRAMREADDATA[10] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[10]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[110] = (MICOMPLETIONRAMREADDATA[110] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[110]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[111] = (MICOMPLETIONRAMREADDATA[111] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[111]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[112] = (MICOMPLETIONRAMREADDATA[112] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[112]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[113] = (MICOMPLETIONRAMREADDATA[113] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[113]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[114] = (MICOMPLETIONRAMREADDATA[114] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[114]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[115] = (MICOMPLETIONRAMREADDATA[115] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[115]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[116] = (MICOMPLETIONRAMREADDATA[116] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[116]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[117] = (MICOMPLETIONRAMREADDATA[117] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[117]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[118] = (MICOMPLETIONRAMREADDATA[118] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[118]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[119] = (MICOMPLETIONRAMREADDATA[119] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[119]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[11] = (MICOMPLETIONRAMREADDATA[11] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[11]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[120] = (MICOMPLETIONRAMREADDATA[120] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[120]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[121] = (MICOMPLETIONRAMREADDATA[121] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[121]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[122] = (MICOMPLETIONRAMREADDATA[122] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[122]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[123] = (MICOMPLETIONRAMREADDATA[123] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[123]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[124] = (MICOMPLETIONRAMREADDATA[124] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[124]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[125] = (MICOMPLETIONRAMREADDATA[125] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[125]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[126] = (MICOMPLETIONRAMREADDATA[126] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[126]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[127] = (MICOMPLETIONRAMREADDATA[127] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[127]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[128] = (MICOMPLETIONRAMREADDATA[128] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[128]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[129] = (MICOMPLETIONRAMREADDATA[129] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[129]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[12] = (MICOMPLETIONRAMREADDATA[12] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[12]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[130] = (MICOMPLETIONRAMREADDATA[130] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[130]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[131] = (MICOMPLETIONRAMREADDATA[131] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[131]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[132] = (MICOMPLETIONRAMREADDATA[132] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[132]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[133] = (MICOMPLETIONRAMREADDATA[133] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[133]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[134] = (MICOMPLETIONRAMREADDATA[134] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[134]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[135] = (MICOMPLETIONRAMREADDATA[135] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[135]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[136] = (MICOMPLETIONRAMREADDATA[136] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[136]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[137] = (MICOMPLETIONRAMREADDATA[137] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[137]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[138] = (MICOMPLETIONRAMREADDATA[138] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[138]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[139] = (MICOMPLETIONRAMREADDATA[139] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[139]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[13] = (MICOMPLETIONRAMREADDATA[13] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[13]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[140] = (MICOMPLETIONRAMREADDATA[140] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[140]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[141] = (MICOMPLETIONRAMREADDATA[141] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[141]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[142] = (MICOMPLETIONRAMREADDATA[142] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[142]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[143] = (MICOMPLETIONRAMREADDATA[143] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[143]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[14] = (MICOMPLETIONRAMREADDATA[14] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[14]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[15] = (MICOMPLETIONRAMREADDATA[15] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[15]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[16] = (MICOMPLETIONRAMREADDATA[16] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[16]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[17] = (MICOMPLETIONRAMREADDATA[17] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[17]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[18] = (MICOMPLETIONRAMREADDATA[18] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[18]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[19] = (MICOMPLETIONRAMREADDATA[19] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[19]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[1] = (MICOMPLETIONRAMREADDATA[1] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[1]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[20] = (MICOMPLETIONRAMREADDATA[20] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[20]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[21] = (MICOMPLETIONRAMREADDATA[21] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[21]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[22] = (MICOMPLETIONRAMREADDATA[22] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[22]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[23] = (MICOMPLETIONRAMREADDATA[23] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[23]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[24] = (MICOMPLETIONRAMREADDATA[24] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[24]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[25] = (MICOMPLETIONRAMREADDATA[25] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[25]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[26] = (MICOMPLETIONRAMREADDATA[26] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[26]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[27] = (MICOMPLETIONRAMREADDATA[27] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[27]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[28] = (MICOMPLETIONRAMREADDATA[28] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[28]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[29] = (MICOMPLETIONRAMREADDATA[29] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[29]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[2] = (MICOMPLETIONRAMREADDATA[2] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[2]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[30] = (MICOMPLETIONRAMREADDATA[30] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[30]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[31] = (MICOMPLETIONRAMREADDATA[31] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[31]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[32] = (MICOMPLETIONRAMREADDATA[32] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[32]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[33] = (MICOMPLETIONRAMREADDATA[33] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[33]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[34] = (MICOMPLETIONRAMREADDATA[34] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[34]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[35] = (MICOMPLETIONRAMREADDATA[35] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[35]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[36] = (MICOMPLETIONRAMREADDATA[36] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[36]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[37] = (MICOMPLETIONRAMREADDATA[37] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[37]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[38] = (MICOMPLETIONRAMREADDATA[38] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[38]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[39] = (MICOMPLETIONRAMREADDATA[39] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[39]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[3] = (MICOMPLETIONRAMREADDATA[3] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[3]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[40] = (MICOMPLETIONRAMREADDATA[40] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[40]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[41] = (MICOMPLETIONRAMREADDATA[41] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[41]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[42] = (MICOMPLETIONRAMREADDATA[42] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[42]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[43] = (MICOMPLETIONRAMREADDATA[43] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[43]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[44] = (MICOMPLETIONRAMREADDATA[44] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[44]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[45] = (MICOMPLETIONRAMREADDATA[45] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[45]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[46] = (MICOMPLETIONRAMREADDATA[46] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[46]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[47] = (MICOMPLETIONRAMREADDATA[47] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[47]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[48] = (MICOMPLETIONRAMREADDATA[48] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[48]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[49] = (MICOMPLETIONRAMREADDATA[49] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[49]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[4] = (MICOMPLETIONRAMREADDATA[4] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[4]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[50] = (MICOMPLETIONRAMREADDATA[50] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[50]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[51] = (MICOMPLETIONRAMREADDATA[51] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[51]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[52] = (MICOMPLETIONRAMREADDATA[52] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[52]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[53] = (MICOMPLETIONRAMREADDATA[53] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[53]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[54] = (MICOMPLETIONRAMREADDATA[54] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[54]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[55] = (MICOMPLETIONRAMREADDATA[55] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[55]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[56] = (MICOMPLETIONRAMREADDATA[56] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[56]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[57] = (MICOMPLETIONRAMREADDATA[57] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[57]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[58] = (MICOMPLETIONRAMREADDATA[58] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[58]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[59] = (MICOMPLETIONRAMREADDATA[59] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[59]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[5] = (MICOMPLETIONRAMREADDATA[5] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[5]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[60] = (MICOMPLETIONRAMREADDATA[60] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[60]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[61] = (MICOMPLETIONRAMREADDATA[61] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[61]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[62] = (MICOMPLETIONRAMREADDATA[62] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[62]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[63] = (MICOMPLETIONRAMREADDATA[63] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[63]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[64] = (MICOMPLETIONRAMREADDATA[64] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[64]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[65] = (MICOMPLETIONRAMREADDATA[65] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[65]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[66] = (MICOMPLETIONRAMREADDATA[66] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[66]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[67] = (MICOMPLETIONRAMREADDATA[67] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[67]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[68] = (MICOMPLETIONRAMREADDATA[68] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[68]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[69] = (MICOMPLETIONRAMREADDATA[69] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[69]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[6] = (MICOMPLETIONRAMREADDATA[6] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[6]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[70] = (MICOMPLETIONRAMREADDATA[70] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[70]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[71] = (MICOMPLETIONRAMREADDATA[71] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[71]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[72] = (MICOMPLETIONRAMREADDATA[72] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[72]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[73] = (MICOMPLETIONRAMREADDATA[73] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[73]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[74] = (MICOMPLETIONRAMREADDATA[74] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[74]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[75] = (MICOMPLETIONRAMREADDATA[75] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[75]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[76] = (MICOMPLETIONRAMREADDATA[76] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[76]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[77] = (MICOMPLETIONRAMREADDATA[77] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[77]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[78] = (MICOMPLETIONRAMREADDATA[78] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[78]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[79] = (MICOMPLETIONRAMREADDATA[79] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[79]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[7] = (MICOMPLETIONRAMREADDATA[7] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[7]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[80] = (MICOMPLETIONRAMREADDATA[80] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[80]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[81] = (MICOMPLETIONRAMREADDATA[81] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[81]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[82] = (MICOMPLETIONRAMREADDATA[82] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[82]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[83] = (MICOMPLETIONRAMREADDATA[83] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[83]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[84] = (MICOMPLETIONRAMREADDATA[84] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[84]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[85] = (MICOMPLETIONRAMREADDATA[85] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[85]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[86] = (MICOMPLETIONRAMREADDATA[86] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[86]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[87] = (MICOMPLETIONRAMREADDATA[87] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[87]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[88] = (MICOMPLETIONRAMREADDATA[88] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[88]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[89] = (MICOMPLETIONRAMREADDATA[89] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[89]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[8] = (MICOMPLETIONRAMREADDATA[8] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[8]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[90] = (MICOMPLETIONRAMREADDATA[90] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[90]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[91] = (MICOMPLETIONRAMREADDATA[91] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[91]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[92] = (MICOMPLETIONRAMREADDATA[92] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[92]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[93] = (MICOMPLETIONRAMREADDATA[93] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[93]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[94] = (MICOMPLETIONRAMREADDATA[94] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[94]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[95] = (MICOMPLETIONRAMREADDATA[95] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[95]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[96] = (MICOMPLETIONRAMREADDATA[96] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[96]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[97] = (MICOMPLETIONRAMREADDATA[97] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[97]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[98] = (MICOMPLETIONRAMREADDATA[98] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[98]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[99] = (MICOMPLETIONRAMREADDATA[99] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[99]; // rv 0
  assign MICOMPLETIONRAMREADDATA_in[9] = (MICOMPLETIONRAMREADDATA[9] !== 1'bz) && MICOMPLETIONRAMREADDATA_delay[9]; // rv 0
  assign MIREPLAYRAMREADDATA_in[0] = (MIREPLAYRAMREADDATA[0] !== 1'bz) && MIREPLAYRAMREADDATA_delay[0]; // rv 0
  assign MIREPLAYRAMREADDATA_in[100] = (MIREPLAYRAMREADDATA[100] !== 1'bz) && MIREPLAYRAMREADDATA_delay[100]; // rv 0
  assign MIREPLAYRAMREADDATA_in[101] = (MIREPLAYRAMREADDATA[101] !== 1'bz) && MIREPLAYRAMREADDATA_delay[101]; // rv 0
  assign MIREPLAYRAMREADDATA_in[102] = (MIREPLAYRAMREADDATA[102] !== 1'bz) && MIREPLAYRAMREADDATA_delay[102]; // rv 0
  assign MIREPLAYRAMREADDATA_in[103] = (MIREPLAYRAMREADDATA[103] !== 1'bz) && MIREPLAYRAMREADDATA_delay[103]; // rv 0
  assign MIREPLAYRAMREADDATA_in[104] = (MIREPLAYRAMREADDATA[104] !== 1'bz) && MIREPLAYRAMREADDATA_delay[104]; // rv 0
  assign MIREPLAYRAMREADDATA_in[105] = (MIREPLAYRAMREADDATA[105] !== 1'bz) && MIREPLAYRAMREADDATA_delay[105]; // rv 0
  assign MIREPLAYRAMREADDATA_in[106] = (MIREPLAYRAMREADDATA[106] !== 1'bz) && MIREPLAYRAMREADDATA_delay[106]; // rv 0
  assign MIREPLAYRAMREADDATA_in[107] = (MIREPLAYRAMREADDATA[107] !== 1'bz) && MIREPLAYRAMREADDATA_delay[107]; // rv 0
  assign MIREPLAYRAMREADDATA_in[108] = (MIREPLAYRAMREADDATA[108] !== 1'bz) && MIREPLAYRAMREADDATA_delay[108]; // rv 0
  assign MIREPLAYRAMREADDATA_in[109] = (MIREPLAYRAMREADDATA[109] !== 1'bz) && MIREPLAYRAMREADDATA_delay[109]; // rv 0
  assign MIREPLAYRAMREADDATA_in[10] = (MIREPLAYRAMREADDATA[10] !== 1'bz) && MIREPLAYRAMREADDATA_delay[10]; // rv 0
  assign MIREPLAYRAMREADDATA_in[110] = (MIREPLAYRAMREADDATA[110] !== 1'bz) && MIREPLAYRAMREADDATA_delay[110]; // rv 0
  assign MIREPLAYRAMREADDATA_in[111] = (MIREPLAYRAMREADDATA[111] !== 1'bz) && MIREPLAYRAMREADDATA_delay[111]; // rv 0
  assign MIREPLAYRAMREADDATA_in[112] = (MIREPLAYRAMREADDATA[112] !== 1'bz) && MIREPLAYRAMREADDATA_delay[112]; // rv 0
  assign MIREPLAYRAMREADDATA_in[113] = (MIREPLAYRAMREADDATA[113] !== 1'bz) && MIREPLAYRAMREADDATA_delay[113]; // rv 0
  assign MIREPLAYRAMREADDATA_in[114] = (MIREPLAYRAMREADDATA[114] !== 1'bz) && MIREPLAYRAMREADDATA_delay[114]; // rv 0
  assign MIREPLAYRAMREADDATA_in[115] = (MIREPLAYRAMREADDATA[115] !== 1'bz) && MIREPLAYRAMREADDATA_delay[115]; // rv 0
  assign MIREPLAYRAMREADDATA_in[116] = (MIREPLAYRAMREADDATA[116] !== 1'bz) && MIREPLAYRAMREADDATA_delay[116]; // rv 0
  assign MIREPLAYRAMREADDATA_in[117] = (MIREPLAYRAMREADDATA[117] !== 1'bz) && MIREPLAYRAMREADDATA_delay[117]; // rv 0
  assign MIREPLAYRAMREADDATA_in[118] = (MIREPLAYRAMREADDATA[118] !== 1'bz) && MIREPLAYRAMREADDATA_delay[118]; // rv 0
  assign MIREPLAYRAMREADDATA_in[119] = (MIREPLAYRAMREADDATA[119] !== 1'bz) && MIREPLAYRAMREADDATA_delay[119]; // rv 0
  assign MIREPLAYRAMREADDATA_in[11] = (MIREPLAYRAMREADDATA[11] !== 1'bz) && MIREPLAYRAMREADDATA_delay[11]; // rv 0
  assign MIREPLAYRAMREADDATA_in[120] = (MIREPLAYRAMREADDATA[120] !== 1'bz) && MIREPLAYRAMREADDATA_delay[120]; // rv 0
  assign MIREPLAYRAMREADDATA_in[121] = (MIREPLAYRAMREADDATA[121] !== 1'bz) && MIREPLAYRAMREADDATA_delay[121]; // rv 0
  assign MIREPLAYRAMREADDATA_in[122] = (MIREPLAYRAMREADDATA[122] !== 1'bz) && MIREPLAYRAMREADDATA_delay[122]; // rv 0
  assign MIREPLAYRAMREADDATA_in[123] = (MIREPLAYRAMREADDATA[123] !== 1'bz) && MIREPLAYRAMREADDATA_delay[123]; // rv 0
  assign MIREPLAYRAMREADDATA_in[124] = (MIREPLAYRAMREADDATA[124] !== 1'bz) && MIREPLAYRAMREADDATA_delay[124]; // rv 0
  assign MIREPLAYRAMREADDATA_in[125] = (MIREPLAYRAMREADDATA[125] !== 1'bz) && MIREPLAYRAMREADDATA_delay[125]; // rv 0
  assign MIREPLAYRAMREADDATA_in[126] = (MIREPLAYRAMREADDATA[126] !== 1'bz) && MIREPLAYRAMREADDATA_delay[126]; // rv 0
  assign MIREPLAYRAMREADDATA_in[127] = (MIREPLAYRAMREADDATA[127] !== 1'bz) && MIREPLAYRAMREADDATA_delay[127]; // rv 0
  assign MIREPLAYRAMREADDATA_in[128] = (MIREPLAYRAMREADDATA[128] !== 1'bz) && MIREPLAYRAMREADDATA_delay[128]; // rv 0
  assign MIREPLAYRAMREADDATA_in[129] = (MIREPLAYRAMREADDATA[129] !== 1'bz) && MIREPLAYRAMREADDATA_delay[129]; // rv 0
  assign MIREPLAYRAMREADDATA_in[12] = (MIREPLAYRAMREADDATA[12] !== 1'bz) && MIREPLAYRAMREADDATA_delay[12]; // rv 0
  assign MIREPLAYRAMREADDATA_in[130] = (MIREPLAYRAMREADDATA[130] !== 1'bz) && MIREPLAYRAMREADDATA_delay[130]; // rv 0
  assign MIREPLAYRAMREADDATA_in[131] = (MIREPLAYRAMREADDATA[131] !== 1'bz) && MIREPLAYRAMREADDATA_delay[131]; // rv 0
  assign MIREPLAYRAMREADDATA_in[132] = (MIREPLAYRAMREADDATA[132] !== 1'bz) && MIREPLAYRAMREADDATA_delay[132]; // rv 0
  assign MIREPLAYRAMREADDATA_in[133] = (MIREPLAYRAMREADDATA[133] !== 1'bz) && MIREPLAYRAMREADDATA_delay[133]; // rv 0
  assign MIREPLAYRAMREADDATA_in[134] = (MIREPLAYRAMREADDATA[134] !== 1'bz) && MIREPLAYRAMREADDATA_delay[134]; // rv 0
  assign MIREPLAYRAMREADDATA_in[135] = (MIREPLAYRAMREADDATA[135] !== 1'bz) && MIREPLAYRAMREADDATA_delay[135]; // rv 0
  assign MIREPLAYRAMREADDATA_in[136] = (MIREPLAYRAMREADDATA[136] !== 1'bz) && MIREPLAYRAMREADDATA_delay[136]; // rv 0
  assign MIREPLAYRAMREADDATA_in[137] = (MIREPLAYRAMREADDATA[137] !== 1'bz) && MIREPLAYRAMREADDATA_delay[137]; // rv 0
  assign MIREPLAYRAMREADDATA_in[138] = (MIREPLAYRAMREADDATA[138] !== 1'bz) && MIREPLAYRAMREADDATA_delay[138]; // rv 0
  assign MIREPLAYRAMREADDATA_in[139] = (MIREPLAYRAMREADDATA[139] !== 1'bz) && MIREPLAYRAMREADDATA_delay[139]; // rv 0
  assign MIREPLAYRAMREADDATA_in[13] = (MIREPLAYRAMREADDATA[13] !== 1'bz) && MIREPLAYRAMREADDATA_delay[13]; // rv 0
  assign MIREPLAYRAMREADDATA_in[140] = (MIREPLAYRAMREADDATA[140] !== 1'bz) && MIREPLAYRAMREADDATA_delay[140]; // rv 0
  assign MIREPLAYRAMREADDATA_in[141] = (MIREPLAYRAMREADDATA[141] !== 1'bz) && MIREPLAYRAMREADDATA_delay[141]; // rv 0
  assign MIREPLAYRAMREADDATA_in[142] = (MIREPLAYRAMREADDATA[142] !== 1'bz) && MIREPLAYRAMREADDATA_delay[142]; // rv 0
  assign MIREPLAYRAMREADDATA_in[143] = (MIREPLAYRAMREADDATA[143] !== 1'bz) && MIREPLAYRAMREADDATA_delay[143]; // rv 0
  assign MIREPLAYRAMREADDATA_in[14] = (MIREPLAYRAMREADDATA[14] !== 1'bz) && MIREPLAYRAMREADDATA_delay[14]; // rv 0
  assign MIREPLAYRAMREADDATA_in[15] = (MIREPLAYRAMREADDATA[15] !== 1'bz) && MIREPLAYRAMREADDATA_delay[15]; // rv 0
  assign MIREPLAYRAMREADDATA_in[16] = (MIREPLAYRAMREADDATA[16] !== 1'bz) && MIREPLAYRAMREADDATA_delay[16]; // rv 0
  assign MIREPLAYRAMREADDATA_in[17] = (MIREPLAYRAMREADDATA[17] !== 1'bz) && MIREPLAYRAMREADDATA_delay[17]; // rv 0
  assign MIREPLAYRAMREADDATA_in[18] = (MIREPLAYRAMREADDATA[18] !== 1'bz) && MIREPLAYRAMREADDATA_delay[18]; // rv 0
  assign MIREPLAYRAMREADDATA_in[19] = (MIREPLAYRAMREADDATA[19] !== 1'bz) && MIREPLAYRAMREADDATA_delay[19]; // rv 0
  assign MIREPLAYRAMREADDATA_in[1] = (MIREPLAYRAMREADDATA[1] !== 1'bz) && MIREPLAYRAMREADDATA_delay[1]; // rv 0
  assign MIREPLAYRAMREADDATA_in[20] = (MIREPLAYRAMREADDATA[20] !== 1'bz) && MIREPLAYRAMREADDATA_delay[20]; // rv 0
  assign MIREPLAYRAMREADDATA_in[21] = (MIREPLAYRAMREADDATA[21] !== 1'bz) && MIREPLAYRAMREADDATA_delay[21]; // rv 0
  assign MIREPLAYRAMREADDATA_in[22] = (MIREPLAYRAMREADDATA[22] !== 1'bz) && MIREPLAYRAMREADDATA_delay[22]; // rv 0
  assign MIREPLAYRAMREADDATA_in[23] = (MIREPLAYRAMREADDATA[23] !== 1'bz) && MIREPLAYRAMREADDATA_delay[23]; // rv 0
  assign MIREPLAYRAMREADDATA_in[24] = (MIREPLAYRAMREADDATA[24] !== 1'bz) && MIREPLAYRAMREADDATA_delay[24]; // rv 0
  assign MIREPLAYRAMREADDATA_in[25] = (MIREPLAYRAMREADDATA[25] !== 1'bz) && MIREPLAYRAMREADDATA_delay[25]; // rv 0
  assign MIREPLAYRAMREADDATA_in[26] = (MIREPLAYRAMREADDATA[26] !== 1'bz) && MIREPLAYRAMREADDATA_delay[26]; // rv 0
  assign MIREPLAYRAMREADDATA_in[27] = (MIREPLAYRAMREADDATA[27] !== 1'bz) && MIREPLAYRAMREADDATA_delay[27]; // rv 0
  assign MIREPLAYRAMREADDATA_in[28] = (MIREPLAYRAMREADDATA[28] !== 1'bz) && MIREPLAYRAMREADDATA_delay[28]; // rv 0
  assign MIREPLAYRAMREADDATA_in[29] = (MIREPLAYRAMREADDATA[29] !== 1'bz) && MIREPLAYRAMREADDATA_delay[29]; // rv 0
  assign MIREPLAYRAMREADDATA_in[2] = (MIREPLAYRAMREADDATA[2] !== 1'bz) && MIREPLAYRAMREADDATA_delay[2]; // rv 0
  assign MIREPLAYRAMREADDATA_in[30] = (MIREPLAYRAMREADDATA[30] !== 1'bz) && MIREPLAYRAMREADDATA_delay[30]; // rv 0
  assign MIREPLAYRAMREADDATA_in[31] = (MIREPLAYRAMREADDATA[31] !== 1'bz) && MIREPLAYRAMREADDATA_delay[31]; // rv 0
  assign MIREPLAYRAMREADDATA_in[32] = (MIREPLAYRAMREADDATA[32] !== 1'bz) && MIREPLAYRAMREADDATA_delay[32]; // rv 0
  assign MIREPLAYRAMREADDATA_in[33] = (MIREPLAYRAMREADDATA[33] !== 1'bz) && MIREPLAYRAMREADDATA_delay[33]; // rv 0
  assign MIREPLAYRAMREADDATA_in[34] = (MIREPLAYRAMREADDATA[34] !== 1'bz) && MIREPLAYRAMREADDATA_delay[34]; // rv 0
  assign MIREPLAYRAMREADDATA_in[35] = (MIREPLAYRAMREADDATA[35] !== 1'bz) && MIREPLAYRAMREADDATA_delay[35]; // rv 0
  assign MIREPLAYRAMREADDATA_in[36] = (MIREPLAYRAMREADDATA[36] !== 1'bz) && MIREPLAYRAMREADDATA_delay[36]; // rv 0
  assign MIREPLAYRAMREADDATA_in[37] = (MIREPLAYRAMREADDATA[37] !== 1'bz) && MIREPLAYRAMREADDATA_delay[37]; // rv 0
  assign MIREPLAYRAMREADDATA_in[38] = (MIREPLAYRAMREADDATA[38] !== 1'bz) && MIREPLAYRAMREADDATA_delay[38]; // rv 0
  assign MIREPLAYRAMREADDATA_in[39] = (MIREPLAYRAMREADDATA[39] !== 1'bz) && MIREPLAYRAMREADDATA_delay[39]; // rv 0
  assign MIREPLAYRAMREADDATA_in[3] = (MIREPLAYRAMREADDATA[3] !== 1'bz) && MIREPLAYRAMREADDATA_delay[3]; // rv 0
  assign MIREPLAYRAMREADDATA_in[40] = (MIREPLAYRAMREADDATA[40] !== 1'bz) && MIREPLAYRAMREADDATA_delay[40]; // rv 0
  assign MIREPLAYRAMREADDATA_in[41] = (MIREPLAYRAMREADDATA[41] !== 1'bz) && MIREPLAYRAMREADDATA_delay[41]; // rv 0
  assign MIREPLAYRAMREADDATA_in[42] = (MIREPLAYRAMREADDATA[42] !== 1'bz) && MIREPLAYRAMREADDATA_delay[42]; // rv 0
  assign MIREPLAYRAMREADDATA_in[43] = (MIREPLAYRAMREADDATA[43] !== 1'bz) && MIREPLAYRAMREADDATA_delay[43]; // rv 0
  assign MIREPLAYRAMREADDATA_in[44] = (MIREPLAYRAMREADDATA[44] !== 1'bz) && MIREPLAYRAMREADDATA_delay[44]; // rv 0
  assign MIREPLAYRAMREADDATA_in[45] = (MIREPLAYRAMREADDATA[45] !== 1'bz) && MIREPLAYRAMREADDATA_delay[45]; // rv 0
  assign MIREPLAYRAMREADDATA_in[46] = (MIREPLAYRAMREADDATA[46] !== 1'bz) && MIREPLAYRAMREADDATA_delay[46]; // rv 0
  assign MIREPLAYRAMREADDATA_in[47] = (MIREPLAYRAMREADDATA[47] !== 1'bz) && MIREPLAYRAMREADDATA_delay[47]; // rv 0
  assign MIREPLAYRAMREADDATA_in[48] = (MIREPLAYRAMREADDATA[48] !== 1'bz) && MIREPLAYRAMREADDATA_delay[48]; // rv 0
  assign MIREPLAYRAMREADDATA_in[49] = (MIREPLAYRAMREADDATA[49] !== 1'bz) && MIREPLAYRAMREADDATA_delay[49]; // rv 0
  assign MIREPLAYRAMREADDATA_in[4] = (MIREPLAYRAMREADDATA[4] !== 1'bz) && MIREPLAYRAMREADDATA_delay[4]; // rv 0
  assign MIREPLAYRAMREADDATA_in[50] = (MIREPLAYRAMREADDATA[50] !== 1'bz) && MIREPLAYRAMREADDATA_delay[50]; // rv 0
  assign MIREPLAYRAMREADDATA_in[51] = (MIREPLAYRAMREADDATA[51] !== 1'bz) && MIREPLAYRAMREADDATA_delay[51]; // rv 0
  assign MIREPLAYRAMREADDATA_in[52] = (MIREPLAYRAMREADDATA[52] !== 1'bz) && MIREPLAYRAMREADDATA_delay[52]; // rv 0
  assign MIREPLAYRAMREADDATA_in[53] = (MIREPLAYRAMREADDATA[53] !== 1'bz) && MIREPLAYRAMREADDATA_delay[53]; // rv 0
  assign MIREPLAYRAMREADDATA_in[54] = (MIREPLAYRAMREADDATA[54] !== 1'bz) && MIREPLAYRAMREADDATA_delay[54]; // rv 0
  assign MIREPLAYRAMREADDATA_in[55] = (MIREPLAYRAMREADDATA[55] !== 1'bz) && MIREPLAYRAMREADDATA_delay[55]; // rv 0
  assign MIREPLAYRAMREADDATA_in[56] = (MIREPLAYRAMREADDATA[56] !== 1'bz) && MIREPLAYRAMREADDATA_delay[56]; // rv 0
  assign MIREPLAYRAMREADDATA_in[57] = (MIREPLAYRAMREADDATA[57] !== 1'bz) && MIREPLAYRAMREADDATA_delay[57]; // rv 0
  assign MIREPLAYRAMREADDATA_in[58] = (MIREPLAYRAMREADDATA[58] !== 1'bz) && MIREPLAYRAMREADDATA_delay[58]; // rv 0
  assign MIREPLAYRAMREADDATA_in[59] = (MIREPLAYRAMREADDATA[59] !== 1'bz) && MIREPLAYRAMREADDATA_delay[59]; // rv 0
  assign MIREPLAYRAMREADDATA_in[5] = (MIREPLAYRAMREADDATA[5] !== 1'bz) && MIREPLAYRAMREADDATA_delay[5]; // rv 0
  assign MIREPLAYRAMREADDATA_in[60] = (MIREPLAYRAMREADDATA[60] !== 1'bz) && MIREPLAYRAMREADDATA_delay[60]; // rv 0
  assign MIREPLAYRAMREADDATA_in[61] = (MIREPLAYRAMREADDATA[61] !== 1'bz) && MIREPLAYRAMREADDATA_delay[61]; // rv 0
  assign MIREPLAYRAMREADDATA_in[62] = (MIREPLAYRAMREADDATA[62] !== 1'bz) && MIREPLAYRAMREADDATA_delay[62]; // rv 0
  assign MIREPLAYRAMREADDATA_in[63] = (MIREPLAYRAMREADDATA[63] !== 1'bz) && MIREPLAYRAMREADDATA_delay[63]; // rv 0
  assign MIREPLAYRAMREADDATA_in[64] = (MIREPLAYRAMREADDATA[64] !== 1'bz) && MIREPLAYRAMREADDATA_delay[64]; // rv 0
  assign MIREPLAYRAMREADDATA_in[65] = (MIREPLAYRAMREADDATA[65] !== 1'bz) && MIREPLAYRAMREADDATA_delay[65]; // rv 0
  assign MIREPLAYRAMREADDATA_in[66] = (MIREPLAYRAMREADDATA[66] !== 1'bz) && MIREPLAYRAMREADDATA_delay[66]; // rv 0
  assign MIREPLAYRAMREADDATA_in[67] = (MIREPLAYRAMREADDATA[67] !== 1'bz) && MIREPLAYRAMREADDATA_delay[67]; // rv 0
  assign MIREPLAYRAMREADDATA_in[68] = (MIREPLAYRAMREADDATA[68] !== 1'bz) && MIREPLAYRAMREADDATA_delay[68]; // rv 0
  assign MIREPLAYRAMREADDATA_in[69] = (MIREPLAYRAMREADDATA[69] !== 1'bz) && MIREPLAYRAMREADDATA_delay[69]; // rv 0
  assign MIREPLAYRAMREADDATA_in[6] = (MIREPLAYRAMREADDATA[6] !== 1'bz) && MIREPLAYRAMREADDATA_delay[6]; // rv 0
  assign MIREPLAYRAMREADDATA_in[70] = (MIREPLAYRAMREADDATA[70] !== 1'bz) && MIREPLAYRAMREADDATA_delay[70]; // rv 0
  assign MIREPLAYRAMREADDATA_in[71] = (MIREPLAYRAMREADDATA[71] !== 1'bz) && MIREPLAYRAMREADDATA_delay[71]; // rv 0
  assign MIREPLAYRAMREADDATA_in[72] = (MIREPLAYRAMREADDATA[72] !== 1'bz) && MIREPLAYRAMREADDATA_delay[72]; // rv 0
  assign MIREPLAYRAMREADDATA_in[73] = (MIREPLAYRAMREADDATA[73] !== 1'bz) && MIREPLAYRAMREADDATA_delay[73]; // rv 0
  assign MIREPLAYRAMREADDATA_in[74] = (MIREPLAYRAMREADDATA[74] !== 1'bz) && MIREPLAYRAMREADDATA_delay[74]; // rv 0
  assign MIREPLAYRAMREADDATA_in[75] = (MIREPLAYRAMREADDATA[75] !== 1'bz) && MIREPLAYRAMREADDATA_delay[75]; // rv 0
  assign MIREPLAYRAMREADDATA_in[76] = (MIREPLAYRAMREADDATA[76] !== 1'bz) && MIREPLAYRAMREADDATA_delay[76]; // rv 0
  assign MIREPLAYRAMREADDATA_in[77] = (MIREPLAYRAMREADDATA[77] !== 1'bz) && MIREPLAYRAMREADDATA_delay[77]; // rv 0
  assign MIREPLAYRAMREADDATA_in[78] = (MIREPLAYRAMREADDATA[78] !== 1'bz) && MIREPLAYRAMREADDATA_delay[78]; // rv 0
  assign MIREPLAYRAMREADDATA_in[79] = (MIREPLAYRAMREADDATA[79] !== 1'bz) && MIREPLAYRAMREADDATA_delay[79]; // rv 0
  assign MIREPLAYRAMREADDATA_in[7] = (MIREPLAYRAMREADDATA[7] !== 1'bz) && MIREPLAYRAMREADDATA_delay[7]; // rv 0
  assign MIREPLAYRAMREADDATA_in[80] = (MIREPLAYRAMREADDATA[80] !== 1'bz) && MIREPLAYRAMREADDATA_delay[80]; // rv 0
  assign MIREPLAYRAMREADDATA_in[81] = (MIREPLAYRAMREADDATA[81] !== 1'bz) && MIREPLAYRAMREADDATA_delay[81]; // rv 0
  assign MIREPLAYRAMREADDATA_in[82] = (MIREPLAYRAMREADDATA[82] !== 1'bz) && MIREPLAYRAMREADDATA_delay[82]; // rv 0
  assign MIREPLAYRAMREADDATA_in[83] = (MIREPLAYRAMREADDATA[83] !== 1'bz) && MIREPLAYRAMREADDATA_delay[83]; // rv 0
  assign MIREPLAYRAMREADDATA_in[84] = (MIREPLAYRAMREADDATA[84] !== 1'bz) && MIREPLAYRAMREADDATA_delay[84]; // rv 0
  assign MIREPLAYRAMREADDATA_in[85] = (MIREPLAYRAMREADDATA[85] !== 1'bz) && MIREPLAYRAMREADDATA_delay[85]; // rv 0
  assign MIREPLAYRAMREADDATA_in[86] = (MIREPLAYRAMREADDATA[86] !== 1'bz) && MIREPLAYRAMREADDATA_delay[86]; // rv 0
  assign MIREPLAYRAMREADDATA_in[87] = (MIREPLAYRAMREADDATA[87] !== 1'bz) && MIREPLAYRAMREADDATA_delay[87]; // rv 0
  assign MIREPLAYRAMREADDATA_in[88] = (MIREPLAYRAMREADDATA[88] !== 1'bz) && MIREPLAYRAMREADDATA_delay[88]; // rv 0
  assign MIREPLAYRAMREADDATA_in[89] = (MIREPLAYRAMREADDATA[89] !== 1'bz) && MIREPLAYRAMREADDATA_delay[89]; // rv 0
  assign MIREPLAYRAMREADDATA_in[8] = (MIREPLAYRAMREADDATA[8] !== 1'bz) && MIREPLAYRAMREADDATA_delay[8]; // rv 0
  assign MIREPLAYRAMREADDATA_in[90] = (MIREPLAYRAMREADDATA[90] !== 1'bz) && MIREPLAYRAMREADDATA_delay[90]; // rv 0
  assign MIREPLAYRAMREADDATA_in[91] = (MIREPLAYRAMREADDATA[91] !== 1'bz) && MIREPLAYRAMREADDATA_delay[91]; // rv 0
  assign MIREPLAYRAMREADDATA_in[92] = (MIREPLAYRAMREADDATA[92] !== 1'bz) && MIREPLAYRAMREADDATA_delay[92]; // rv 0
  assign MIREPLAYRAMREADDATA_in[93] = (MIREPLAYRAMREADDATA[93] !== 1'bz) && MIREPLAYRAMREADDATA_delay[93]; // rv 0
  assign MIREPLAYRAMREADDATA_in[94] = (MIREPLAYRAMREADDATA[94] !== 1'bz) && MIREPLAYRAMREADDATA_delay[94]; // rv 0
  assign MIREPLAYRAMREADDATA_in[95] = (MIREPLAYRAMREADDATA[95] !== 1'bz) && MIREPLAYRAMREADDATA_delay[95]; // rv 0
  assign MIREPLAYRAMREADDATA_in[96] = (MIREPLAYRAMREADDATA[96] !== 1'bz) && MIREPLAYRAMREADDATA_delay[96]; // rv 0
  assign MIREPLAYRAMREADDATA_in[97] = (MIREPLAYRAMREADDATA[97] !== 1'bz) && MIREPLAYRAMREADDATA_delay[97]; // rv 0
  assign MIREPLAYRAMREADDATA_in[98] = (MIREPLAYRAMREADDATA[98] !== 1'bz) && MIREPLAYRAMREADDATA_delay[98]; // rv 0
  assign MIREPLAYRAMREADDATA_in[99] = (MIREPLAYRAMREADDATA[99] !== 1'bz) && MIREPLAYRAMREADDATA_delay[99]; // rv 0
  assign MIREPLAYRAMREADDATA_in[9] = (MIREPLAYRAMREADDATA[9] !== 1'bz) && MIREPLAYRAMREADDATA_delay[9]; // rv 0
  assign MIREQUESTRAMREADDATA_in[0] = (MIREQUESTRAMREADDATA[0] !== 1'bz) && MIREQUESTRAMREADDATA_delay[0]; // rv 0
  assign MIREQUESTRAMREADDATA_in[100] = (MIREQUESTRAMREADDATA[100] !== 1'bz) && MIREQUESTRAMREADDATA_delay[100]; // rv 0
  assign MIREQUESTRAMREADDATA_in[101] = (MIREQUESTRAMREADDATA[101] !== 1'bz) && MIREQUESTRAMREADDATA_delay[101]; // rv 0
  assign MIREQUESTRAMREADDATA_in[102] = (MIREQUESTRAMREADDATA[102] !== 1'bz) && MIREQUESTRAMREADDATA_delay[102]; // rv 0
  assign MIREQUESTRAMREADDATA_in[103] = (MIREQUESTRAMREADDATA[103] !== 1'bz) && MIREQUESTRAMREADDATA_delay[103]; // rv 0
  assign MIREQUESTRAMREADDATA_in[104] = (MIREQUESTRAMREADDATA[104] !== 1'bz) && MIREQUESTRAMREADDATA_delay[104]; // rv 0
  assign MIREQUESTRAMREADDATA_in[105] = (MIREQUESTRAMREADDATA[105] !== 1'bz) && MIREQUESTRAMREADDATA_delay[105]; // rv 0
  assign MIREQUESTRAMREADDATA_in[106] = (MIREQUESTRAMREADDATA[106] !== 1'bz) && MIREQUESTRAMREADDATA_delay[106]; // rv 0
  assign MIREQUESTRAMREADDATA_in[107] = (MIREQUESTRAMREADDATA[107] !== 1'bz) && MIREQUESTRAMREADDATA_delay[107]; // rv 0
  assign MIREQUESTRAMREADDATA_in[108] = (MIREQUESTRAMREADDATA[108] !== 1'bz) && MIREQUESTRAMREADDATA_delay[108]; // rv 0
  assign MIREQUESTRAMREADDATA_in[109] = (MIREQUESTRAMREADDATA[109] !== 1'bz) && MIREQUESTRAMREADDATA_delay[109]; // rv 0
  assign MIREQUESTRAMREADDATA_in[10] = (MIREQUESTRAMREADDATA[10] !== 1'bz) && MIREQUESTRAMREADDATA_delay[10]; // rv 0
  assign MIREQUESTRAMREADDATA_in[110] = (MIREQUESTRAMREADDATA[110] !== 1'bz) && MIREQUESTRAMREADDATA_delay[110]; // rv 0
  assign MIREQUESTRAMREADDATA_in[111] = (MIREQUESTRAMREADDATA[111] !== 1'bz) && MIREQUESTRAMREADDATA_delay[111]; // rv 0
  assign MIREQUESTRAMREADDATA_in[112] = (MIREQUESTRAMREADDATA[112] !== 1'bz) && MIREQUESTRAMREADDATA_delay[112]; // rv 0
  assign MIREQUESTRAMREADDATA_in[113] = (MIREQUESTRAMREADDATA[113] !== 1'bz) && MIREQUESTRAMREADDATA_delay[113]; // rv 0
  assign MIREQUESTRAMREADDATA_in[114] = (MIREQUESTRAMREADDATA[114] !== 1'bz) && MIREQUESTRAMREADDATA_delay[114]; // rv 0
  assign MIREQUESTRAMREADDATA_in[115] = (MIREQUESTRAMREADDATA[115] !== 1'bz) && MIREQUESTRAMREADDATA_delay[115]; // rv 0
  assign MIREQUESTRAMREADDATA_in[116] = (MIREQUESTRAMREADDATA[116] !== 1'bz) && MIREQUESTRAMREADDATA_delay[116]; // rv 0
  assign MIREQUESTRAMREADDATA_in[117] = (MIREQUESTRAMREADDATA[117] !== 1'bz) && MIREQUESTRAMREADDATA_delay[117]; // rv 0
  assign MIREQUESTRAMREADDATA_in[118] = (MIREQUESTRAMREADDATA[118] !== 1'bz) && MIREQUESTRAMREADDATA_delay[118]; // rv 0
  assign MIREQUESTRAMREADDATA_in[119] = (MIREQUESTRAMREADDATA[119] !== 1'bz) && MIREQUESTRAMREADDATA_delay[119]; // rv 0
  assign MIREQUESTRAMREADDATA_in[11] = (MIREQUESTRAMREADDATA[11] !== 1'bz) && MIREQUESTRAMREADDATA_delay[11]; // rv 0
  assign MIREQUESTRAMREADDATA_in[120] = (MIREQUESTRAMREADDATA[120] !== 1'bz) && MIREQUESTRAMREADDATA_delay[120]; // rv 0
  assign MIREQUESTRAMREADDATA_in[121] = (MIREQUESTRAMREADDATA[121] !== 1'bz) && MIREQUESTRAMREADDATA_delay[121]; // rv 0
  assign MIREQUESTRAMREADDATA_in[122] = (MIREQUESTRAMREADDATA[122] !== 1'bz) && MIREQUESTRAMREADDATA_delay[122]; // rv 0
  assign MIREQUESTRAMREADDATA_in[123] = (MIREQUESTRAMREADDATA[123] !== 1'bz) && MIREQUESTRAMREADDATA_delay[123]; // rv 0
  assign MIREQUESTRAMREADDATA_in[124] = (MIREQUESTRAMREADDATA[124] !== 1'bz) && MIREQUESTRAMREADDATA_delay[124]; // rv 0
  assign MIREQUESTRAMREADDATA_in[125] = (MIREQUESTRAMREADDATA[125] !== 1'bz) && MIREQUESTRAMREADDATA_delay[125]; // rv 0
  assign MIREQUESTRAMREADDATA_in[126] = (MIREQUESTRAMREADDATA[126] !== 1'bz) && MIREQUESTRAMREADDATA_delay[126]; // rv 0
  assign MIREQUESTRAMREADDATA_in[127] = (MIREQUESTRAMREADDATA[127] !== 1'bz) && MIREQUESTRAMREADDATA_delay[127]; // rv 0
  assign MIREQUESTRAMREADDATA_in[128] = (MIREQUESTRAMREADDATA[128] !== 1'bz) && MIREQUESTRAMREADDATA_delay[128]; // rv 0
  assign MIREQUESTRAMREADDATA_in[129] = (MIREQUESTRAMREADDATA[129] !== 1'bz) && MIREQUESTRAMREADDATA_delay[129]; // rv 0
  assign MIREQUESTRAMREADDATA_in[12] = (MIREQUESTRAMREADDATA[12] !== 1'bz) && MIREQUESTRAMREADDATA_delay[12]; // rv 0
  assign MIREQUESTRAMREADDATA_in[130] = (MIREQUESTRAMREADDATA[130] !== 1'bz) && MIREQUESTRAMREADDATA_delay[130]; // rv 0
  assign MIREQUESTRAMREADDATA_in[131] = (MIREQUESTRAMREADDATA[131] !== 1'bz) && MIREQUESTRAMREADDATA_delay[131]; // rv 0
  assign MIREQUESTRAMREADDATA_in[132] = (MIREQUESTRAMREADDATA[132] !== 1'bz) && MIREQUESTRAMREADDATA_delay[132]; // rv 0
  assign MIREQUESTRAMREADDATA_in[133] = (MIREQUESTRAMREADDATA[133] !== 1'bz) && MIREQUESTRAMREADDATA_delay[133]; // rv 0
  assign MIREQUESTRAMREADDATA_in[134] = (MIREQUESTRAMREADDATA[134] !== 1'bz) && MIREQUESTRAMREADDATA_delay[134]; // rv 0
  assign MIREQUESTRAMREADDATA_in[135] = (MIREQUESTRAMREADDATA[135] !== 1'bz) && MIREQUESTRAMREADDATA_delay[135]; // rv 0
  assign MIREQUESTRAMREADDATA_in[136] = (MIREQUESTRAMREADDATA[136] !== 1'bz) && MIREQUESTRAMREADDATA_delay[136]; // rv 0
  assign MIREQUESTRAMREADDATA_in[137] = (MIREQUESTRAMREADDATA[137] !== 1'bz) && MIREQUESTRAMREADDATA_delay[137]; // rv 0
  assign MIREQUESTRAMREADDATA_in[138] = (MIREQUESTRAMREADDATA[138] !== 1'bz) && MIREQUESTRAMREADDATA_delay[138]; // rv 0
  assign MIREQUESTRAMREADDATA_in[139] = (MIREQUESTRAMREADDATA[139] !== 1'bz) && MIREQUESTRAMREADDATA_delay[139]; // rv 0
  assign MIREQUESTRAMREADDATA_in[13] = (MIREQUESTRAMREADDATA[13] !== 1'bz) && MIREQUESTRAMREADDATA_delay[13]; // rv 0
  assign MIREQUESTRAMREADDATA_in[140] = (MIREQUESTRAMREADDATA[140] !== 1'bz) && MIREQUESTRAMREADDATA_delay[140]; // rv 0
  assign MIREQUESTRAMREADDATA_in[141] = (MIREQUESTRAMREADDATA[141] !== 1'bz) && MIREQUESTRAMREADDATA_delay[141]; // rv 0
  assign MIREQUESTRAMREADDATA_in[142] = (MIREQUESTRAMREADDATA[142] !== 1'bz) && MIREQUESTRAMREADDATA_delay[142]; // rv 0
  assign MIREQUESTRAMREADDATA_in[143] = (MIREQUESTRAMREADDATA[143] !== 1'bz) && MIREQUESTRAMREADDATA_delay[143]; // rv 0
  assign MIREQUESTRAMREADDATA_in[14] = (MIREQUESTRAMREADDATA[14] !== 1'bz) && MIREQUESTRAMREADDATA_delay[14]; // rv 0
  assign MIREQUESTRAMREADDATA_in[15] = (MIREQUESTRAMREADDATA[15] !== 1'bz) && MIREQUESTRAMREADDATA_delay[15]; // rv 0
  assign MIREQUESTRAMREADDATA_in[16] = (MIREQUESTRAMREADDATA[16] !== 1'bz) && MIREQUESTRAMREADDATA_delay[16]; // rv 0
  assign MIREQUESTRAMREADDATA_in[17] = (MIREQUESTRAMREADDATA[17] !== 1'bz) && MIREQUESTRAMREADDATA_delay[17]; // rv 0
  assign MIREQUESTRAMREADDATA_in[18] = (MIREQUESTRAMREADDATA[18] !== 1'bz) && MIREQUESTRAMREADDATA_delay[18]; // rv 0
  assign MIREQUESTRAMREADDATA_in[19] = (MIREQUESTRAMREADDATA[19] !== 1'bz) && MIREQUESTRAMREADDATA_delay[19]; // rv 0
  assign MIREQUESTRAMREADDATA_in[1] = (MIREQUESTRAMREADDATA[1] !== 1'bz) && MIREQUESTRAMREADDATA_delay[1]; // rv 0
  assign MIREQUESTRAMREADDATA_in[20] = (MIREQUESTRAMREADDATA[20] !== 1'bz) && MIREQUESTRAMREADDATA_delay[20]; // rv 0
  assign MIREQUESTRAMREADDATA_in[21] = (MIREQUESTRAMREADDATA[21] !== 1'bz) && MIREQUESTRAMREADDATA_delay[21]; // rv 0
  assign MIREQUESTRAMREADDATA_in[22] = (MIREQUESTRAMREADDATA[22] !== 1'bz) && MIREQUESTRAMREADDATA_delay[22]; // rv 0
  assign MIREQUESTRAMREADDATA_in[23] = (MIREQUESTRAMREADDATA[23] !== 1'bz) && MIREQUESTRAMREADDATA_delay[23]; // rv 0
  assign MIREQUESTRAMREADDATA_in[24] = (MIREQUESTRAMREADDATA[24] !== 1'bz) && MIREQUESTRAMREADDATA_delay[24]; // rv 0
  assign MIREQUESTRAMREADDATA_in[25] = (MIREQUESTRAMREADDATA[25] !== 1'bz) && MIREQUESTRAMREADDATA_delay[25]; // rv 0
  assign MIREQUESTRAMREADDATA_in[26] = (MIREQUESTRAMREADDATA[26] !== 1'bz) && MIREQUESTRAMREADDATA_delay[26]; // rv 0
  assign MIREQUESTRAMREADDATA_in[27] = (MIREQUESTRAMREADDATA[27] !== 1'bz) && MIREQUESTRAMREADDATA_delay[27]; // rv 0
  assign MIREQUESTRAMREADDATA_in[28] = (MIREQUESTRAMREADDATA[28] !== 1'bz) && MIREQUESTRAMREADDATA_delay[28]; // rv 0
  assign MIREQUESTRAMREADDATA_in[29] = (MIREQUESTRAMREADDATA[29] !== 1'bz) && MIREQUESTRAMREADDATA_delay[29]; // rv 0
  assign MIREQUESTRAMREADDATA_in[2] = (MIREQUESTRAMREADDATA[2] !== 1'bz) && MIREQUESTRAMREADDATA_delay[2]; // rv 0
  assign MIREQUESTRAMREADDATA_in[30] = (MIREQUESTRAMREADDATA[30] !== 1'bz) && MIREQUESTRAMREADDATA_delay[30]; // rv 0
  assign MIREQUESTRAMREADDATA_in[31] = (MIREQUESTRAMREADDATA[31] !== 1'bz) && MIREQUESTRAMREADDATA_delay[31]; // rv 0
  assign MIREQUESTRAMREADDATA_in[32] = (MIREQUESTRAMREADDATA[32] !== 1'bz) && MIREQUESTRAMREADDATA_delay[32]; // rv 0
  assign MIREQUESTRAMREADDATA_in[33] = (MIREQUESTRAMREADDATA[33] !== 1'bz) && MIREQUESTRAMREADDATA_delay[33]; // rv 0
  assign MIREQUESTRAMREADDATA_in[34] = (MIREQUESTRAMREADDATA[34] !== 1'bz) && MIREQUESTRAMREADDATA_delay[34]; // rv 0
  assign MIREQUESTRAMREADDATA_in[35] = (MIREQUESTRAMREADDATA[35] !== 1'bz) && MIREQUESTRAMREADDATA_delay[35]; // rv 0
  assign MIREQUESTRAMREADDATA_in[36] = (MIREQUESTRAMREADDATA[36] !== 1'bz) && MIREQUESTRAMREADDATA_delay[36]; // rv 0
  assign MIREQUESTRAMREADDATA_in[37] = (MIREQUESTRAMREADDATA[37] !== 1'bz) && MIREQUESTRAMREADDATA_delay[37]; // rv 0
  assign MIREQUESTRAMREADDATA_in[38] = (MIREQUESTRAMREADDATA[38] !== 1'bz) && MIREQUESTRAMREADDATA_delay[38]; // rv 0
  assign MIREQUESTRAMREADDATA_in[39] = (MIREQUESTRAMREADDATA[39] !== 1'bz) && MIREQUESTRAMREADDATA_delay[39]; // rv 0
  assign MIREQUESTRAMREADDATA_in[3] = (MIREQUESTRAMREADDATA[3] !== 1'bz) && MIREQUESTRAMREADDATA_delay[3]; // rv 0
  assign MIREQUESTRAMREADDATA_in[40] = (MIREQUESTRAMREADDATA[40] !== 1'bz) && MIREQUESTRAMREADDATA_delay[40]; // rv 0
  assign MIREQUESTRAMREADDATA_in[41] = (MIREQUESTRAMREADDATA[41] !== 1'bz) && MIREQUESTRAMREADDATA_delay[41]; // rv 0
  assign MIREQUESTRAMREADDATA_in[42] = (MIREQUESTRAMREADDATA[42] !== 1'bz) && MIREQUESTRAMREADDATA_delay[42]; // rv 0
  assign MIREQUESTRAMREADDATA_in[43] = (MIREQUESTRAMREADDATA[43] !== 1'bz) && MIREQUESTRAMREADDATA_delay[43]; // rv 0
  assign MIREQUESTRAMREADDATA_in[44] = (MIREQUESTRAMREADDATA[44] !== 1'bz) && MIREQUESTRAMREADDATA_delay[44]; // rv 0
  assign MIREQUESTRAMREADDATA_in[45] = (MIREQUESTRAMREADDATA[45] !== 1'bz) && MIREQUESTRAMREADDATA_delay[45]; // rv 0
  assign MIREQUESTRAMREADDATA_in[46] = (MIREQUESTRAMREADDATA[46] !== 1'bz) && MIREQUESTRAMREADDATA_delay[46]; // rv 0
  assign MIREQUESTRAMREADDATA_in[47] = (MIREQUESTRAMREADDATA[47] !== 1'bz) && MIREQUESTRAMREADDATA_delay[47]; // rv 0
  assign MIREQUESTRAMREADDATA_in[48] = (MIREQUESTRAMREADDATA[48] !== 1'bz) && MIREQUESTRAMREADDATA_delay[48]; // rv 0
  assign MIREQUESTRAMREADDATA_in[49] = (MIREQUESTRAMREADDATA[49] !== 1'bz) && MIREQUESTRAMREADDATA_delay[49]; // rv 0
  assign MIREQUESTRAMREADDATA_in[4] = (MIREQUESTRAMREADDATA[4] !== 1'bz) && MIREQUESTRAMREADDATA_delay[4]; // rv 0
  assign MIREQUESTRAMREADDATA_in[50] = (MIREQUESTRAMREADDATA[50] !== 1'bz) && MIREQUESTRAMREADDATA_delay[50]; // rv 0
  assign MIREQUESTRAMREADDATA_in[51] = (MIREQUESTRAMREADDATA[51] !== 1'bz) && MIREQUESTRAMREADDATA_delay[51]; // rv 0
  assign MIREQUESTRAMREADDATA_in[52] = (MIREQUESTRAMREADDATA[52] !== 1'bz) && MIREQUESTRAMREADDATA_delay[52]; // rv 0
  assign MIREQUESTRAMREADDATA_in[53] = (MIREQUESTRAMREADDATA[53] !== 1'bz) && MIREQUESTRAMREADDATA_delay[53]; // rv 0
  assign MIREQUESTRAMREADDATA_in[54] = (MIREQUESTRAMREADDATA[54] !== 1'bz) && MIREQUESTRAMREADDATA_delay[54]; // rv 0
  assign MIREQUESTRAMREADDATA_in[55] = (MIREQUESTRAMREADDATA[55] !== 1'bz) && MIREQUESTRAMREADDATA_delay[55]; // rv 0
  assign MIREQUESTRAMREADDATA_in[56] = (MIREQUESTRAMREADDATA[56] !== 1'bz) && MIREQUESTRAMREADDATA_delay[56]; // rv 0
  assign MIREQUESTRAMREADDATA_in[57] = (MIREQUESTRAMREADDATA[57] !== 1'bz) && MIREQUESTRAMREADDATA_delay[57]; // rv 0
  assign MIREQUESTRAMREADDATA_in[58] = (MIREQUESTRAMREADDATA[58] !== 1'bz) && MIREQUESTRAMREADDATA_delay[58]; // rv 0
  assign MIREQUESTRAMREADDATA_in[59] = (MIREQUESTRAMREADDATA[59] !== 1'bz) && MIREQUESTRAMREADDATA_delay[59]; // rv 0
  assign MIREQUESTRAMREADDATA_in[5] = (MIREQUESTRAMREADDATA[5] !== 1'bz) && MIREQUESTRAMREADDATA_delay[5]; // rv 0
  assign MIREQUESTRAMREADDATA_in[60] = (MIREQUESTRAMREADDATA[60] !== 1'bz) && MIREQUESTRAMREADDATA_delay[60]; // rv 0
  assign MIREQUESTRAMREADDATA_in[61] = (MIREQUESTRAMREADDATA[61] !== 1'bz) && MIREQUESTRAMREADDATA_delay[61]; // rv 0
  assign MIREQUESTRAMREADDATA_in[62] = (MIREQUESTRAMREADDATA[62] !== 1'bz) && MIREQUESTRAMREADDATA_delay[62]; // rv 0
  assign MIREQUESTRAMREADDATA_in[63] = (MIREQUESTRAMREADDATA[63] !== 1'bz) && MIREQUESTRAMREADDATA_delay[63]; // rv 0
  assign MIREQUESTRAMREADDATA_in[64] = (MIREQUESTRAMREADDATA[64] !== 1'bz) && MIREQUESTRAMREADDATA_delay[64]; // rv 0
  assign MIREQUESTRAMREADDATA_in[65] = (MIREQUESTRAMREADDATA[65] !== 1'bz) && MIREQUESTRAMREADDATA_delay[65]; // rv 0
  assign MIREQUESTRAMREADDATA_in[66] = (MIREQUESTRAMREADDATA[66] !== 1'bz) && MIREQUESTRAMREADDATA_delay[66]; // rv 0
  assign MIREQUESTRAMREADDATA_in[67] = (MIREQUESTRAMREADDATA[67] !== 1'bz) && MIREQUESTRAMREADDATA_delay[67]; // rv 0
  assign MIREQUESTRAMREADDATA_in[68] = (MIREQUESTRAMREADDATA[68] !== 1'bz) && MIREQUESTRAMREADDATA_delay[68]; // rv 0
  assign MIREQUESTRAMREADDATA_in[69] = (MIREQUESTRAMREADDATA[69] !== 1'bz) && MIREQUESTRAMREADDATA_delay[69]; // rv 0
  assign MIREQUESTRAMREADDATA_in[6] = (MIREQUESTRAMREADDATA[6] !== 1'bz) && MIREQUESTRAMREADDATA_delay[6]; // rv 0
  assign MIREQUESTRAMREADDATA_in[70] = (MIREQUESTRAMREADDATA[70] !== 1'bz) && MIREQUESTRAMREADDATA_delay[70]; // rv 0
  assign MIREQUESTRAMREADDATA_in[71] = (MIREQUESTRAMREADDATA[71] !== 1'bz) && MIREQUESTRAMREADDATA_delay[71]; // rv 0
  assign MIREQUESTRAMREADDATA_in[72] = (MIREQUESTRAMREADDATA[72] !== 1'bz) && MIREQUESTRAMREADDATA_delay[72]; // rv 0
  assign MIREQUESTRAMREADDATA_in[73] = (MIREQUESTRAMREADDATA[73] !== 1'bz) && MIREQUESTRAMREADDATA_delay[73]; // rv 0
  assign MIREQUESTRAMREADDATA_in[74] = (MIREQUESTRAMREADDATA[74] !== 1'bz) && MIREQUESTRAMREADDATA_delay[74]; // rv 0
  assign MIREQUESTRAMREADDATA_in[75] = (MIREQUESTRAMREADDATA[75] !== 1'bz) && MIREQUESTRAMREADDATA_delay[75]; // rv 0
  assign MIREQUESTRAMREADDATA_in[76] = (MIREQUESTRAMREADDATA[76] !== 1'bz) && MIREQUESTRAMREADDATA_delay[76]; // rv 0
  assign MIREQUESTRAMREADDATA_in[77] = (MIREQUESTRAMREADDATA[77] !== 1'bz) && MIREQUESTRAMREADDATA_delay[77]; // rv 0
  assign MIREQUESTRAMREADDATA_in[78] = (MIREQUESTRAMREADDATA[78] !== 1'bz) && MIREQUESTRAMREADDATA_delay[78]; // rv 0
  assign MIREQUESTRAMREADDATA_in[79] = (MIREQUESTRAMREADDATA[79] !== 1'bz) && MIREQUESTRAMREADDATA_delay[79]; // rv 0
  assign MIREQUESTRAMREADDATA_in[7] = (MIREQUESTRAMREADDATA[7] !== 1'bz) && MIREQUESTRAMREADDATA_delay[7]; // rv 0
  assign MIREQUESTRAMREADDATA_in[80] = (MIREQUESTRAMREADDATA[80] !== 1'bz) && MIREQUESTRAMREADDATA_delay[80]; // rv 0
  assign MIREQUESTRAMREADDATA_in[81] = (MIREQUESTRAMREADDATA[81] !== 1'bz) && MIREQUESTRAMREADDATA_delay[81]; // rv 0
  assign MIREQUESTRAMREADDATA_in[82] = (MIREQUESTRAMREADDATA[82] !== 1'bz) && MIREQUESTRAMREADDATA_delay[82]; // rv 0
  assign MIREQUESTRAMREADDATA_in[83] = (MIREQUESTRAMREADDATA[83] !== 1'bz) && MIREQUESTRAMREADDATA_delay[83]; // rv 0
  assign MIREQUESTRAMREADDATA_in[84] = (MIREQUESTRAMREADDATA[84] !== 1'bz) && MIREQUESTRAMREADDATA_delay[84]; // rv 0
  assign MIREQUESTRAMREADDATA_in[85] = (MIREQUESTRAMREADDATA[85] !== 1'bz) && MIREQUESTRAMREADDATA_delay[85]; // rv 0
  assign MIREQUESTRAMREADDATA_in[86] = (MIREQUESTRAMREADDATA[86] !== 1'bz) && MIREQUESTRAMREADDATA_delay[86]; // rv 0
  assign MIREQUESTRAMREADDATA_in[87] = (MIREQUESTRAMREADDATA[87] !== 1'bz) && MIREQUESTRAMREADDATA_delay[87]; // rv 0
  assign MIREQUESTRAMREADDATA_in[88] = (MIREQUESTRAMREADDATA[88] !== 1'bz) && MIREQUESTRAMREADDATA_delay[88]; // rv 0
  assign MIREQUESTRAMREADDATA_in[89] = (MIREQUESTRAMREADDATA[89] !== 1'bz) && MIREQUESTRAMREADDATA_delay[89]; // rv 0
  assign MIREQUESTRAMREADDATA_in[8] = (MIREQUESTRAMREADDATA[8] !== 1'bz) && MIREQUESTRAMREADDATA_delay[8]; // rv 0
  assign MIREQUESTRAMREADDATA_in[90] = (MIREQUESTRAMREADDATA[90] !== 1'bz) && MIREQUESTRAMREADDATA_delay[90]; // rv 0
  assign MIREQUESTRAMREADDATA_in[91] = (MIREQUESTRAMREADDATA[91] !== 1'bz) && MIREQUESTRAMREADDATA_delay[91]; // rv 0
  assign MIREQUESTRAMREADDATA_in[92] = (MIREQUESTRAMREADDATA[92] !== 1'bz) && MIREQUESTRAMREADDATA_delay[92]; // rv 0
  assign MIREQUESTRAMREADDATA_in[93] = (MIREQUESTRAMREADDATA[93] !== 1'bz) && MIREQUESTRAMREADDATA_delay[93]; // rv 0
  assign MIREQUESTRAMREADDATA_in[94] = (MIREQUESTRAMREADDATA[94] !== 1'bz) && MIREQUESTRAMREADDATA_delay[94]; // rv 0
  assign MIREQUESTRAMREADDATA_in[95] = (MIREQUESTRAMREADDATA[95] !== 1'bz) && MIREQUESTRAMREADDATA_delay[95]; // rv 0
  assign MIREQUESTRAMREADDATA_in[96] = (MIREQUESTRAMREADDATA[96] !== 1'bz) && MIREQUESTRAMREADDATA_delay[96]; // rv 0
  assign MIREQUESTRAMREADDATA_in[97] = (MIREQUESTRAMREADDATA[97] !== 1'bz) && MIREQUESTRAMREADDATA_delay[97]; // rv 0
  assign MIREQUESTRAMREADDATA_in[98] = (MIREQUESTRAMREADDATA[98] !== 1'bz) && MIREQUESTRAMREADDATA_delay[98]; // rv 0
  assign MIREQUESTRAMREADDATA_in[99] = (MIREQUESTRAMREADDATA[99] !== 1'bz) && MIREQUESTRAMREADDATA_delay[99]; // rv 0
  assign MIREQUESTRAMREADDATA_in[9] = (MIREQUESTRAMREADDATA[9] !== 1'bz) && MIREQUESTRAMREADDATA_delay[9]; // rv 0
  assign PCIECQNPREQ_in = (PCIECQNPREQ === 1'bz) || PCIECQNPREQ_delay; // rv 1
  assign PIPECLK_in = (PIPECLK !== 1'bz) && PIPECLK_delay; // rv 0
  assign PIPEEQFS_in[0] = (PIPEEQFS[0] !== 1'bz) && PIPEEQFS_delay[0]; // rv 0
  assign PIPEEQFS_in[1] = (PIPEEQFS[1] !== 1'bz) && PIPEEQFS_delay[1]; // rv 0
  assign PIPEEQFS_in[2] = (PIPEEQFS[2] !== 1'bz) && PIPEEQFS_delay[2]; // rv 0
  assign PIPEEQFS_in[3] = (PIPEEQFS[3] !== 1'bz) && PIPEEQFS_delay[3]; // rv 0
  assign PIPEEQFS_in[4] = (PIPEEQFS[4] !== 1'bz) && PIPEEQFS_delay[4]; // rv 0
  assign PIPEEQFS_in[5] = (PIPEEQFS[5] !== 1'bz) && PIPEEQFS_delay[5]; // rv 0
  assign PIPEEQLF_in[0] = (PIPEEQLF[0] !== 1'bz) && PIPEEQLF_delay[0]; // rv 0
  assign PIPEEQLF_in[1] = (PIPEEQLF[1] !== 1'bz) && PIPEEQLF_delay[1]; // rv 0
  assign PIPEEQLF_in[2] = (PIPEEQLF[2] !== 1'bz) && PIPEEQLF_delay[2]; // rv 0
  assign PIPEEQLF_in[3] = (PIPEEQLF[3] !== 1'bz) && PIPEEQLF_delay[3]; // rv 0
  assign PIPEEQLF_in[4] = (PIPEEQLF[4] !== 1'bz) && PIPEEQLF_delay[4]; // rv 0
  assign PIPEEQLF_in[5] = (PIPEEQLF[5] !== 1'bz) && PIPEEQLF_delay[5]; // rv 0
  assign PIPERESETN_in = (PIPERESETN !== 1'bz) && PIPERESETN_delay; // rv 0
  assign PIPERX0CHARISK_in[0] = (PIPERX0CHARISK[0] === 1'bz) || PIPERX0CHARISK_delay[0]; // rv 1
  assign PIPERX0CHARISK_in[1] = (PIPERX0CHARISK[1] === 1'bz) || PIPERX0CHARISK_delay[1]; // rv 1
  assign PIPERX0DATAVALID_in = (PIPERX0DATAVALID !== 1'bz) && PIPERX0DATAVALID_delay; // rv 0
  assign PIPERX0DATA_in[0] = (PIPERX0DATA[0] !== 1'bz) && PIPERX0DATA_delay[0]; // rv 0
  assign PIPERX0DATA_in[10] = (PIPERX0DATA[10] !== 1'bz) && PIPERX0DATA_delay[10]; // rv 0
  assign PIPERX0DATA_in[11] = (PIPERX0DATA[11] !== 1'bz) && PIPERX0DATA_delay[11]; // rv 0
  assign PIPERX0DATA_in[12] = (PIPERX0DATA[12] !== 1'bz) && PIPERX0DATA_delay[12]; // rv 0
  assign PIPERX0DATA_in[13] = (PIPERX0DATA[13] !== 1'bz) && PIPERX0DATA_delay[13]; // rv 0
  assign PIPERX0DATA_in[14] = (PIPERX0DATA[14] !== 1'bz) && PIPERX0DATA_delay[14]; // rv 0
  assign PIPERX0DATA_in[15] = (PIPERX0DATA[15] !== 1'bz) && PIPERX0DATA_delay[15]; // rv 0
  assign PIPERX0DATA_in[16] = (PIPERX0DATA[16] !== 1'bz) && PIPERX0DATA_delay[16]; // rv 0
  assign PIPERX0DATA_in[17] = (PIPERX0DATA[17] !== 1'bz) && PIPERX0DATA_delay[17]; // rv 0
  assign PIPERX0DATA_in[18] = (PIPERX0DATA[18] !== 1'bz) && PIPERX0DATA_delay[18]; // rv 0
  assign PIPERX0DATA_in[19] = (PIPERX0DATA[19] !== 1'bz) && PIPERX0DATA_delay[19]; // rv 0
  assign PIPERX0DATA_in[1] = (PIPERX0DATA[1] !== 1'bz) && PIPERX0DATA_delay[1]; // rv 0
  assign PIPERX0DATA_in[20] = (PIPERX0DATA[20] !== 1'bz) && PIPERX0DATA_delay[20]; // rv 0
  assign PIPERX0DATA_in[21] = (PIPERX0DATA[21] !== 1'bz) && PIPERX0DATA_delay[21]; // rv 0
  assign PIPERX0DATA_in[22] = (PIPERX0DATA[22] !== 1'bz) && PIPERX0DATA_delay[22]; // rv 0
  assign PIPERX0DATA_in[23] = (PIPERX0DATA[23] !== 1'bz) && PIPERX0DATA_delay[23]; // rv 0
  assign PIPERX0DATA_in[24] = (PIPERX0DATA[24] !== 1'bz) && PIPERX0DATA_delay[24]; // rv 0
  assign PIPERX0DATA_in[25] = (PIPERX0DATA[25] !== 1'bz) && PIPERX0DATA_delay[25]; // rv 0
  assign PIPERX0DATA_in[26] = (PIPERX0DATA[26] !== 1'bz) && PIPERX0DATA_delay[26]; // rv 0
  assign PIPERX0DATA_in[27] = (PIPERX0DATA[27] !== 1'bz) && PIPERX0DATA_delay[27]; // rv 0
  assign PIPERX0DATA_in[28] = (PIPERX0DATA[28] !== 1'bz) && PIPERX0DATA_delay[28]; // rv 0
  assign PIPERX0DATA_in[29] = (PIPERX0DATA[29] !== 1'bz) && PIPERX0DATA_delay[29]; // rv 0
  assign PIPERX0DATA_in[2] = (PIPERX0DATA[2] !== 1'bz) && PIPERX0DATA_delay[2]; // rv 0
  assign PIPERX0DATA_in[30] = (PIPERX0DATA[30] !== 1'bz) && PIPERX0DATA_delay[30]; // rv 0
  assign PIPERX0DATA_in[31] = (PIPERX0DATA[31] !== 1'bz) && PIPERX0DATA_delay[31]; // rv 0
  assign PIPERX0DATA_in[3] = (PIPERX0DATA[3] !== 1'bz) && PIPERX0DATA_delay[3]; // rv 0
  assign PIPERX0DATA_in[4] = (PIPERX0DATA[4] !== 1'bz) && PIPERX0DATA_delay[4]; // rv 0
  assign PIPERX0DATA_in[5] = (PIPERX0DATA[5] !== 1'bz) && PIPERX0DATA_delay[5]; // rv 0
  assign PIPERX0DATA_in[6] = (PIPERX0DATA[6] !== 1'bz) && PIPERX0DATA_delay[6]; // rv 0
  assign PIPERX0DATA_in[7] = (PIPERX0DATA[7] !== 1'bz) && PIPERX0DATA_delay[7]; // rv 0
  assign PIPERX0DATA_in[8] = (PIPERX0DATA[8] !== 1'bz) && PIPERX0DATA_delay[8]; // rv 0
  assign PIPERX0DATA_in[9] = (PIPERX0DATA[9] !== 1'bz) && PIPERX0DATA_delay[9]; // rv 0
  assign PIPERX0ELECIDLE_in = (PIPERX0ELECIDLE === 1'bz) || PIPERX0ELECIDLE_delay; // rv 1
  assign PIPERX0EQDONE_in = (PIPERX0EQDONE !== 1'bz) && PIPERX0EQDONE_delay; // rv 0
  assign PIPERX0EQLPADAPTDONE_in = (PIPERX0EQLPADAPTDONE !== 1'bz) && PIPERX0EQLPADAPTDONE_delay; // rv 0
  assign PIPERX0EQLPLFFSSEL_in = (PIPERX0EQLPLFFSSEL !== 1'bz) && PIPERX0EQLPLFFSSEL_delay; // rv 0
  assign PIPERX0EQLPNEWTXCOEFFORPRESET_in[0] = (PIPERX0EQLPNEWTXCOEFFORPRESET[0] !== 1'bz) && PIPERX0EQLPNEWTXCOEFFORPRESET_delay[0]; // rv 0
  assign PIPERX0EQLPNEWTXCOEFFORPRESET_in[10] = (PIPERX0EQLPNEWTXCOEFFORPRESET[10] !== 1'bz) && PIPERX0EQLPNEWTXCOEFFORPRESET_delay[10]; // rv 0
  assign PIPERX0EQLPNEWTXCOEFFORPRESET_in[11] = (PIPERX0EQLPNEWTXCOEFFORPRESET[11] !== 1'bz) && PIPERX0EQLPNEWTXCOEFFORPRESET_delay[11]; // rv 0
  assign PIPERX0EQLPNEWTXCOEFFORPRESET_in[12] = (PIPERX0EQLPNEWTXCOEFFORPRESET[12] !== 1'bz) && PIPERX0EQLPNEWTXCOEFFORPRESET_delay[12]; // rv 0
  assign PIPERX0EQLPNEWTXCOEFFORPRESET_in[13] = (PIPERX0EQLPNEWTXCOEFFORPRESET[13] !== 1'bz) && PIPERX0EQLPNEWTXCOEFFORPRESET_delay[13]; // rv 0
  assign PIPERX0EQLPNEWTXCOEFFORPRESET_in[14] = (PIPERX0EQLPNEWTXCOEFFORPRESET[14] !== 1'bz) && PIPERX0EQLPNEWTXCOEFFORPRESET_delay[14]; // rv 0
  assign PIPERX0EQLPNEWTXCOEFFORPRESET_in[15] = (PIPERX0EQLPNEWTXCOEFFORPRESET[15] !== 1'bz) && PIPERX0EQLPNEWTXCOEFFORPRESET_delay[15]; // rv 0
  assign PIPERX0EQLPNEWTXCOEFFORPRESET_in[16] = (PIPERX0EQLPNEWTXCOEFFORPRESET[16] !== 1'bz) && PIPERX0EQLPNEWTXCOEFFORPRESET_delay[16]; // rv 0
  assign PIPERX0EQLPNEWTXCOEFFORPRESET_in[17] = (PIPERX0EQLPNEWTXCOEFFORPRESET[17] !== 1'bz) && PIPERX0EQLPNEWTXCOEFFORPRESET_delay[17]; // rv 0
  assign PIPERX0EQLPNEWTXCOEFFORPRESET_in[1] = (PIPERX0EQLPNEWTXCOEFFORPRESET[1] !== 1'bz) && PIPERX0EQLPNEWTXCOEFFORPRESET_delay[1]; // rv 0
  assign PIPERX0EQLPNEWTXCOEFFORPRESET_in[2] = (PIPERX0EQLPNEWTXCOEFFORPRESET[2] !== 1'bz) && PIPERX0EQLPNEWTXCOEFFORPRESET_delay[2]; // rv 0
  assign PIPERX0EQLPNEWTXCOEFFORPRESET_in[3] = (PIPERX0EQLPNEWTXCOEFFORPRESET[3] !== 1'bz) && PIPERX0EQLPNEWTXCOEFFORPRESET_delay[3]; // rv 0
  assign PIPERX0EQLPNEWTXCOEFFORPRESET_in[4] = (PIPERX0EQLPNEWTXCOEFFORPRESET[4] !== 1'bz) && PIPERX0EQLPNEWTXCOEFFORPRESET_delay[4]; // rv 0
  assign PIPERX0EQLPNEWTXCOEFFORPRESET_in[5] = (PIPERX0EQLPNEWTXCOEFFORPRESET[5] !== 1'bz) && PIPERX0EQLPNEWTXCOEFFORPRESET_delay[5]; // rv 0
  assign PIPERX0EQLPNEWTXCOEFFORPRESET_in[6] = (PIPERX0EQLPNEWTXCOEFFORPRESET[6] !== 1'bz) && PIPERX0EQLPNEWTXCOEFFORPRESET_delay[6]; // rv 0
  assign PIPERX0EQLPNEWTXCOEFFORPRESET_in[7] = (PIPERX0EQLPNEWTXCOEFFORPRESET[7] !== 1'bz) && PIPERX0EQLPNEWTXCOEFFORPRESET_delay[7]; // rv 0
  assign PIPERX0EQLPNEWTXCOEFFORPRESET_in[8] = (PIPERX0EQLPNEWTXCOEFFORPRESET[8] !== 1'bz) && PIPERX0EQLPNEWTXCOEFFORPRESET_delay[8]; // rv 0
  assign PIPERX0EQLPNEWTXCOEFFORPRESET_in[9] = (PIPERX0EQLPNEWTXCOEFFORPRESET[9] !== 1'bz) && PIPERX0EQLPNEWTXCOEFFORPRESET_delay[9]; // rv 0
  assign PIPERX0PHYSTATUS_in = (PIPERX0PHYSTATUS === 1'bz) || PIPERX0PHYSTATUS_delay; // rv 1
  assign PIPERX0STARTBLOCK_in = (PIPERX0STARTBLOCK !== 1'bz) && PIPERX0STARTBLOCK_delay; // rv 0
  assign PIPERX0STATUS_in[0] = (PIPERX0STATUS[0] !== 1'bz) && PIPERX0STATUS_delay[0]; // rv 0
  assign PIPERX0STATUS_in[1] = (PIPERX0STATUS[1] !== 1'bz) && PIPERX0STATUS_delay[1]; // rv 0
  assign PIPERX0STATUS_in[2] = (PIPERX0STATUS[2] !== 1'bz) && PIPERX0STATUS_delay[2]; // rv 0
  assign PIPERX0SYNCHEADER_in[0] = (PIPERX0SYNCHEADER[0] !== 1'bz) && PIPERX0SYNCHEADER_delay[0]; // rv 0
  assign PIPERX0SYNCHEADER_in[1] = (PIPERX0SYNCHEADER[1] !== 1'bz) && PIPERX0SYNCHEADER_delay[1]; // rv 0
  assign PIPERX0VALID_in = (PIPERX0VALID !== 1'bz) && PIPERX0VALID_delay; // rv 0
  assign PIPERX1CHARISK_in[0] = (PIPERX1CHARISK[0] === 1'bz) || PIPERX1CHARISK_delay[0]; // rv 1
  assign PIPERX1CHARISK_in[1] = (PIPERX1CHARISK[1] === 1'bz) || PIPERX1CHARISK_delay[1]; // rv 1
  assign PIPERX1DATAVALID_in = (PIPERX1DATAVALID !== 1'bz) && PIPERX1DATAVALID_delay; // rv 0
  assign PIPERX1DATA_in[0] = (PIPERX1DATA[0] !== 1'bz) && PIPERX1DATA_delay[0]; // rv 0
  assign PIPERX1DATA_in[10] = (PIPERX1DATA[10] !== 1'bz) && PIPERX1DATA_delay[10]; // rv 0
  assign PIPERX1DATA_in[11] = (PIPERX1DATA[11] !== 1'bz) && PIPERX1DATA_delay[11]; // rv 0
  assign PIPERX1DATA_in[12] = (PIPERX1DATA[12] !== 1'bz) && PIPERX1DATA_delay[12]; // rv 0
  assign PIPERX1DATA_in[13] = (PIPERX1DATA[13] !== 1'bz) && PIPERX1DATA_delay[13]; // rv 0
  assign PIPERX1DATA_in[14] = (PIPERX1DATA[14] !== 1'bz) && PIPERX1DATA_delay[14]; // rv 0
  assign PIPERX1DATA_in[15] = (PIPERX1DATA[15] !== 1'bz) && PIPERX1DATA_delay[15]; // rv 0
  assign PIPERX1DATA_in[16] = (PIPERX1DATA[16] !== 1'bz) && PIPERX1DATA_delay[16]; // rv 0
  assign PIPERX1DATA_in[17] = (PIPERX1DATA[17] !== 1'bz) && PIPERX1DATA_delay[17]; // rv 0
  assign PIPERX1DATA_in[18] = (PIPERX1DATA[18] !== 1'bz) && PIPERX1DATA_delay[18]; // rv 0
  assign PIPERX1DATA_in[19] = (PIPERX1DATA[19] !== 1'bz) && PIPERX1DATA_delay[19]; // rv 0
  assign PIPERX1DATA_in[1] = (PIPERX1DATA[1] !== 1'bz) && PIPERX1DATA_delay[1]; // rv 0
  assign PIPERX1DATA_in[20] = (PIPERX1DATA[20] !== 1'bz) && PIPERX1DATA_delay[20]; // rv 0
  assign PIPERX1DATA_in[21] = (PIPERX1DATA[21] !== 1'bz) && PIPERX1DATA_delay[21]; // rv 0
  assign PIPERX1DATA_in[22] = (PIPERX1DATA[22] !== 1'bz) && PIPERX1DATA_delay[22]; // rv 0
  assign PIPERX1DATA_in[23] = (PIPERX1DATA[23] !== 1'bz) && PIPERX1DATA_delay[23]; // rv 0
  assign PIPERX1DATA_in[24] = (PIPERX1DATA[24] !== 1'bz) && PIPERX1DATA_delay[24]; // rv 0
  assign PIPERX1DATA_in[25] = (PIPERX1DATA[25] !== 1'bz) && PIPERX1DATA_delay[25]; // rv 0
  assign PIPERX1DATA_in[26] = (PIPERX1DATA[26] !== 1'bz) && PIPERX1DATA_delay[26]; // rv 0
  assign PIPERX1DATA_in[27] = (PIPERX1DATA[27] !== 1'bz) && PIPERX1DATA_delay[27]; // rv 0
  assign PIPERX1DATA_in[28] = (PIPERX1DATA[28] !== 1'bz) && PIPERX1DATA_delay[28]; // rv 0
  assign PIPERX1DATA_in[29] = (PIPERX1DATA[29] !== 1'bz) && PIPERX1DATA_delay[29]; // rv 0
  assign PIPERX1DATA_in[2] = (PIPERX1DATA[2] !== 1'bz) && PIPERX1DATA_delay[2]; // rv 0
  assign PIPERX1DATA_in[30] = (PIPERX1DATA[30] !== 1'bz) && PIPERX1DATA_delay[30]; // rv 0
  assign PIPERX1DATA_in[31] = (PIPERX1DATA[31] !== 1'bz) && PIPERX1DATA_delay[31]; // rv 0
  assign PIPERX1DATA_in[3] = (PIPERX1DATA[3] !== 1'bz) && PIPERX1DATA_delay[3]; // rv 0
  assign PIPERX1DATA_in[4] = (PIPERX1DATA[4] !== 1'bz) && PIPERX1DATA_delay[4]; // rv 0
  assign PIPERX1DATA_in[5] = (PIPERX1DATA[5] !== 1'bz) && PIPERX1DATA_delay[5]; // rv 0
  assign PIPERX1DATA_in[6] = (PIPERX1DATA[6] !== 1'bz) && PIPERX1DATA_delay[6]; // rv 0
  assign PIPERX1DATA_in[7] = (PIPERX1DATA[7] !== 1'bz) && PIPERX1DATA_delay[7]; // rv 0
  assign PIPERX1DATA_in[8] = (PIPERX1DATA[8] !== 1'bz) && PIPERX1DATA_delay[8]; // rv 0
  assign PIPERX1DATA_in[9] = (PIPERX1DATA[9] !== 1'bz) && PIPERX1DATA_delay[9]; // rv 0
  assign PIPERX1ELECIDLE_in = (PIPERX1ELECIDLE === 1'bz) || PIPERX1ELECIDLE_delay; // rv 1
  assign PIPERX1EQDONE_in = (PIPERX1EQDONE !== 1'bz) && PIPERX1EQDONE_delay; // rv 0
  assign PIPERX1EQLPADAPTDONE_in = (PIPERX1EQLPADAPTDONE !== 1'bz) && PIPERX1EQLPADAPTDONE_delay; // rv 0
  assign PIPERX1EQLPLFFSSEL_in = (PIPERX1EQLPLFFSSEL !== 1'bz) && PIPERX1EQLPLFFSSEL_delay; // rv 0
  assign PIPERX1EQLPNEWTXCOEFFORPRESET_in[0] = (PIPERX1EQLPNEWTXCOEFFORPRESET[0] !== 1'bz) && PIPERX1EQLPNEWTXCOEFFORPRESET_delay[0]; // rv 0
  assign PIPERX1EQLPNEWTXCOEFFORPRESET_in[10] = (PIPERX1EQLPNEWTXCOEFFORPRESET[10] !== 1'bz) && PIPERX1EQLPNEWTXCOEFFORPRESET_delay[10]; // rv 0
  assign PIPERX1EQLPNEWTXCOEFFORPRESET_in[11] = (PIPERX1EQLPNEWTXCOEFFORPRESET[11] !== 1'bz) && PIPERX1EQLPNEWTXCOEFFORPRESET_delay[11]; // rv 0
  assign PIPERX1EQLPNEWTXCOEFFORPRESET_in[12] = (PIPERX1EQLPNEWTXCOEFFORPRESET[12] !== 1'bz) && PIPERX1EQLPNEWTXCOEFFORPRESET_delay[12]; // rv 0
  assign PIPERX1EQLPNEWTXCOEFFORPRESET_in[13] = (PIPERX1EQLPNEWTXCOEFFORPRESET[13] !== 1'bz) && PIPERX1EQLPNEWTXCOEFFORPRESET_delay[13]; // rv 0
  assign PIPERX1EQLPNEWTXCOEFFORPRESET_in[14] = (PIPERX1EQLPNEWTXCOEFFORPRESET[14] !== 1'bz) && PIPERX1EQLPNEWTXCOEFFORPRESET_delay[14]; // rv 0
  assign PIPERX1EQLPNEWTXCOEFFORPRESET_in[15] = (PIPERX1EQLPNEWTXCOEFFORPRESET[15] !== 1'bz) && PIPERX1EQLPNEWTXCOEFFORPRESET_delay[15]; // rv 0
  assign PIPERX1EQLPNEWTXCOEFFORPRESET_in[16] = (PIPERX1EQLPNEWTXCOEFFORPRESET[16] !== 1'bz) && PIPERX1EQLPNEWTXCOEFFORPRESET_delay[16]; // rv 0
  assign PIPERX1EQLPNEWTXCOEFFORPRESET_in[17] = (PIPERX1EQLPNEWTXCOEFFORPRESET[17] !== 1'bz) && PIPERX1EQLPNEWTXCOEFFORPRESET_delay[17]; // rv 0
  assign PIPERX1EQLPNEWTXCOEFFORPRESET_in[1] = (PIPERX1EQLPNEWTXCOEFFORPRESET[1] !== 1'bz) && PIPERX1EQLPNEWTXCOEFFORPRESET_delay[1]; // rv 0
  assign PIPERX1EQLPNEWTXCOEFFORPRESET_in[2] = (PIPERX1EQLPNEWTXCOEFFORPRESET[2] !== 1'bz) && PIPERX1EQLPNEWTXCOEFFORPRESET_delay[2]; // rv 0
  assign PIPERX1EQLPNEWTXCOEFFORPRESET_in[3] = (PIPERX1EQLPNEWTXCOEFFORPRESET[3] !== 1'bz) && PIPERX1EQLPNEWTXCOEFFORPRESET_delay[3]; // rv 0
  assign PIPERX1EQLPNEWTXCOEFFORPRESET_in[4] = (PIPERX1EQLPNEWTXCOEFFORPRESET[4] !== 1'bz) && PIPERX1EQLPNEWTXCOEFFORPRESET_delay[4]; // rv 0
  assign PIPERX1EQLPNEWTXCOEFFORPRESET_in[5] = (PIPERX1EQLPNEWTXCOEFFORPRESET[5] !== 1'bz) && PIPERX1EQLPNEWTXCOEFFORPRESET_delay[5]; // rv 0
  assign PIPERX1EQLPNEWTXCOEFFORPRESET_in[6] = (PIPERX1EQLPNEWTXCOEFFORPRESET[6] !== 1'bz) && PIPERX1EQLPNEWTXCOEFFORPRESET_delay[6]; // rv 0
  assign PIPERX1EQLPNEWTXCOEFFORPRESET_in[7] = (PIPERX1EQLPNEWTXCOEFFORPRESET[7] !== 1'bz) && PIPERX1EQLPNEWTXCOEFFORPRESET_delay[7]; // rv 0
  assign PIPERX1EQLPNEWTXCOEFFORPRESET_in[8] = (PIPERX1EQLPNEWTXCOEFFORPRESET[8] !== 1'bz) && PIPERX1EQLPNEWTXCOEFFORPRESET_delay[8]; // rv 0
  assign PIPERX1EQLPNEWTXCOEFFORPRESET_in[9] = (PIPERX1EQLPNEWTXCOEFFORPRESET[9] !== 1'bz) && PIPERX1EQLPNEWTXCOEFFORPRESET_delay[9]; // rv 0
  assign PIPERX1PHYSTATUS_in = (PIPERX1PHYSTATUS === 1'bz) || PIPERX1PHYSTATUS_delay; // rv 1
  assign PIPERX1STARTBLOCK_in = (PIPERX1STARTBLOCK !== 1'bz) && PIPERX1STARTBLOCK_delay; // rv 0
  assign PIPERX1STATUS_in[0] = (PIPERX1STATUS[0] !== 1'bz) && PIPERX1STATUS_delay[0]; // rv 0
  assign PIPERX1STATUS_in[1] = (PIPERX1STATUS[1] !== 1'bz) && PIPERX1STATUS_delay[1]; // rv 0
  assign PIPERX1STATUS_in[2] = (PIPERX1STATUS[2] !== 1'bz) && PIPERX1STATUS_delay[2]; // rv 0
  assign PIPERX1SYNCHEADER_in[0] = (PIPERX1SYNCHEADER[0] !== 1'bz) && PIPERX1SYNCHEADER_delay[0]; // rv 0
  assign PIPERX1SYNCHEADER_in[1] = (PIPERX1SYNCHEADER[1] !== 1'bz) && PIPERX1SYNCHEADER_delay[1]; // rv 0
  assign PIPERX1VALID_in = (PIPERX1VALID !== 1'bz) && PIPERX1VALID_delay; // rv 0
  assign PIPERX2CHARISK_in[0] = (PIPERX2CHARISK[0] === 1'bz) || PIPERX2CHARISK_delay[0]; // rv 1
  assign PIPERX2CHARISK_in[1] = (PIPERX2CHARISK[1] === 1'bz) || PIPERX2CHARISK_delay[1]; // rv 1
  assign PIPERX2DATAVALID_in = (PIPERX2DATAVALID !== 1'bz) && PIPERX2DATAVALID_delay; // rv 0
  assign PIPERX2DATA_in[0] = (PIPERX2DATA[0] !== 1'bz) && PIPERX2DATA_delay[0]; // rv 0
  assign PIPERX2DATA_in[10] = (PIPERX2DATA[10] !== 1'bz) && PIPERX2DATA_delay[10]; // rv 0
  assign PIPERX2DATA_in[11] = (PIPERX2DATA[11] !== 1'bz) && PIPERX2DATA_delay[11]; // rv 0
  assign PIPERX2DATA_in[12] = (PIPERX2DATA[12] !== 1'bz) && PIPERX2DATA_delay[12]; // rv 0
  assign PIPERX2DATA_in[13] = (PIPERX2DATA[13] !== 1'bz) && PIPERX2DATA_delay[13]; // rv 0
  assign PIPERX2DATA_in[14] = (PIPERX2DATA[14] !== 1'bz) && PIPERX2DATA_delay[14]; // rv 0
  assign PIPERX2DATA_in[15] = (PIPERX2DATA[15] !== 1'bz) && PIPERX2DATA_delay[15]; // rv 0
  assign PIPERX2DATA_in[16] = (PIPERX2DATA[16] !== 1'bz) && PIPERX2DATA_delay[16]; // rv 0
  assign PIPERX2DATA_in[17] = (PIPERX2DATA[17] !== 1'bz) && PIPERX2DATA_delay[17]; // rv 0
  assign PIPERX2DATA_in[18] = (PIPERX2DATA[18] !== 1'bz) && PIPERX2DATA_delay[18]; // rv 0
  assign PIPERX2DATA_in[19] = (PIPERX2DATA[19] !== 1'bz) && PIPERX2DATA_delay[19]; // rv 0
  assign PIPERX2DATA_in[1] = (PIPERX2DATA[1] !== 1'bz) && PIPERX2DATA_delay[1]; // rv 0
  assign PIPERX2DATA_in[20] = (PIPERX2DATA[20] !== 1'bz) && PIPERX2DATA_delay[20]; // rv 0
  assign PIPERX2DATA_in[21] = (PIPERX2DATA[21] !== 1'bz) && PIPERX2DATA_delay[21]; // rv 0
  assign PIPERX2DATA_in[22] = (PIPERX2DATA[22] !== 1'bz) && PIPERX2DATA_delay[22]; // rv 0
  assign PIPERX2DATA_in[23] = (PIPERX2DATA[23] !== 1'bz) && PIPERX2DATA_delay[23]; // rv 0
  assign PIPERX2DATA_in[24] = (PIPERX2DATA[24] !== 1'bz) && PIPERX2DATA_delay[24]; // rv 0
  assign PIPERX2DATA_in[25] = (PIPERX2DATA[25] !== 1'bz) && PIPERX2DATA_delay[25]; // rv 0
  assign PIPERX2DATA_in[26] = (PIPERX2DATA[26] !== 1'bz) && PIPERX2DATA_delay[26]; // rv 0
  assign PIPERX2DATA_in[27] = (PIPERX2DATA[27] !== 1'bz) && PIPERX2DATA_delay[27]; // rv 0
  assign PIPERX2DATA_in[28] = (PIPERX2DATA[28] !== 1'bz) && PIPERX2DATA_delay[28]; // rv 0
  assign PIPERX2DATA_in[29] = (PIPERX2DATA[29] !== 1'bz) && PIPERX2DATA_delay[29]; // rv 0
  assign PIPERX2DATA_in[2] = (PIPERX2DATA[2] !== 1'bz) && PIPERX2DATA_delay[2]; // rv 0
  assign PIPERX2DATA_in[30] = (PIPERX2DATA[30] !== 1'bz) && PIPERX2DATA_delay[30]; // rv 0
  assign PIPERX2DATA_in[31] = (PIPERX2DATA[31] !== 1'bz) && PIPERX2DATA_delay[31]; // rv 0
  assign PIPERX2DATA_in[3] = (PIPERX2DATA[3] !== 1'bz) && PIPERX2DATA_delay[3]; // rv 0
  assign PIPERX2DATA_in[4] = (PIPERX2DATA[4] !== 1'bz) && PIPERX2DATA_delay[4]; // rv 0
  assign PIPERX2DATA_in[5] = (PIPERX2DATA[5] !== 1'bz) && PIPERX2DATA_delay[5]; // rv 0
  assign PIPERX2DATA_in[6] = (PIPERX2DATA[6] !== 1'bz) && PIPERX2DATA_delay[6]; // rv 0
  assign PIPERX2DATA_in[7] = (PIPERX2DATA[7] !== 1'bz) && PIPERX2DATA_delay[7]; // rv 0
  assign PIPERX2DATA_in[8] = (PIPERX2DATA[8] !== 1'bz) && PIPERX2DATA_delay[8]; // rv 0
  assign PIPERX2DATA_in[9] = (PIPERX2DATA[9] !== 1'bz) && PIPERX2DATA_delay[9]; // rv 0
  assign PIPERX2ELECIDLE_in = (PIPERX2ELECIDLE === 1'bz) || PIPERX2ELECIDLE_delay; // rv 1
  assign PIPERX2EQDONE_in = (PIPERX2EQDONE !== 1'bz) && PIPERX2EQDONE_delay; // rv 0
  assign PIPERX2EQLPADAPTDONE_in = (PIPERX2EQLPADAPTDONE !== 1'bz) && PIPERX2EQLPADAPTDONE_delay; // rv 0
  assign PIPERX2EQLPLFFSSEL_in = (PIPERX2EQLPLFFSSEL !== 1'bz) && PIPERX2EQLPLFFSSEL_delay; // rv 0
  assign PIPERX2EQLPNEWTXCOEFFORPRESET_in[0] = (PIPERX2EQLPNEWTXCOEFFORPRESET[0] !== 1'bz) && PIPERX2EQLPNEWTXCOEFFORPRESET_delay[0]; // rv 0
  assign PIPERX2EQLPNEWTXCOEFFORPRESET_in[10] = (PIPERX2EQLPNEWTXCOEFFORPRESET[10] !== 1'bz) && PIPERX2EQLPNEWTXCOEFFORPRESET_delay[10]; // rv 0
  assign PIPERX2EQLPNEWTXCOEFFORPRESET_in[11] = (PIPERX2EQLPNEWTXCOEFFORPRESET[11] !== 1'bz) && PIPERX2EQLPNEWTXCOEFFORPRESET_delay[11]; // rv 0
  assign PIPERX2EQLPNEWTXCOEFFORPRESET_in[12] = (PIPERX2EQLPNEWTXCOEFFORPRESET[12] !== 1'bz) && PIPERX2EQLPNEWTXCOEFFORPRESET_delay[12]; // rv 0
  assign PIPERX2EQLPNEWTXCOEFFORPRESET_in[13] = (PIPERX2EQLPNEWTXCOEFFORPRESET[13] !== 1'bz) && PIPERX2EQLPNEWTXCOEFFORPRESET_delay[13]; // rv 0
  assign PIPERX2EQLPNEWTXCOEFFORPRESET_in[14] = (PIPERX2EQLPNEWTXCOEFFORPRESET[14] !== 1'bz) && PIPERX2EQLPNEWTXCOEFFORPRESET_delay[14]; // rv 0
  assign PIPERX2EQLPNEWTXCOEFFORPRESET_in[15] = (PIPERX2EQLPNEWTXCOEFFORPRESET[15] !== 1'bz) && PIPERX2EQLPNEWTXCOEFFORPRESET_delay[15]; // rv 0
  assign PIPERX2EQLPNEWTXCOEFFORPRESET_in[16] = (PIPERX2EQLPNEWTXCOEFFORPRESET[16] !== 1'bz) && PIPERX2EQLPNEWTXCOEFFORPRESET_delay[16]; // rv 0
  assign PIPERX2EQLPNEWTXCOEFFORPRESET_in[17] = (PIPERX2EQLPNEWTXCOEFFORPRESET[17] !== 1'bz) && PIPERX2EQLPNEWTXCOEFFORPRESET_delay[17]; // rv 0
  assign PIPERX2EQLPNEWTXCOEFFORPRESET_in[1] = (PIPERX2EQLPNEWTXCOEFFORPRESET[1] !== 1'bz) && PIPERX2EQLPNEWTXCOEFFORPRESET_delay[1]; // rv 0
  assign PIPERX2EQLPNEWTXCOEFFORPRESET_in[2] = (PIPERX2EQLPNEWTXCOEFFORPRESET[2] !== 1'bz) && PIPERX2EQLPNEWTXCOEFFORPRESET_delay[2]; // rv 0
  assign PIPERX2EQLPNEWTXCOEFFORPRESET_in[3] = (PIPERX2EQLPNEWTXCOEFFORPRESET[3] !== 1'bz) && PIPERX2EQLPNEWTXCOEFFORPRESET_delay[3]; // rv 0
  assign PIPERX2EQLPNEWTXCOEFFORPRESET_in[4] = (PIPERX2EQLPNEWTXCOEFFORPRESET[4] !== 1'bz) && PIPERX2EQLPNEWTXCOEFFORPRESET_delay[4]; // rv 0
  assign PIPERX2EQLPNEWTXCOEFFORPRESET_in[5] = (PIPERX2EQLPNEWTXCOEFFORPRESET[5] !== 1'bz) && PIPERX2EQLPNEWTXCOEFFORPRESET_delay[5]; // rv 0
  assign PIPERX2EQLPNEWTXCOEFFORPRESET_in[6] = (PIPERX2EQLPNEWTXCOEFFORPRESET[6] !== 1'bz) && PIPERX2EQLPNEWTXCOEFFORPRESET_delay[6]; // rv 0
  assign PIPERX2EQLPNEWTXCOEFFORPRESET_in[7] = (PIPERX2EQLPNEWTXCOEFFORPRESET[7] !== 1'bz) && PIPERX2EQLPNEWTXCOEFFORPRESET_delay[7]; // rv 0
  assign PIPERX2EQLPNEWTXCOEFFORPRESET_in[8] = (PIPERX2EQLPNEWTXCOEFFORPRESET[8] !== 1'bz) && PIPERX2EQLPNEWTXCOEFFORPRESET_delay[8]; // rv 0
  assign PIPERX2EQLPNEWTXCOEFFORPRESET_in[9] = (PIPERX2EQLPNEWTXCOEFFORPRESET[9] !== 1'bz) && PIPERX2EQLPNEWTXCOEFFORPRESET_delay[9]; // rv 0
  assign PIPERX2PHYSTATUS_in = (PIPERX2PHYSTATUS === 1'bz) || PIPERX2PHYSTATUS_delay; // rv 1
  assign PIPERX2STARTBLOCK_in = (PIPERX2STARTBLOCK !== 1'bz) && PIPERX2STARTBLOCK_delay; // rv 0
  assign PIPERX2STATUS_in[0] = (PIPERX2STATUS[0] !== 1'bz) && PIPERX2STATUS_delay[0]; // rv 0
  assign PIPERX2STATUS_in[1] = (PIPERX2STATUS[1] !== 1'bz) && PIPERX2STATUS_delay[1]; // rv 0
  assign PIPERX2STATUS_in[2] = (PIPERX2STATUS[2] !== 1'bz) && PIPERX2STATUS_delay[2]; // rv 0
  assign PIPERX2SYNCHEADER_in[0] = (PIPERX2SYNCHEADER[0] !== 1'bz) && PIPERX2SYNCHEADER_delay[0]; // rv 0
  assign PIPERX2SYNCHEADER_in[1] = (PIPERX2SYNCHEADER[1] !== 1'bz) && PIPERX2SYNCHEADER_delay[1]; // rv 0
  assign PIPERX2VALID_in = (PIPERX2VALID !== 1'bz) && PIPERX2VALID_delay; // rv 0
  assign PIPERX3CHARISK_in[0] = (PIPERX3CHARISK[0] === 1'bz) || PIPERX3CHARISK_delay[0]; // rv 1
  assign PIPERX3CHARISK_in[1] = (PIPERX3CHARISK[1] === 1'bz) || PIPERX3CHARISK_delay[1]; // rv 1
  assign PIPERX3DATAVALID_in = (PIPERX3DATAVALID !== 1'bz) && PIPERX3DATAVALID_delay; // rv 0
  assign PIPERX3DATA_in[0] = (PIPERX3DATA[0] !== 1'bz) && PIPERX3DATA_delay[0]; // rv 0
  assign PIPERX3DATA_in[10] = (PIPERX3DATA[10] !== 1'bz) && PIPERX3DATA_delay[10]; // rv 0
  assign PIPERX3DATA_in[11] = (PIPERX3DATA[11] !== 1'bz) && PIPERX3DATA_delay[11]; // rv 0
  assign PIPERX3DATA_in[12] = (PIPERX3DATA[12] !== 1'bz) && PIPERX3DATA_delay[12]; // rv 0
  assign PIPERX3DATA_in[13] = (PIPERX3DATA[13] !== 1'bz) && PIPERX3DATA_delay[13]; // rv 0
  assign PIPERX3DATA_in[14] = (PIPERX3DATA[14] !== 1'bz) && PIPERX3DATA_delay[14]; // rv 0
  assign PIPERX3DATA_in[15] = (PIPERX3DATA[15] !== 1'bz) && PIPERX3DATA_delay[15]; // rv 0
  assign PIPERX3DATA_in[16] = (PIPERX3DATA[16] !== 1'bz) && PIPERX3DATA_delay[16]; // rv 0
  assign PIPERX3DATA_in[17] = (PIPERX3DATA[17] !== 1'bz) && PIPERX3DATA_delay[17]; // rv 0
  assign PIPERX3DATA_in[18] = (PIPERX3DATA[18] !== 1'bz) && PIPERX3DATA_delay[18]; // rv 0
  assign PIPERX3DATA_in[19] = (PIPERX3DATA[19] !== 1'bz) && PIPERX3DATA_delay[19]; // rv 0
  assign PIPERX3DATA_in[1] = (PIPERX3DATA[1] !== 1'bz) && PIPERX3DATA_delay[1]; // rv 0
  assign PIPERX3DATA_in[20] = (PIPERX3DATA[20] !== 1'bz) && PIPERX3DATA_delay[20]; // rv 0
  assign PIPERX3DATA_in[21] = (PIPERX3DATA[21] !== 1'bz) && PIPERX3DATA_delay[21]; // rv 0
  assign PIPERX3DATA_in[22] = (PIPERX3DATA[22] !== 1'bz) && PIPERX3DATA_delay[22]; // rv 0
  assign PIPERX3DATA_in[23] = (PIPERX3DATA[23] !== 1'bz) && PIPERX3DATA_delay[23]; // rv 0
  assign PIPERX3DATA_in[24] = (PIPERX3DATA[24] !== 1'bz) && PIPERX3DATA_delay[24]; // rv 0
  assign PIPERX3DATA_in[25] = (PIPERX3DATA[25] !== 1'bz) && PIPERX3DATA_delay[25]; // rv 0
  assign PIPERX3DATA_in[26] = (PIPERX3DATA[26] !== 1'bz) && PIPERX3DATA_delay[26]; // rv 0
  assign PIPERX3DATA_in[27] = (PIPERX3DATA[27] !== 1'bz) && PIPERX3DATA_delay[27]; // rv 0
  assign PIPERX3DATA_in[28] = (PIPERX3DATA[28] !== 1'bz) && PIPERX3DATA_delay[28]; // rv 0
  assign PIPERX3DATA_in[29] = (PIPERX3DATA[29] !== 1'bz) && PIPERX3DATA_delay[29]; // rv 0
  assign PIPERX3DATA_in[2] = (PIPERX3DATA[2] !== 1'bz) && PIPERX3DATA_delay[2]; // rv 0
  assign PIPERX3DATA_in[30] = (PIPERX3DATA[30] !== 1'bz) && PIPERX3DATA_delay[30]; // rv 0
  assign PIPERX3DATA_in[31] = (PIPERX3DATA[31] !== 1'bz) && PIPERX3DATA_delay[31]; // rv 0
  assign PIPERX3DATA_in[3] = (PIPERX3DATA[3] !== 1'bz) && PIPERX3DATA_delay[3]; // rv 0
  assign PIPERX3DATA_in[4] = (PIPERX3DATA[4] !== 1'bz) && PIPERX3DATA_delay[4]; // rv 0
  assign PIPERX3DATA_in[5] = (PIPERX3DATA[5] !== 1'bz) && PIPERX3DATA_delay[5]; // rv 0
  assign PIPERX3DATA_in[6] = (PIPERX3DATA[6] !== 1'bz) && PIPERX3DATA_delay[6]; // rv 0
  assign PIPERX3DATA_in[7] = (PIPERX3DATA[7] !== 1'bz) && PIPERX3DATA_delay[7]; // rv 0
  assign PIPERX3DATA_in[8] = (PIPERX3DATA[8] !== 1'bz) && PIPERX3DATA_delay[8]; // rv 0
  assign PIPERX3DATA_in[9] = (PIPERX3DATA[9] !== 1'bz) && PIPERX3DATA_delay[9]; // rv 0
  assign PIPERX3ELECIDLE_in = (PIPERX3ELECIDLE === 1'bz) || PIPERX3ELECIDLE_delay; // rv 1
  assign PIPERX3EQDONE_in = (PIPERX3EQDONE !== 1'bz) && PIPERX3EQDONE_delay; // rv 0
  assign PIPERX3EQLPADAPTDONE_in = (PIPERX3EQLPADAPTDONE !== 1'bz) && PIPERX3EQLPADAPTDONE_delay; // rv 0
  assign PIPERX3EQLPLFFSSEL_in = (PIPERX3EQLPLFFSSEL !== 1'bz) && PIPERX3EQLPLFFSSEL_delay; // rv 0
  assign PIPERX3EQLPNEWTXCOEFFORPRESET_in[0] = (PIPERX3EQLPNEWTXCOEFFORPRESET[0] !== 1'bz) && PIPERX3EQLPNEWTXCOEFFORPRESET_delay[0]; // rv 0
  assign PIPERX3EQLPNEWTXCOEFFORPRESET_in[10] = (PIPERX3EQLPNEWTXCOEFFORPRESET[10] !== 1'bz) && PIPERX3EQLPNEWTXCOEFFORPRESET_delay[10]; // rv 0
  assign PIPERX3EQLPNEWTXCOEFFORPRESET_in[11] = (PIPERX3EQLPNEWTXCOEFFORPRESET[11] !== 1'bz) && PIPERX3EQLPNEWTXCOEFFORPRESET_delay[11]; // rv 0
  assign PIPERX3EQLPNEWTXCOEFFORPRESET_in[12] = (PIPERX3EQLPNEWTXCOEFFORPRESET[12] !== 1'bz) && PIPERX3EQLPNEWTXCOEFFORPRESET_delay[12]; // rv 0
  assign PIPERX3EQLPNEWTXCOEFFORPRESET_in[13] = (PIPERX3EQLPNEWTXCOEFFORPRESET[13] !== 1'bz) && PIPERX3EQLPNEWTXCOEFFORPRESET_delay[13]; // rv 0
  assign PIPERX3EQLPNEWTXCOEFFORPRESET_in[14] = (PIPERX3EQLPNEWTXCOEFFORPRESET[14] !== 1'bz) && PIPERX3EQLPNEWTXCOEFFORPRESET_delay[14]; // rv 0
  assign PIPERX3EQLPNEWTXCOEFFORPRESET_in[15] = (PIPERX3EQLPNEWTXCOEFFORPRESET[15] !== 1'bz) && PIPERX3EQLPNEWTXCOEFFORPRESET_delay[15]; // rv 0
  assign PIPERX3EQLPNEWTXCOEFFORPRESET_in[16] = (PIPERX3EQLPNEWTXCOEFFORPRESET[16] !== 1'bz) && PIPERX3EQLPNEWTXCOEFFORPRESET_delay[16]; // rv 0
  assign PIPERX3EQLPNEWTXCOEFFORPRESET_in[17] = (PIPERX3EQLPNEWTXCOEFFORPRESET[17] !== 1'bz) && PIPERX3EQLPNEWTXCOEFFORPRESET_delay[17]; // rv 0
  assign PIPERX3EQLPNEWTXCOEFFORPRESET_in[1] = (PIPERX3EQLPNEWTXCOEFFORPRESET[1] !== 1'bz) && PIPERX3EQLPNEWTXCOEFFORPRESET_delay[1]; // rv 0
  assign PIPERX3EQLPNEWTXCOEFFORPRESET_in[2] = (PIPERX3EQLPNEWTXCOEFFORPRESET[2] !== 1'bz) && PIPERX3EQLPNEWTXCOEFFORPRESET_delay[2]; // rv 0
  assign PIPERX3EQLPNEWTXCOEFFORPRESET_in[3] = (PIPERX3EQLPNEWTXCOEFFORPRESET[3] !== 1'bz) && PIPERX3EQLPNEWTXCOEFFORPRESET_delay[3]; // rv 0
  assign PIPERX3EQLPNEWTXCOEFFORPRESET_in[4] = (PIPERX3EQLPNEWTXCOEFFORPRESET[4] !== 1'bz) && PIPERX3EQLPNEWTXCOEFFORPRESET_delay[4]; // rv 0
  assign PIPERX3EQLPNEWTXCOEFFORPRESET_in[5] = (PIPERX3EQLPNEWTXCOEFFORPRESET[5] !== 1'bz) && PIPERX3EQLPNEWTXCOEFFORPRESET_delay[5]; // rv 0
  assign PIPERX3EQLPNEWTXCOEFFORPRESET_in[6] = (PIPERX3EQLPNEWTXCOEFFORPRESET[6] !== 1'bz) && PIPERX3EQLPNEWTXCOEFFORPRESET_delay[6]; // rv 0
  assign PIPERX3EQLPNEWTXCOEFFORPRESET_in[7] = (PIPERX3EQLPNEWTXCOEFFORPRESET[7] !== 1'bz) && PIPERX3EQLPNEWTXCOEFFORPRESET_delay[7]; // rv 0
  assign PIPERX3EQLPNEWTXCOEFFORPRESET_in[8] = (PIPERX3EQLPNEWTXCOEFFORPRESET[8] !== 1'bz) && PIPERX3EQLPNEWTXCOEFFORPRESET_delay[8]; // rv 0
  assign PIPERX3EQLPNEWTXCOEFFORPRESET_in[9] = (PIPERX3EQLPNEWTXCOEFFORPRESET[9] !== 1'bz) && PIPERX3EQLPNEWTXCOEFFORPRESET_delay[9]; // rv 0
  assign PIPERX3PHYSTATUS_in = (PIPERX3PHYSTATUS === 1'bz) || PIPERX3PHYSTATUS_delay; // rv 1
  assign PIPERX3STARTBLOCK_in = (PIPERX3STARTBLOCK !== 1'bz) && PIPERX3STARTBLOCK_delay; // rv 0
  assign PIPERX3STATUS_in[0] = (PIPERX3STATUS[0] !== 1'bz) && PIPERX3STATUS_delay[0]; // rv 0
  assign PIPERX3STATUS_in[1] = (PIPERX3STATUS[1] !== 1'bz) && PIPERX3STATUS_delay[1]; // rv 0
  assign PIPERX3STATUS_in[2] = (PIPERX3STATUS[2] !== 1'bz) && PIPERX3STATUS_delay[2]; // rv 0
  assign PIPERX3SYNCHEADER_in[0] = (PIPERX3SYNCHEADER[0] !== 1'bz) && PIPERX3SYNCHEADER_delay[0]; // rv 0
  assign PIPERX3SYNCHEADER_in[1] = (PIPERX3SYNCHEADER[1] !== 1'bz) && PIPERX3SYNCHEADER_delay[1]; // rv 0
  assign PIPERX3VALID_in = (PIPERX3VALID !== 1'bz) && PIPERX3VALID_delay; // rv 0
  assign PIPERX4CHARISK_in[0] = (PIPERX4CHARISK[0] === 1'bz) || PIPERX4CHARISK_delay[0]; // rv 1
  assign PIPERX4CHARISK_in[1] = (PIPERX4CHARISK[1] === 1'bz) || PIPERX4CHARISK_delay[1]; // rv 1
  assign PIPERX4DATAVALID_in = (PIPERX4DATAVALID !== 1'bz) && PIPERX4DATAVALID_delay; // rv 0
  assign PIPERX4DATA_in[0] = (PIPERX4DATA[0] !== 1'bz) && PIPERX4DATA_delay[0]; // rv 0
  assign PIPERX4DATA_in[10] = (PIPERX4DATA[10] !== 1'bz) && PIPERX4DATA_delay[10]; // rv 0
  assign PIPERX4DATA_in[11] = (PIPERX4DATA[11] !== 1'bz) && PIPERX4DATA_delay[11]; // rv 0
  assign PIPERX4DATA_in[12] = (PIPERX4DATA[12] !== 1'bz) && PIPERX4DATA_delay[12]; // rv 0
  assign PIPERX4DATA_in[13] = (PIPERX4DATA[13] !== 1'bz) && PIPERX4DATA_delay[13]; // rv 0
  assign PIPERX4DATA_in[14] = (PIPERX4DATA[14] !== 1'bz) && PIPERX4DATA_delay[14]; // rv 0
  assign PIPERX4DATA_in[15] = (PIPERX4DATA[15] !== 1'bz) && PIPERX4DATA_delay[15]; // rv 0
  assign PIPERX4DATA_in[16] = (PIPERX4DATA[16] !== 1'bz) && PIPERX4DATA_delay[16]; // rv 0
  assign PIPERX4DATA_in[17] = (PIPERX4DATA[17] !== 1'bz) && PIPERX4DATA_delay[17]; // rv 0
  assign PIPERX4DATA_in[18] = (PIPERX4DATA[18] !== 1'bz) && PIPERX4DATA_delay[18]; // rv 0
  assign PIPERX4DATA_in[19] = (PIPERX4DATA[19] !== 1'bz) && PIPERX4DATA_delay[19]; // rv 0
  assign PIPERX4DATA_in[1] = (PIPERX4DATA[1] !== 1'bz) && PIPERX4DATA_delay[1]; // rv 0
  assign PIPERX4DATA_in[20] = (PIPERX4DATA[20] !== 1'bz) && PIPERX4DATA_delay[20]; // rv 0
  assign PIPERX4DATA_in[21] = (PIPERX4DATA[21] !== 1'bz) && PIPERX4DATA_delay[21]; // rv 0
  assign PIPERX4DATA_in[22] = (PIPERX4DATA[22] !== 1'bz) && PIPERX4DATA_delay[22]; // rv 0
  assign PIPERX4DATA_in[23] = (PIPERX4DATA[23] !== 1'bz) && PIPERX4DATA_delay[23]; // rv 0
  assign PIPERX4DATA_in[24] = (PIPERX4DATA[24] !== 1'bz) && PIPERX4DATA_delay[24]; // rv 0
  assign PIPERX4DATA_in[25] = (PIPERX4DATA[25] !== 1'bz) && PIPERX4DATA_delay[25]; // rv 0
  assign PIPERX4DATA_in[26] = (PIPERX4DATA[26] !== 1'bz) && PIPERX4DATA_delay[26]; // rv 0
  assign PIPERX4DATA_in[27] = (PIPERX4DATA[27] !== 1'bz) && PIPERX4DATA_delay[27]; // rv 0
  assign PIPERX4DATA_in[28] = (PIPERX4DATA[28] !== 1'bz) && PIPERX4DATA_delay[28]; // rv 0
  assign PIPERX4DATA_in[29] = (PIPERX4DATA[29] !== 1'bz) && PIPERX4DATA_delay[29]; // rv 0
  assign PIPERX4DATA_in[2] = (PIPERX4DATA[2] !== 1'bz) && PIPERX4DATA_delay[2]; // rv 0
  assign PIPERX4DATA_in[30] = (PIPERX4DATA[30] !== 1'bz) && PIPERX4DATA_delay[30]; // rv 0
  assign PIPERX4DATA_in[31] = (PIPERX4DATA[31] !== 1'bz) && PIPERX4DATA_delay[31]; // rv 0
  assign PIPERX4DATA_in[3] = (PIPERX4DATA[3] !== 1'bz) && PIPERX4DATA_delay[3]; // rv 0
  assign PIPERX4DATA_in[4] = (PIPERX4DATA[4] !== 1'bz) && PIPERX4DATA_delay[4]; // rv 0
  assign PIPERX4DATA_in[5] = (PIPERX4DATA[5] !== 1'bz) && PIPERX4DATA_delay[5]; // rv 0
  assign PIPERX4DATA_in[6] = (PIPERX4DATA[6] !== 1'bz) && PIPERX4DATA_delay[6]; // rv 0
  assign PIPERX4DATA_in[7] = (PIPERX4DATA[7] !== 1'bz) && PIPERX4DATA_delay[7]; // rv 0
  assign PIPERX4DATA_in[8] = (PIPERX4DATA[8] !== 1'bz) && PIPERX4DATA_delay[8]; // rv 0
  assign PIPERX4DATA_in[9] = (PIPERX4DATA[9] !== 1'bz) && PIPERX4DATA_delay[9]; // rv 0
  assign PIPERX4ELECIDLE_in = (PIPERX4ELECIDLE === 1'bz) || PIPERX4ELECIDLE_delay; // rv 1
  assign PIPERX4EQDONE_in = (PIPERX4EQDONE !== 1'bz) && PIPERX4EQDONE_delay; // rv 0
  assign PIPERX4EQLPADAPTDONE_in = (PIPERX4EQLPADAPTDONE !== 1'bz) && PIPERX4EQLPADAPTDONE_delay; // rv 0
  assign PIPERX4EQLPLFFSSEL_in = (PIPERX4EQLPLFFSSEL !== 1'bz) && PIPERX4EQLPLFFSSEL_delay; // rv 0
  assign PIPERX4EQLPNEWTXCOEFFORPRESET_in[0] = (PIPERX4EQLPNEWTXCOEFFORPRESET[0] !== 1'bz) && PIPERX4EQLPNEWTXCOEFFORPRESET_delay[0]; // rv 0
  assign PIPERX4EQLPNEWTXCOEFFORPRESET_in[10] = (PIPERX4EQLPNEWTXCOEFFORPRESET[10] !== 1'bz) && PIPERX4EQLPNEWTXCOEFFORPRESET_delay[10]; // rv 0
  assign PIPERX4EQLPNEWTXCOEFFORPRESET_in[11] = (PIPERX4EQLPNEWTXCOEFFORPRESET[11] !== 1'bz) && PIPERX4EQLPNEWTXCOEFFORPRESET_delay[11]; // rv 0
  assign PIPERX4EQLPNEWTXCOEFFORPRESET_in[12] = (PIPERX4EQLPNEWTXCOEFFORPRESET[12] !== 1'bz) && PIPERX4EQLPNEWTXCOEFFORPRESET_delay[12]; // rv 0
  assign PIPERX4EQLPNEWTXCOEFFORPRESET_in[13] = (PIPERX4EQLPNEWTXCOEFFORPRESET[13] !== 1'bz) && PIPERX4EQLPNEWTXCOEFFORPRESET_delay[13]; // rv 0
  assign PIPERX4EQLPNEWTXCOEFFORPRESET_in[14] = (PIPERX4EQLPNEWTXCOEFFORPRESET[14] !== 1'bz) && PIPERX4EQLPNEWTXCOEFFORPRESET_delay[14]; // rv 0
  assign PIPERX4EQLPNEWTXCOEFFORPRESET_in[15] = (PIPERX4EQLPNEWTXCOEFFORPRESET[15] !== 1'bz) && PIPERX4EQLPNEWTXCOEFFORPRESET_delay[15]; // rv 0
  assign PIPERX4EQLPNEWTXCOEFFORPRESET_in[16] = (PIPERX4EQLPNEWTXCOEFFORPRESET[16] !== 1'bz) && PIPERX4EQLPNEWTXCOEFFORPRESET_delay[16]; // rv 0
  assign PIPERX4EQLPNEWTXCOEFFORPRESET_in[17] = (PIPERX4EQLPNEWTXCOEFFORPRESET[17] !== 1'bz) && PIPERX4EQLPNEWTXCOEFFORPRESET_delay[17]; // rv 0
  assign PIPERX4EQLPNEWTXCOEFFORPRESET_in[1] = (PIPERX4EQLPNEWTXCOEFFORPRESET[1] !== 1'bz) && PIPERX4EQLPNEWTXCOEFFORPRESET_delay[1]; // rv 0
  assign PIPERX4EQLPNEWTXCOEFFORPRESET_in[2] = (PIPERX4EQLPNEWTXCOEFFORPRESET[2] !== 1'bz) && PIPERX4EQLPNEWTXCOEFFORPRESET_delay[2]; // rv 0
  assign PIPERX4EQLPNEWTXCOEFFORPRESET_in[3] = (PIPERX4EQLPNEWTXCOEFFORPRESET[3] !== 1'bz) && PIPERX4EQLPNEWTXCOEFFORPRESET_delay[3]; // rv 0
  assign PIPERX4EQLPNEWTXCOEFFORPRESET_in[4] = (PIPERX4EQLPNEWTXCOEFFORPRESET[4] !== 1'bz) && PIPERX4EQLPNEWTXCOEFFORPRESET_delay[4]; // rv 0
  assign PIPERX4EQLPNEWTXCOEFFORPRESET_in[5] = (PIPERX4EQLPNEWTXCOEFFORPRESET[5] !== 1'bz) && PIPERX4EQLPNEWTXCOEFFORPRESET_delay[5]; // rv 0
  assign PIPERX4EQLPNEWTXCOEFFORPRESET_in[6] = (PIPERX4EQLPNEWTXCOEFFORPRESET[6] !== 1'bz) && PIPERX4EQLPNEWTXCOEFFORPRESET_delay[6]; // rv 0
  assign PIPERX4EQLPNEWTXCOEFFORPRESET_in[7] = (PIPERX4EQLPNEWTXCOEFFORPRESET[7] !== 1'bz) && PIPERX4EQLPNEWTXCOEFFORPRESET_delay[7]; // rv 0
  assign PIPERX4EQLPNEWTXCOEFFORPRESET_in[8] = (PIPERX4EQLPNEWTXCOEFFORPRESET[8] !== 1'bz) && PIPERX4EQLPNEWTXCOEFFORPRESET_delay[8]; // rv 0
  assign PIPERX4EQLPNEWTXCOEFFORPRESET_in[9] = (PIPERX4EQLPNEWTXCOEFFORPRESET[9] !== 1'bz) && PIPERX4EQLPNEWTXCOEFFORPRESET_delay[9]; // rv 0
  assign PIPERX4PHYSTATUS_in = (PIPERX4PHYSTATUS === 1'bz) || PIPERX4PHYSTATUS_delay; // rv 1
  assign PIPERX4STARTBLOCK_in = (PIPERX4STARTBLOCK !== 1'bz) && PIPERX4STARTBLOCK_delay; // rv 0
  assign PIPERX4STATUS_in[0] = (PIPERX4STATUS[0] !== 1'bz) && PIPERX4STATUS_delay[0]; // rv 0
  assign PIPERX4STATUS_in[1] = (PIPERX4STATUS[1] !== 1'bz) && PIPERX4STATUS_delay[1]; // rv 0
  assign PIPERX4STATUS_in[2] = (PIPERX4STATUS[2] !== 1'bz) && PIPERX4STATUS_delay[2]; // rv 0
  assign PIPERX4SYNCHEADER_in[0] = (PIPERX4SYNCHEADER[0] !== 1'bz) && PIPERX4SYNCHEADER_delay[0]; // rv 0
  assign PIPERX4SYNCHEADER_in[1] = (PIPERX4SYNCHEADER[1] !== 1'bz) && PIPERX4SYNCHEADER_delay[1]; // rv 0
  assign PIPERX4VALID_in = (PIPERX4VALID !== 1'bz) && PIPERX4VALID_delay; // rv 0
  assign PIPERX5CHARISK_in[0] = (PIPERX5CHARISK[0] === 1'bz) || PIPERX5CHARISK_delay[0]; // rv 1
  assign PIPERX5CHARISK_in[1] = (PIPERX5CHARISK[1] === 1'bz) || PIPERX5CHARISK_delay[1]; // rv 1
  assign PIPERX5DATAVALID_in = (PIPERX5DATAVALID !== 1'bz) && PIPERX5DATAVALID_delay; // rv 0
  assign PIPERX5DATA_in[0] = (PIPERX5DATA[0] !== 1'bz) && PIPERX5DATA_delay[0]; // rv 0
  assign PIPERX5DATA_in[10] = (PIPERX5DATA[10] !== 1'bz) && PIPERX5DATA_delay[10]; // rv 0
  assign PIPERX5DATA_in[11] = (PIPERX5DATA[11] !== 1'bz) && PIPERX5DATA_delay[11]; // rv 0
  assign PIPERX5DATA_in[12] = (PIPERX5DATA[12] !== 1'bz) && PIPERX5DATA_delay[12]; // rv 0
  assign PIPERX5DATA_in[13] = (PIPERX5DATA[13] !== 1'bz) && PIPERX5DATA_delay[13]; // rv 0
  assign PIPERX5DATA_in[14] = (PIPERX5DATA[14] !== 1'bz) && PIPERX5DATA_delay[14]; // rv 0
  assign PIPERX5DATA_in[15] = (PIPERX5DATA[15] !== 1'bz) && PIPERX5DATA_delay[15]; // rv 0
  assign PIPERX5DATA_in[16] = (PIPERX5DATA[16] !== 1'bz) && PIPERX5DATA_delay[16]; // rv 0
  assign PIPERX5DATA_in[17] = (PIPERX5DATA[17] !== 1'bz) && PIPERX5DATA_delay[17]; // rv 0
  assign PIPERX5DATA_in[18] = (PIPERX5DATA[18] !== 1'bz) && PIPERX5DATA_delay[18]; // rv 0
  assign PIPERX5DATA_in[19] = (PIPERX5DATA[19] !== 1'bz) && PIPERX5DATA_delay[19]; // rv 0
  assign PIPERX5DATA_in[1] = (PIPERX5DATA[1] !== 1'bz) && PIPERX5DATA_delay[1]; // rv 0
  assign PIPERX5DATA_in[20] = (PIPERX5DATA[20] !== 1'bz) && PIPERX5DATA_delay[20]; // rv 0
  assign PIPERX5DATA_in[21] = (PIPERX5DATA[21] !== 1'bz) && PIPERX5DATA_delay[21]; // rv 0
  assign PIPERX5DATA_in[22] = (PIPERX5DATA[22] !== 1'bz) && PIPERX5DATA_delay[22]; // rv 0
  assign PIPERX5DATA_in[23] = (PIPERX5DATA[23] !== 1'bz) && PIPERX5DATA_delay[23]; // rv 0
  assign PIPERX5DATA_in[24] = (PIPERX5DATA[24] !== 1'bz) && PIPERX5DATA_delay[24]; // rv 0
  assign PIPERX5DATA_in[25] = (PIPERX5DATA[25] !== 1'bz) && PIPERX5DATA_delay[25]; // rv 0
  assign PIPERX5DATA_in[26] = (PIPERX5DATA[26] !== 1'bz) && PIPERX5DATA_delay[26]; // rv 0
  assign PIPERX5DATA_in[27] = (PIPERX5DATA[27] !== 1'bz) && PIPERX5DATA_delay[27]; // rv 0
  assign PIPERX5DATA_in[28] = (PIPERX5DATA[28] !== 1'bz) && PIPERX5DATA_delay[28]; // rv 0
  assign PIPERX5DATA_in[29] = (PIPERX5DATA[29] !== 1'bz) && PIPERX5DATA_delay[29]; // rv 0
  assign PIPERX5DATA_in[2] = (PIPERX5DATA[2] !== 1'bz) && PIPERX5DATA_delay[2]; // rv 0
  assign PIPERX5DATA_in[30] = (PIPERX5DATA[30] !== 1'bz) && PIPERX5DATA_delay[30]; // rv 0
  assign PIPERX5DATA_in[31] = (PIPERX5DATA[31] !== 1'bz) && PIPERX5DATA_delay[31]; // rv 0
  assign PIPERX5DATA_in[3] = (PIPERX5DATA[3] !== 1'bz) && PIPERX5DATA_delay[3]; // rv 0
  assign PIPERX5DATA_in[4] = (PIPERX5DATA[4] !== 1'bz) && PIPERX5DATA_delay[4]; // rv 0
  assign PIPERX5DATA_in[5] = (PIPERX5DATA[5] !== 1'bz) && PIPERX5DATA_delay[5]; // rv 0
  assign PIPERX5DATA_in[6] = (PIPERX5DATA[6] !== 1'bz) && PIPERX5DATA_delay[6]; // rv 0
  assign PIPERX5DATA_in[7] = (PIPERX5DATA[7] !== 1'bz) && PIPERX5DATA_delay[7]; // rv 0
  assign PIPERX5DATA_in[8] = (PIPERX5DATA[8] !== 1'bz) && PIPERX5DATA_delay[8]; // rv 0
  assign PIPERX5DATA_in[9] = (PIPERX5DATA[9] !== 1'bz) && PIPERX5DATA_delay[9]; // rv 0
  assign PIPERX5ELECIDLE_in = (PIPERX5ELECIDLE === 1'bz) || PIPERX5ELECIDLE_delay; // rv 1
  assign PIPERX5EQDONE_in = (PIPERX5EQDONE !== 1'bz) && PIPERX5EQDONE_delay; // rv 0
  assign PIPERX5EQLPADAPTDONE_in = (PIPERX5EQLPADAPTDONE !== 1'bz) && PIPERX5EQLPADAPTDONE_delay; // rv 0
  assign PIPERX5EQLPLFFSSEL_in = (PIPERX5EQLPLFFSSEL !== 1'bz) && PIPERX5EQLPLFFSSEL_delay; // rv 0
  assign PIPERX5EQLPNEWTXCOEFFORPRESET_in[0] = (PIPERX5EQLPNEWTXCOEFFORPRESET[0] !== 1'bz) && PIPERX5EQLPNEWTXCOEFFORPRESET_delay[0]; // rv 0
  assign PIPERX5EQLPNEWTXCOEFFORPRESET_in[10] = (PIPERX5EQLPNEWTXCOEFFORPRESET[10] !== 1'bz) && PIPERX5EQLPNEWTXCOEFFORPRESET_delay[10]; // rv 0
  assign PIPERX5EQLPNEWTXCOEFFORPRESET_in[11] = (PIPERX5EQLPNEWTXCOEFFORPRESET[11] !== 1'bz) && PIPERX5EQLPNEWTXCOEFFORPRESET_delay[11]; // rv 0
  assign PIPERX5EQLPNEWTXCOEFFORPRESET_in[12] = (PIPERX5EQLPNEWTXCOEFFORPRESET[12] !== 1'bz) && PIPERX5EQLPNEWTXCOEFFORPRESET_delay[12]; // rv 0
  assign PIPERX5EQLPNEWTXCOEFFORPRESET_in[13] = (PIPERX5EQLPNEWTXCOEFFORPRESET[13] !== 1'bz) && PIPERX5EQLPNEWTXCOEFFORPRESET_delay[13]; // rv 0
  assign PIPERX5EQLPNEWTXCOEFFORPRESET_in[14] = (PIPERX5EQLPNEWTXCOEFFORPRESET[14] !== 1'bz) && PIPERX5EQLPNEWTXCOEFFORPRESET_delay[14]; // rv 0
  assign PIPERX5EQLPNEWTXCOEFFORPRESET_in[15] = (PIPERX5EQLPNEWTXCOEFFORPRESET[15] !== 1'bz) && PIPERX5EQLPNEWTXCOEFFORPRESET_delay[15]; // rv 0
  assign PIPERX5EQLPNEWTXCOEFFORPRESET_in[16] = (PIPERX5EQLPNEWTXCOEFFORPRESET[16] !== 1'bz) && PIPERX5EQLPNEWTXCOEFFORPRESET_delay[16]; // rv 0
  assign PIPERX5EQLPNEWTXCOEFFORPRESET_in[17] = (PIPERX5EQLPNEWTXCOEFFORPRESET[17] !== 1'bz) && PIPERX5EQLPNEWTXCOEFFORPRESET_delay[17]; // rv 0
  assign PIPERX5EQLPNEWTXCOEFFORPRESET_in[1] = (PIPERX5EQLPNEWTXCOEFFORPRESET[1] !== 1'bz) && PIPERX5EQLPNEWTXCOEFFORPRESET_delay[1]; // rv 0
  assign PIPERX5EQLPNEWTXCOEFFORPRESET_in[2] = (PIPERX5EQLPNEWTXCOEFFORPRESET[2] !== 1'bz) && PIPERX5EQLPNEWTXCOEFFORPRESET_delay[2]; // rv 0
  assign PIPERX5EQLPNEWTXCOEFFORPRESET_in[3] = (PIPERX5EQLPNEWTXCOEFFORPRESET[3] !== 1'bz) && PIPERX5EQLPNEWTXCOEFFORPRESET_delay[3]; // rv 0
  assign PIPERX5EQLPNEWTXCOEFFORPRESET_in[4] = (PIPERX5EQLPNEWTXCOEFFORPRESET[4] !== 1'bz) && PIPERX5EQLPNEWTXCOEFFORPRESET_delay[4]; // rv 0
  assign PIPERX5EQLPNEWTXCOEFFORPRESET_in[5] = (PIPERX5EQLPNEWTXCOEFFORPRESET[5] !== 1'bz) && PIPERX5EQLPNEWTXCOEFFORPRESET_delay[5]; // rv 0
  assign PIPERX5EQLPNEWTXCOEFFORPRESET_in[6] = (PIPERX5EQLPNEWTXCOEFFORPRESET[6] !== 1'bz) && PIPERX5EQLPNEWTXCOEFFORPRESET_delay[6]; // rv 0
  assign PIPERX5EQLPNEWTXCOEFFORPRESET_in[7] = (PIPERX5EQLPNEWTXCOEFFORPRESET[7] !== 1'bz) && PIPERX5EQLPNEWTXCOEFFORPRESET_delay[7]; // rv 0
  assign PIPERX5EQLPNEWTXCOEFFORPRESET_in[8] = (PIPERX5EQLPNEWTXCOEFFORPRESET[8] !== 1'bz) && PIPERX5EQLPNEWTXCOEFFORPRESET_delay[8]; // rv 0
  assign PIPERX5EQLPNEWTXCOEFFORPRESET_in[9] = (PIPERX5EQLPNEWTXCOEFFORPRESET[9] !== 1'bz) && PIPERX5EQLPNEWTXCOEFFORPRESET_delay[9]; // rv 0
  assign PIPERX5PHYSTATUS_in = (PIPERX5PHYSTATUS === 1'bz) || PIPERX5PHYSTATUS_delay; // rv 1
  assign PIPERX5STARTBLOCK_in = (PIPERX5STARTBLOCK !== 1'bz) && PIPERX5STARTBLOCK_delay; // rv 0
  assign PIPERX5STATUS_in[0] = (PIPERX5STATUS[0] !== 1'bz) && PIPERX5STATUS_delay[0]; // rv 0
  assign PIPERX5STATUS_in[1] = (PIPERX5STATUS[1] !== 1'bz) && PIPERX5STATUS_delay[1]; // rv 0
  assign PIPERX5STATUS_in[2] = (PIPERX5STATUS[2] !== 1'bz) && PIPERX5STATUS_delay[2]; // rv 0
  assign PIPERX5SYNCHEADER_in[0] = (PIPERX5SYNCHEADER[0] !== 1'bz) && PIPERX5SYNCHEADER_delay[0]; // rv 0
  assign PIPERX5SYNCHEADER_in[1] = (PIPERX5SYNCHEADER[1] !== 1'bz) && PIPERX5SYNCHEADER_delay[1]; // rv 0
  assign PIPERX5VALID_in = (PIPERX5VALID !== 1'bz) && PIPERX5VALID_delay; // rv 0
  assign PIPERX6CHARISK_in[0] = (PIPERX6CHARISK[0] === 1'bz) || PIPERX6CHARISK_delay[0]; // rv 1
  assign PIPERX6CHARISK_in[1] = (PIPERX6CHARISK[1] === 1'bz) || PIPERX6CHARISK_delay[1]; // rv 1
  assign PIPERX6DATAVALID_in = (PIPERX6DATAVALID !== 1'bz) && PIPERX6DATAVALID_delay; // rv 0
  assign PIPERX6DATA_in[0] = (PIPERX6DATA[0] !== 1'bz) && PIPERX6DATA_delay[0]; // rv 0
  assign PIPERX6DATA_in[10] = (PIPERX6DATA[10] !== 1'bz) && PIPERX6DATA_delay[10]; // rv 0
  assign PIPERX6DATA_in[11] = (PIPERX6DATA[11] !== 1'bz) && PIPERX6DATA_delay[11]; // rv 0
  assign PIPERX6DATA_in[12] = (PIPERX6DATA[12] !== 1'bz) && PIPERX6DATA_delay[12]; // rv 0
  assign PIPERX6DATA_in[13] = (PIPERX6DATA[13] !== 1'bz) && PIPERX6DATA_delay[13]; // rv 0
  assign PIPERX6DATA_in[14] = (PIPERX6DATA[14] !== 1'bz) && PIPERX6DATA_delay[14]; // rv 0
  assign PIPERX6DATA_in[15] = (PIPERX6DATA[15] !== 1'bz) && PIPERX6DATA_delay[15]; // rv 0
  assign PIPERX6DATA_in[16] = (PIPERX6DATA[16] !== 1'bz) && PIPERX6DATA_delay[16]; // rv 0
  assign PIPERX6DATA_in[17] = (PIPERX6DATA[17] !== 1'bz) && PIPERX6DATA_delay[17]; // rv 0
  assign PIPERX6DATA_in[18] = (PIPERX6DATA[18] !== 1'bz) && PIPERX6DATA_delay[18]; // rv 0
  assign PIPERX6DATA_in[19] = (PIPERX6DATA[19] !== 1'bz) && PIPERX6DATA_delay[19]; // rv 0
  assign PIPERX6DATA_in[1] = (PIPERX6DATA[1] !== 1'bz) && PIPERX6DATA_delay[1]; // rv 0
  assign PIPERX6DATA_in[20] = (PIPERX6DATA[20] !== 1'bz) && PIPERX6DATA_delay[20]; // rv 0
  assign PIPERX6DATA_in[21] = (PIPERX6DATA[21] !== 1'bz) && PIPERX6DATA_delay[21]; // rv 0
  assign PIPERX6DATA_in[22] = (PIPERX6DATA[22] !== 1'bz) && PIPERX6DATA_delay[22]; // rv 0
  assign PIPERX6DATA_in[23] = (PIPERX6DATA[23] !== 1'bz) && PIPERX6DATA_delay[23]; // rv 0
  assign PIPERX6DATA_in[24] = (PIPERX6DATA[24] !== 1'bz) && PIPERX6DATA_delay[24]; // rv 0
  assign PIPERX6DATA_in[25] = (PIPERX6DATA[25] !== 1'bz) && PIPERX6DATA_delay[25]; // rv 0
  assign PIPERX6DATA_in[26] = (PIPERX6DATA[26] !== 1'bz) && PIPERX6DATA_delay[26]; // rv 0
  assign PIPERX6DATA_in[27] = (PIPERX6DATA[27] !== 1'bz) && PIPERX6DATA_delay[27]; // rv 0
  assign PIPERX6DATA_in[28] = (PIPERX6DATA[28] !== 1'bz) && PIPERX6DATA_delay[28]; // rv 0
  assign PIPERX6DATA_in[29] = (PIPERX6DATA[29] !== 1'bz) && PIPERX6DATA_delay[29]; // rv 0
  assign PIPERX6DATA_in[2] = (PIPERX6DATA[2] !== 1'bz) && PIPERX6DATA_delay[2]; // rv 0
  assign PIPERX6DATA_in[30] = (PIPERX6DATA[30] !== 1'bz) && PIPERX6DATA_delay[30]; // rv 0
  assign PIPERX6DATA_in[31] = (PIPERX6DATA[31] !== 1'bz) && PIPERX6DATA_delay[31]; // rv 0
  assign PIPERX6DATA_in[3] = (PIPERX6DATA[3] !== 1'bz) && PIPERX6DATA_delay[3]; // rv 0
  assign PIPERX6DATA_in[4] = (PIPERX6DATA[4] !== 1'bz) && PIPERX6DATA_delay[4]; // rv 0
  assign PIPERX6DATA_in[5] = (PIPERX6DATA[5] !== 1'bz) && PIPERX6DATA_delay[5]; // rv 0
  assign PIPERX6DATA_in[6] = (PIPERX6DATA[6] !== 1'bz) && PIPERX6DATA_delay[6]; // rv 0
  assign PIPERX6DATA_in[7] = (PIPERX6DATA[7] !== 1'bz) && PIPERX6DATA_delay[7]; // rv 0
  assign PIPERX6DATA_in[8] = (PIPERX6DATA[8] !== 1'bz) && PIPERX6DATA_delay[8]; // rv 0
  assign PIPERX6DATA_in[9] = (PIPERX6DATA[9] !== 1'bz) && PIPERX6DATA_delay[9]; // rv 0
  assign PIPERX6ELECIDLE_in = (PIPERX6ELECIDLE === 1'bz) || PIPERX6ELECIDLE_delay; // rv 1
  assign PIPERX6EQDONE_in = (PIPERX6EQDONE !== 1'bz) && PIPERX6EQDONE_delay; // rv 0
  assign PIPERX6EQLPADAPTDONE_in = (PIPERX6EQLPADAPTDONE !== 1'bz) && PIPERX6EQLPADAPTDONE_delay; // rv 0
  assign PIPERX6EQLPLFFSSEL_in = (PIPERX6EQLPLFFSSEL !== 1'bz) && PIPERX6EQLPLFFSSEL_delay; // rv 0
  assign PIPERX6EQLPNEWTXCOEFFORPRESET_in[0] = (PIPERX6EQLPNEWTXCOEFFORPRESET[0] !== 1'bz) && PIPERX6EQLPNEWTXCOEFFORPRESET_delay[0]; // rv 0
  assign PIPERX6EQLPNEWTXCOEFFORPRESET_in[10] = (PIPERX6EQLPNEWTXCOEFFORPRESET[10] !== 1'bz) && PIPERX6EQLPNEWTXCOEFFORPRESET_delay[10]; // rv 0
  assign PIPERX6EQLPNEWTXCOEFFORPRESET_in[11] = (PIPERX6EQLPNEWTXCOEFFORPRESET[11] !== 1'bz) && PIPERX6EQLPNEWTXCOEFFORPRESET_delay[11]; // rv 0
  assign PIPERX6EQLPNEWTXCOEFFORPRESET_in[12] = (PIPERX6EQLPNEWTXCOEFFORPRESET[12] !== 1'bz) && PIPERX6EQLPNEWTXCOEFFORPRESET_delay[12]; // rv 0
  assign PIPERX6EQLPNEWTXCOEFFORPRESET_in[13] = (PIPERX6EQLPNEWTXCOEFFORPRESET[13] !== 1'bz) && PIPERX6EQLPNEWTXCOEFFORPRESET_delay[13]; // rv 0
  assign PIPERX6EQLPNEWTXCOEFFORPRESET_in[14] = (PIPERX6EQLPNEWTXCOEFFORPRESET[14] !== 1'bz) && PIPERX6EQLPNEWTXCOEFFORPRESET_delay[14]; // rv 0
  assign PIPERX6EQLPNEWTXCOEFFORPRESET_in[15] = (PIPERX6EQLPNEWTXCOEFFORPRESET[15] !== 1'bz) && PIPERX6EQLPNEWTXCOEFFORPRESET_delay[15]; // rv 0
  assign PIPERX6EQLPNEWTXCOEFFORPRESET_in[16] = (PIPERX6EQLPNEWTXCOEFFORPRESET[16] !== 1'bz) && PIPERX6EQLPNEWTXCOEFFORPRESET_delay[16]; // rv 0
  assign PIPERX6EQLPNEWTXCOEFFORPRESET_in[17] = (PIPERX6EQLPNEWTXCOEFFORPRESET[17] !== 1'bz) && PIPERX6EQLPNEWTXCOEFFORPRESET_delay[17]; // rv 0
  assign PIPERX6EQLPNEWTXCOEFFORPRESET_in[1] = (PIPERX6EQLPNEWTXCOEFFORPRESET[1] !== 1'bz) && PIPERX6EQLPNEWTXCOEFFORPRESET_delay[1]; // rv 0
  assign PIPERX6EQLPNEWTXCOEFFORPRESET_in[2] = (PIPERX6EQLPNEWTXCOEFFORPRESET[2] !== 1'bz) && PIPERX6EQLPNEWTXCOEFFORPRESET_delay[2]; // rv 0
  assign PIPERX6EQLPNEWTXCOEFFORPRESET_in[3] = (PIPERX6EQLPNEWTXCOEFFORPRESET[3] !== 1'bz) && PIPERX6EQLPNEWTXCOEFFORPRESET_delay[3]; // rv 0
  assign PIPERX6EQLPNEWTXCOEFFORPRESET_in[4] = (PIPERX6EQLPNEWTXCOEFFORPRESET[4] !== 1'bz) && PIPERX6EQLPNEWTXCOEFFORPRESET_delay[4]; // rv 0
  assign PIPERX6EQLPNEWTXCOEFFORPRESET_in[5] = (PIPERX6EQLPNEWTXCOEFFORPRESET[5] !== 1'bz) && PIPERX6EQLPNEWTXCOEFFORPRESET_delay[5]; // rv 0
  assign PIPERX6EQLPNEWTXCOEFFORPRESET_in[6] = (PIPERX6EQLPNEWTXCOEFFORPRESET[6] !== 1'bz) && PIPERX6EQLPNEWTXCOEFFORPRESET_delay[6]; // rv 0
  assign PIPERX6EQLPNEWTXCOEFFORPRESET_in[7] = (PIPERX6EQLPNEWTXCOEFFORPRESET[7] !== 1'bz) && PIPERX6EQLPNEWTXCOEFFORPRESET_delay[7]; // rv 0
  assign PIPERX6EQLPNEWTXCOEFFORPRESET_in[8] = (PIPERX6EQLPNEWTXCOEFFORPRESET[8] !== 1'bz) && PIPERX6EQLPNEWTXCOEFFORPRESET_delay[8]; // rv 0
  assign PIPERX6EQLPNEWTXCOEFFORPRESET_in[9] = (PIPERX6EQLPNEWTXCOEFFORPRESET[9] !== 1'bz) && PIPERX6EQLPNEWTXCOEFFORPRESET_delay[9]; // rv 0
  assign PIPERX6PHYSTATUS_in = (PIPERX6PHYSTATUS === 1'bz) || PIPERX6PHYSTATUS_delay; // rv 1
  assign PIPERX6STARTBLOCK_in = (PIPERX6STARTBLOCK !== 1'bz) && PIPERX6STARTBLOCK_delay; // rv 0
  assign PIPERX6STATUS_in[0] = (PIPERX6STATUS[0] !== 1'bz) && PIPERX6STATUS_delay[0]; // rv 0
  assign PIPERX6STATUS_in[1] = (PIPERX6STATUS[1] !== 1'bz) && PIPERX6STATUS_delay[1]; // rv 0
  assign PIPERX6STATUS_in[2] = (PIPERX6STATUS[2] !== 1'bz) && PIPERX6STATUS_delay[2]; // rv 0
  assign PIPERX6SYNCHEADER_in[0] = (PIPERX6SYNCHEADER[0] !== 1'bz) && PIPERX6SYNCHEADER_delay[0]; // rv 0
  assign PIPERX6SYNCHEADER_in[1] = (PIPERX6SYNCHEADER[1] !== 1'bz) && PIPERX6SYNCHEADER_delay[1]; // rv 0
  assign PIPERX6VALID_in = (PIPERX6VALID !== 1'bz) && PIPERX6VALID_delay; // rv 0
  assign PIPERX7CHARISK_in[0] = (PIPERX7CHARISK[0] === 1'bz) || PIPERX7CHARISK_delay[0]; // rv 1
  assign PIPERX7CHARISK_in[1] = (PIPERX7CHARISK[1] === 1'bz) || PIPERX7CHARISK_delay[1]; // rv 1
  assign PIPERX7DATAVALID_in = (PIPERX7DATAVALID !== 1'bz) && PIPERX7DATAVALID_delay; // rv 0
  assign PIPERX7DATA_in[0] = (PIPERX7DATA[0] !== 1'bz) && PIPERX7DATA_delay[0]; // rv 0
  assign PIPERX7DATA_in[10] = (PIPERX7DATA[10] !== 1'bz) && PIPERX7DATA_delay[10]; // rv 0
  assign PIPERX7DATA_in[11] = (PIPERX7DATA[11] !== 1'bz) && PIPERX7DATA_delay[11]; // rv 0
  assign PIPERX7DATA_in[12] = (PIPERX7DATA[12] !== 1'bz) && PIPERX7DATA_delay[12]; // rv 0
  assign PIPERX7DATA_in[13] = (PIPERX7DATA[13] !== 1'bz) && PIPERX7DATA_delay[13]; // rv 0
  assign PIPERX7DATA_in[14] = (PIPERX7DATA[14] !== 1'bz) && PIPERX7DATA_delay[14]; // rv 0
  assign PIPERX7DATA_in[15] = (PIPERX7DATA[15] !== 1'bz) && PIPERX7DATA_delay[15]; // rv 0
  assign PIPERX7DATA_in[16] = (PIPERX7DATA[16] !== 1'bz) && PIPERX7DATA_delay[16]; // rv 0
  assign PIPERX7DATA_in[17] = (PIPERX7DATA[17] !== 1'bz) && PIPERX7DATA_delay[17]; // rv 0
  assign PIPERX7DATA_in[18] = (PIPERX7DATA[18] !== 1'bz) && PIPERX7DATA_delay[18]; // rv 0
  assign PIPERX7DATA_in[19] = (PIPERX7DATA[19] !== 1'bz) && PIPERX7DATA_delay[19]; // rv 0
  assign PIPERX7DATA_in[1] = (PIPERX7DATA[1] !== 1'bz) && PIPERX7DATA_delay[1]; // rv 0
  assign PIPERX7DATA_in[20] = (PIPERX7DATA[20] !== 1'bz) && PIPERX7DATA_delay[20]; // rv 0
  assign PIPERX7DATA_in[21] = (PIPERX7DATA[21] !== 1'bz) && PIPERX7DATA_delay[21]; // rv 0
  assign PIPERX7DATA_in[22] = (PIPERX7DATA[22] !== 1'bz) && PIPERX7DATA_delay[22]; // rv 0
  assign PIPERX7DATA_in[23] = (PIPERX7DATA[23] !== 1'bz) && PIPERX7DATA_delay[23]; // rv 0
  assign PIPERX7DATA_in[24] = (PIPERX7DATA[24] !== 1'bz) && PIPERX7DATA_delay[24]; // rv 0
  assign PIPERX7DATA_in[25] = (PIPERX7DATA[25] !== 1'bz) && PIPERX7DATA_delay[25]; // rv 0
  assign PIPERX7DATA_in[26] = (PIPERX7DATA[26] !== 1'bz) && PIPERX7DATA_delay[26]; // rv 0
  assign PIPERX7DATA_in[27] = (PIPERX7DATA[27] !== 1'bz) && PIPERX7DATA_delay[27]; // rv 0
  assign PIPERX7DATA_in[28] = (PIPERX7DATA[28] !== 1'bz) && PIPERX7DATA_delay[28]; // rv 0
  assign PIPERX7DATA_in[29] = (PIPERX7DATA[29] !== 1'bz) && PIPERX7DATA_delay[29]; // rv 0
  assign PIPERX7DATA_in[2] = (PIPERX7DATA[2] !== 1'bz) && PIPERX7DATA_delay[2]; // rv 0
  assign PIPERX7DATA_in[30] = (PIPERX7DATA[30] !== 1'bz) && PIPERX7DATA_delay[30]; // rv 0
  assign PIPERX7DATA_in[31] = (PIPERX7DATA[31] !== 1'bz) && PIPERX7DATA_delay[31]; // rv 0
  assign PIPERX7DATA_in[3] = (PIPERX7DATA[3] !== 1'bz) && PIPERX7DATA_delay[3]; // rv 0
  assign PIPERX7DATA_in[4] = (PIPERX7DATA[4] !== 1'bz) && PIPERX7DATA_delay[4]; // rv 0
  assign PIPERX7DATA_in[5] = (PIPERX7DATA[5] !== 1'bz) && PIPERX7DATA_delay[5]; // rv 0
  assign PIPERX7DATA_in[6] = (PIPERX7DATA[6] !== 1'bz) && PIPERX7DATA_delay[6]; // rv 0
  assign PIPERX7DATA_in[7] = (PIPERX7DATA[7] !== 1'bz) && PIPERX7DATA_delay[7]; // rv 0
  assign PIPERX7DATA_in[8] = (PIPERX7DATA[8] !== 1'bz) && PIPERX7DATA_delay[8]; // rv 0
  assign PIPERX7DATA_in[9] = (PIPERX7DATA[9] !== 1'bz) && PIPERX7DATA_delay[9]; // rv 0
  assign PIPERX7ELECIDLE_in = (PIPERX7ELECIDLE === 1'bz) || PIPERX7ELECIDLE_delay; // rv 1
  assign PIPERX7EQDONE_in = (PIPERX7EQDONE !== 1'bz) && PIPERX7EQDONE_delay; // rv 0
  assign PIPERX7EQLPADAPTDONE_in = (PIPERX7EQLPADAPTDONE !== 1'bz) && PIPERX7EQLPADAPTDONE_delay; // rv 0
  assign PIPERX7EQLPLFFSSEL_in = (PIPERX7EQLPLFFSSEL !== 1'bz) && PIPERX7EQLPLFFSSEL_delay; // rv 0
  assign PIPERX7EQLPNEWTXCOEFFORPRESET_in[0] = (PIPERX7EQLPNEWTXCOEFFORPRESET[0] !== 1'bz) && PIPERX7EQLPNEWTXCOEFFORPRESET_delay[0]; // rv 0
  assign PIPERX7EQLPNEWTXCOEFFORPRESET_in[10] = (PIPERX7EQLPNEWTXCOEFFORPRESET[10] !== 1'bz) && PIPERX7EQLPNEWTXCOEFFORPRESET_delay[10]; // rv 0
  assign PIPERX7EQLPNEWTXCOEFFORPRESET_in[11] = (PIPERX7EQLPNEWTXCOEFFORPRESET[11] !== 1'bz) && PIPERX7EQLPNEWTXCOEFFORPRESET_delay[11]; // rv 0
  assign PIPERX7EQLPNEWTXCOEFFORPRESET_in[12] = (PIPERX7EQLPNEWTXCOEFFORPRESET[12] !== 1'bz) && PIPERX7EQLPNEWTXCOEFFORPRESET_delay[12]; // rv 0
  assign PIPERX7EQLPNEWTXCOEFFORPRESET_in[13] = (PIPERX7EQLPNEWTXCOEFFORPRESET[13] !== 1'bz) && PIPERX7EQLPNEWTXCOEFFORPRESET_delay[13]; // rv 0
  assign PIPERX7EQLPNEWTXCOEFFORPRESET_in[14] = (PIPERX7EQLPNEWTXCOEFFORPRESET[14] !== 1'bz) && PIPERX7EQLPNEWTXCOEFFORPRESET_delay[14]; // rv 0
  assign PIPERX7EQLPNEWTXCOEFFORPRESET_in[15] = (PIPERX7EQLPNEWTXCOEFFORPRESET[15] !== 1'bz) && PIPERX7EQLPNEWTXCOEFFORPRESET_delay[15]; // rv 0
  assign PIPERX7EQLPNEWTXCOEFFORPRESET_in[16] = (PIPERX7EQLPNEWTXCOEFFORPRESET[16] !== 1'bz) && PIPERX7EQLPNEWTXCOEFFORPRESET_delay[16]; // rv 0
  assign PIPERX7EQLPNEWTXCOEFFORPRESET_in[17] = (PIPERX7EQLPNEWTXCOEFFORPRESET[17] !== 1'bz) && PIPERX7EQLPNEWTXCOEFFORPRESET_delay[17]; // rv 0
  assign PIPERX7EQLPNEWTXCOEFFORPRESET_in[1] = (PIPERX7EQLPNEWTXCOEFFORPRESET[1] !== 1'bz) && PIPERX7EQLPNEWTXCOEFFORPRESET_delay[1]; // rv 0
  assign PIPERX7EQLPNEWTXCOEFFORPRESET_in[2] = (PIPERX7EQLPNEWTXCOEFFORPRESET[2] !== 1'bz) && PIPERX7EQLPNEWTXCOEFFORPRESET_delay[2]; // rv 0
  assign PIPERX7EQLPNEWTXCOEFFORPRESET_in[3] = (PIPERX7EQLPNEWTXCOEFFORPRESET[3] !== 1'bz) && PIPERX7EQLPNEWTXCOEFFORPRESET_delay[3]; // rv 0
  assign PIPERX7EQLPNEWTXCOEFFORPRESET_in[4] = (PIPERX7EQLPNEWTXCOEFFORPRESET[4] !== 1'bz) && PIPERX7EQLPNEWTXCOEFFORPRESET_delay[4]; // rv 0
  assign PIPERX7EQLPNEWTXCOEFFORPRESET_in[5] = (PIPERX7EQLPNEWTXCOEFFORPRESET[5] !== 1'bz) && PIPERX7EQLPNEWTXCOEFFORPRESET_delay[5]; // rv 0
  assign PIPERX7EQLPNEWTXCOEFFORPRESET_in[6] = (PIPERX7EQLPNEWTXCOEFFORPRESET[6] !== 1'bz) && PIPERX7EQLPNEWTXCOEFFORPRESET_delay[6]; // rv 0
  assign PIPERX7EQLPNEWTXCOEFFORPRESET_in[7] = (PIPERX7EQLPNEWTXCOEFFORPRESET[7] !== 1'bz) && PIPERX7EQLPNEWTXCOEFFORPRESET_delay[7]; // rv 0
  assign PIPERX7EQLPNEWTXCOEFFORPRESET_in[8] = (PIPERX7EQLPNEWTXCOEFFORPRESET[8] !== 1'bz) && PIPERX7EQLPNEWTXCOEFFORPRESET_delay[8]; // rv 0
  assign PIPERX7EQLPNEWTXCOEFFORPRESET_in[9] = (PIPERX7EQLPNEWTXCOEFFORPRESET[9] !== 1'bz) && PIPERX7EQLPNEWTXCOEFFORPRESET_delay[9]; // rv 0
  assign PIPERX7PHYSTATUS_in = (PIPERX7PHYSTATUS === 1'bz) || PIPERX7PHYSTATUS_delay; // rv 1
  assign PIPERX7STARTBLOCK_in = (PIPERX7STARTBLOCK !== 1'bz) && PIPERX7STARTBLOCK_delay; // rv 0
  assign PIPERX7STATUS_in[0] = (PIPERX7STATUS[0] !== 1'bz) && PIPERX7STATUS_delay[0]; // rv 0
  assign PIPERX7STATUS_in[1] = (PIPERX7STATUS[1] !== 1'bz) && PIPERX7STATUS_delay[1]; // rv 0
  assign PIPERX7STATUS_in[2] = (PIPERX7STATUS[2] !== 1'bz) && PIPERX7STATUS_delay[2]; // rv 0
  assign PIPERX7SYNCHEADER_in[0] = (PIPERX7SYNCHEADER[0] !== 1'bz) && PIPERX7SYNCHEADER_delay[0]; // rv 0
  assign PIPERX7SYNCHEADER_in[1] = (PIPERX7SYNCHEADER[1] !== 1'bz) && PIPERX7SYNCHEADER_delay[1]; // rv 0
  assign PIPERX7VALID_in = (PIPERX7VALID !== 1'bz) && PIPERX7VALID_delay; // rv 0
  assign PIPETX0EQCOEFF_in[0] = (PIPETX0EQCOEFF[0] !== 1'bz) && PIPETX0EQCOEFF_delay[0]; // rv 0
  assign PIPETX0EQCOEFF_in[10] = (PIPETX0EQCOEFF[10] !== 1'bz) && PIPETX0EQCOEFF_delay[10]; // rv 0
  assign PIPETX0EQCOEFF_in[11] = (PIPETX0EQCOEFF[11] !== 1'bz) && PIPETX0EQCOEFF_delay[11]; // rv 0
  assign PIPETX0EQCOEFF_in[12] = (PIPETX0EQCOEFF[12] !== 1'bz) && PIPETX0EQCOEFF_delay[12]; // rv 0
  assign PIPETX0EQCOEFF_in[13] = (PIPETX0EQCOEFF[13] !== 1'bz) && PIPETX0EQCOEFF_delay[13]; // rv 0
  assign PIPETX0EQCOEFF_in[14] = (PIPETX0EQCOEFF[14] !== 1'bz) && PIPETX0EQCOEFF_delay[14]; // rv 0
  assign PIPETX0EQCOEFF_in[15] = (PIPETX0EQCOEFF[15] !== 1'bz) && PIPETX0EQCOEFF_delay[15]; // rv 0
  assign PIPETX0EQCOEFF_in[16] = (PIPETX0EQCOEFF[16] !== 1'bz) && PIPETX0EQCOEFF_delay[16]; // rv 0
  assign PIPETX0EQCOEFF_in[17] = (PIPETX0EQCOEFF[17] !== 1'bz) && PIPETX0EQCOEFF_delay[17]; // rv 0
  assign PIPETX0EQCOEFF_in[1] = (PIPETX0EQCOEFF[1] !== 1'bz) && PIPETX0EQCOEFF_delay[1]; // rv 0
  assign PIPETX0EQCOEFF_in[2] = (PIPETX0EQCOEFF[2] !== 1'bz) && PIPETX0EQCOEFF_delay[2]; // rv 0
  assign PIPETX0EQCOEFF_in[3] = (PIPETX0EQCOEFF[3] !== 1'bz) && PIPETX0EQCOEFF_delay[3]; // rv 0
  assign PIPETX0EQCOEFF_in[4] = (PIPETX0EQCOEFF[4] !== 1'bz) && PIPETX0EQCOEFF_delay[4]; // rv 0
  assign PIPETX0EQCOEFF_in[5] = (PIPETX0EQCOEFF[5] !== 1'bz) && PIPETX0EQCOEFF_delay[5]; // rv 0
  assign PIPETX0EQCOEFF_in[6] = (PIPETX0EQCOEFF[6] !== 1'bz) && PIPETX0EQCOEFF_delay[6]; // rv 0
  assign PIPETX0EQCOEFF_in[7] = (PIPETX0EQCOEFF[7] !== 1'bz) && PIPETX0EQCOEFF_delay[7]; // rv 0
  assign PIPETX0EQCOEFF_in[8] = (PIPETX0EQCOEFF[8] !== 1'bz) && PIPETX0EQCOEFF_delay[8]; // rv 0
  assign PIPETX0EQCOEFF_in[9] = (PIPETX0EQCOEFF[9] !== 1'bz) && PIPETX0EQCOEFF_delay[9]; // rv 0
  assign PIPETX0EQDONE_in = (PIPETX0EQDONE !== 1'bz) && PIPETX0EQDONE_delay; // rv 0
  assign PIPETX1EQCOEFF_in[0] = (PIPETX1EQCOEFF[0] !== 1'bz) && PIPETX1EQCOEFF_delay[0]; // rv 0
  assign PIPETX1EQCOEFF_in[10] = (PIPETX1EQCOEFF[10] !== 1'bz) && PIPETX1EQCOEFF_delay[10]; // rv 0
  assign PIPETX1EQCOEFF_in[11] = (PIPETX1EQCOEFF[11] !== 1'bz) && PIPETX1EQCOEFF_delay[11]; // rv 0
  assign PIPETX1EQCOEFF_in[12] = (PIPETX1EQCOEFF[12] !== 1'bz) && PIPETX1EQCOEFF_delay[12]; // rv 0
  assign PIPETX1EQCOEFF_in[13] = (PIPETX1EQCOEFF[13] !== 1'bz) && PIPETX1EQCOEFF_delay[13]; // rv 0
  assign PIPETX1EQCOEFF_in[14] = (PIPETX1EQCOEFF[14] !== 1'bz) && PIPETX1EQCOEFF_delay[14]; // rv 0
  assign PIPETX1EQCOEFF_in[15] = (PIPETX1EQCOEFF[15] !== 1'bz) && PIPETX1EQCOEFF_delay[15]; // rv 0
  assign PIPETX1EQCOEFF_in[16] = (PIPETX1EQCOEFF[16] !== 1'bz) && PIPETX1EQCOEFF_delay[16]; // rv 0
  assign PIPETX1EQCOEFF_in[17] = (PIPETX1EQCOEFF[17] !== 1'bz) && PIPETX1EQCOEFF_delay[17]; // rv 0
  assign PIPETX1EQCOEFF_in[1] = (PIPETX1EQCOEFF[1] !== 1'bz) && PIPETX1EQCOEFF_delay[1]; // rv 0
  assign PIPETX1EQCOEFF_in[2] = (PIPETX1EQCOEFF[2] !== 1'bz) && PIPETX1EQCOEFF_delay[2]; // rv 0
  assign PIPETX1EQCOEFF_in[3] = (PIPETX1EQCOEFF[3] !== 1'bz) && PIPETX1EQCOEFF_delay[3]; // rv 0
  assign PIPETX1EQCOEFF_in[4] = (PIPETX1EQCOEFF[4] !== 1'bz) && PIPETX1EQCOEFF_delay[4]; // rv 0
  assign PIPETX1EQCOEFF_in[5] = (PIPETX1EQCOEFF[5] !== 1'bz) && PIPETX1EQCOEFF_delay[5]; // rv 0
  assign PIPETX1EQCOEFF_in[6] = (PIPETX1EQCOEFF[6] !== 1'bz) && PIPETX1EQCOEFF_delay[6]; // rv 0
  assign PIPETX1EQCOEFF_in[7] = (PIPETX1EQCOEFF[7] !== 1'bz) && PIPETX1EQCOEFF_delay[7]; // rv 0
  assign PIPETX1EQCOEFF_in[8] = (PIPETX1EQCOEFF[8] !== 1'bz) && PIPETX1EQCOEFF_delay[8]; // rv 0
  assign PIPETX1EQCOEFF_in[9] = (PIPETX1EQCOEFF[9] !== 1'bz) && PIPETX1EQCOEFF_delay[9]; // rv 0
  assign PIPETX1EQDONE_in = (PIPETX1EQDONE !== 1'bz) && PIPETX1EQDONE_delay; // rv 0
  assign PIPETX2EQCOEFF_in[0] = (PIPETX2EQCOEFF[0] !== 1'bz) && PIPETX2EQCOEFF_delay[0]; // rv 0
  assign PIPETX2EQCOEFF_in[10] = (PIPETX2EQCOEFF[10] !== 1'bz) && PIPETX2EQCOEFF_delay[10]; // rv 0
  assign PIPETX2EQCOEFF_in[11] = (PIPETX2EQCOEFF[11] !== 1'bz) && PIPETX2EQCOEFF_delay[11]; // rv 0
  assign PIPETX2EQCOEFF_in[12] = (PIPETX2EQCOEFF[12] !== 1'bz) && PIPETX2EQCOEFF_delay[12]; // rv 0
  assign PIPETX2EQCOEFF_in[13] = (PIPETX2EQCOEFF[13] !== 1'bz) && PIPETX2EQCOEFF_delay[13]; // rv 0
  assign PIPETX2EQCOEFF_in[14] = (PIPETX2EQCOEFF[14] !== 1'bz) && PIPETX2EQCOEFF_delay[14]; // rv 0
  assign PIPETX2EQCOEFF_in[15] = (PIPETX2EQCOEFF[15] !== 1'bz) && PIPETX2EQCOEFF_delay[15]; // rv 0
  assign PIPETX2EQCOEFF_in[16] = (PIPETX2EQCOEFF[16] !== 1'bz) && PIPETX2EQCOEFF_delay[16]; // rv 0
  assign PIPETX2EQCOEFF_in[17] = (PIPETX2EQCOEFF[17] !== 1'bz) && PIPETX2EQCOEFF_delay[17]; // rv 0
  assign PIPETX2EQCOEFF_in[1] = (PIPETX2EQCOEFF[1] !== 1'bz) && PIPETX2EQCOEFF_delay[1]; // rv 0
  assign PIPETX2EQCOEFF_in[2] = (PIPETX2EQCOEFF[2] !== 1'bz) && PIPETX2EQCOEFF_delay[2]; // rv 0
  assign PIPETX2EQCOEFF_in[3] = (PIPETX2EQCOEFF[3] !== 1'bz) && PIPETX2EQCOEFF_delay[3]; // rv 0
  assign PIPETX2EQCOEFF_in[4] = (PIPETX2EQCOEFF[4] !== 1'bz) && PIPETX2EQCOEFF_delay[4]; // rv 0
  assign PIPETX2EQCOEFF_in[5] = (PIPETX2EQCOEFF[5] !== 1'bz) && PIPETX2EQCOEFF_delay[5]; // rv 0
  assign PIPETX2EQCOEFF_in[6] = (PIPETX2EQCOEFF[6] !== 1'bz) && PIPETX2EQCOEFF_delay[6]; // rv 0
  assign PIPETX2EQCOEFF_in[7] = (PIPETX2EQCOEFF[7] !== 1'bz) && PIPETX2EQCOEFF_delay[7]; // rv 0
  assign PIPETX2EQCOEFF_in[8] = (PIPETX2EQCOEFF[8] !== 1'bz) && PIPETX2EQCOEFF_delay[8]; // rv 0
  assign PIPETX2EQCOEFF_in[9] = (PIPETX2EQCOEFF[9] !== 1'bz) && PIPETX2EQCOEFF_delay[9]; // rv 0
  assign PIPETX2EQDONE_in = (PIPETX2EQDONE !== 1'bz) && PIPETX2EQDONE_delay; // rv 0
  assign PIPETX3EQCOEFF_in[0] = (PIPETX3EQCOEFF[0] !== 1'bz) && PIPETX3EQCOEFF_delay[0]; // rv 0
  assign PIPETX3EQCOEFF_in[10] = (PIPETX3EQCOEFF[10] !== 1'bz) && PIPETX3EQCOEFF_delay[10]; // rv 0
  assign PIPETX3EQCOEFF_in[11] = (PIPETX3EQCOEFF[11] !== 1'bz) && PIPETX3EQCOEFF_delay[11]; // rv 0
  assign PIPETX3EQCOEFF_in[12] = (PIPETX3EQCOEFF[12] !== 1'bz) && PIPETX3EQCOEFF_delay[12]; // rv 0
  assign PIPETX3EQCOEFF_in[13] = (PIPETX3EQCOEFF[13] !== 1'bz) && PIPETX3EQCOEFF_delay[13]; // rv 0
  assign PIPETX3EQCOEFF_in[14] = (PIPETX3EQCOEFF[14] !== 1'bz) && PIPETX3EQCOEFF_delay[14]; // rv 0
  assign PIPETX3EQCOEFF_in[15] = (PIPETX3EQCOEFF[15] !== 1'bz) && PIPETX3EQCOEFF_delay[15]; // rv 0
  assign PIPETX3EQCOEFF_in[16] = (PIPETX3EQCOEFF[16] !== 1'bz) && PIPETX3EQCOEFF_delay[16]; // rv 0
  assign PIPETX3EQCOEFF_in[17] = (PIPETX3EQCOEFF[17] !== 1'bz) && PIPETX3EQCOEFF_delay[17]; // rv 0
  assign PIPETX3EQCOEFF_in[1] = (PIPETX3EQCOEFF[1] !== 1'bz) && PIPETX3EQCOEFF_delay[1]; // rv 0
  assign PIPETX3EQCOEFF_in[2] = (PIPETX3EQCOEFF[2] !== 1'bz) && PIPETX3EQCOEFF_delay[2]; // rv 0
  assign PIPETX3EQCOEFF_in[3] = (PIPETX3EQCOEFF[3] !== 1'bz) && PIPETX3EQCOEFF_delay[3]; // rv 0
  assign PIPETX3EQCOEFF_in[4] = (PIPETX3EQCOEFF[4] !== 1'bz) && PIPETX3EQCOEFF_delay[4]; // rv 0
  assign PIPETX3EQCOEFF_in[5] = (PIPETX3EQCOEFF[5] !== 1'bz) && PIPETX3EQCOEFF_delay[5]; // rv 0
  assign PIPETX3EQCOEFF_in[6] = (PIPETX3EQCOEFF[6] !== 1'bz) && PIPETX3EQCOEFF_delay[6]; // rv 0
  assign PIPETX3EQCOEFF_in[7] = (PIPETX3EQCOEFF[7] !== 1'bz) && PIPETX3EQCOEFF_delay[7]; // rv 0
  assign PIPETX3EQCOEFF_in[8] = (PIPETX3EQCOEFF[8] !== 1'bz) && PIPETX3EQCOEFF_delay[8]; // rv 0
  assign PIPETX3EQCOEFF_in[9] = (PIPETX3EQCOEFF[9] !== 1'bz) && PIPETX3EQCOEFF_delay[9]; // rv 0
  assign PIPETX3EQDONE_in = (PIPETX3EQDONE !== 1'bz) && PIPETX3EQDONE_delay; // rv 0
  assign PIPETX4EQCOEFF_in[0] = (PIPETX4EQCOEFF[0] !== 1'bz) && PIPETX4EQCOEFF_delay[0]; // rv 0
  assign PIPETX4EQCOEFF_in[10] = (PIPETX4EQCOEFF[10] !== 1'bz) && PIPETX4EQCOEFF_delay[10]; // rv 0
  assign PIPETX4EQCOEFF_in[11] = (PIPETX4EQCOEFF[11] !== 1'bz) && PIPETX4EQCOEFF_delay[11]; // rv 0
  assign PIPETX4EQCOEFF_in[12] = (PIPETX4EQCOEFF[12] !== 1'bz) && PIPETX4EQCOEFF_delay[12]; // rv 0
  assign PIPETX4EQCOEFF_in[13] = (PIPETX4EQCOEFF[13] !== 1'bz) && PIPETX4EQCOEFF_delay[13]; // rv 0
  assign PIPETX4EQCOEFF_in[14] = (PIPETX4EQCOEFF[14] !== 1'bz) && PIPETX4EQCOEFF_delay[14]; // rv 0
  assign PIPETX4EQCOEFF_in[15] = (PIPETX4EQCOEFF[15] !== 1'bz) && PIPETX4EQCOEFF_delay[15]; // rv 0
  assign PIPETX4EQCOEFF_in[16] = (PIPETX4EQCOEFF[16] !== 1'bz) && PIPETX4EQCOEFF_delay[16]; // rv 0
  assign PIPETX4EQCOEFF_in[17] = (PIPETX4EQCOEFF[17] !== 1'bz) && PIPETX4EQCOEFF_delay[17]; // rv 0
  assign PIPETX4EQCOEFF_in[1] = (PIPETX4EQCOEFF[1] !== 1'bz) && PIPETX4EQCOEFF_delay[1]; // rv 0
  assign PIPETX4EQCOEFF_in[2] = (PIPETX4EQCOEFF[2] !== 1'bz) && PIPETX4EQCOEFF_delay[2]; // rv 0
  assign PIPETX4EQCOEFF_in[3] = (PIPETX4EQCOEFF[3] !== 1'bz) && PIPETX4EQCOEFF_delay[3]; // rv 0
  assign PIPETX4EQCOEFF_in[4] = (PIPETX4EQCOEFF[4] !== 1'bz) && PIPETX4EQCOEFF_delay[4]; // rv 0
  assign PIPETX4EQCOEFF_in[5] = (PIPETX4EQCOEFF[5] !== 1'bz) && PIPETX4EQCOEFF_delay[5]; // rv 0
  assign PIPETX4EQCOEFF_in[6] = (PIPETX4EQCOEFF[6] !== 1'bz) && PIPETX4EQCOEFF_delay[6]; // rv 0
  assign PIPETX4EQCOEFF_in[7] = (PIPETX4EQCOEFF[7] !== 1'bz) && PIPETX4EQCOEFF_delay[7]; // rv 0
  assign PIPETX4EQCOEFF_in[8] = (PIPETX4EQCOEFF[8] !== 1'bz) && PIPETX4EQCOEFF_delay[8]; // rv 0
  assign PIPETX4EQCOEFF_in[9] = (PIPETX4EQCOEFF[9] !== 1'bz) && PIPETX4EQCOEFF_delay[9]; // rv 0
  assign PIPETX4EQDONE_in = (PIPETX4EQDONE !== 1'bz) && PIPETX4EQDONE_delay; // rv 0
  assign PIPETX5EQCOEFF_in[0] = (PIPETX5EQCOEFF[0] !== 1'bz) && PIPETX5EQCOEFF_delay[0]; // rv 0
  assign PIPETX5EQCOEFF_in[10] = (PIPETX5EQCOEFF[10] !== 1'bz) && PIPETX5EQCOEFF_delay[10]; // rv 0
  assign PIPETX5EQCOEFF_in[11] = (PIPETX5EQCOEFF[11] !== 1'bz) && PIPETX5EQCOEFF_delay[11]; // rv 0
  assign PIPETX5EQCOEFF_in[12] = (PIPETX5EQCOEFF[12] !== 1'bz) && PIPETX5EQCOEFF_delay[12]; // rv 0
  assign PIPETX5EQCOEFF_in[13] = (PIPETX5EQCOEFF[13] !== 1'bz) && PIPETX5EQCOEFF_delay[13]; // rv 0
  assign PIPETX5EQCOEFF_in[14] = (PIPETX5EQCOEFF[14] !== 1'bz) && PIPETX5EQCOEFF_delay[14]; // rv 0
  assign PIPETX5EQCOEFF_in[15] = (PIPETX5EQCOEFF[15] !== 1'bz) && PIPETX5EQCOEFF_delay[15]; // rv 0
  assign PIPETX5EQCOEFF_in[16] = (PIPETX5EQCOEFF[16] !== 1'bz) && PIPETX5EQCOEFF_delay[16]; // rv 0
  assign PIPETX5EQCOEFF_in[17] = (PIPETX5EQCOEFF[17] !== 1'bz) && PIPETX5EQCOEFF_delay[17]; // rv 0
  assign PIPETX5EQCOEFF_in[1] = (PIPETX5EQCOEFF[1] !== 1'bz) && PIPETX5EQCOEFF_delay[1]; // rv 0
  assign PIPETX5EQCOEFF_in[2] = (PIPETX5EQCOEFF[2] !== 1'bz) && PIPETX5EQCOEFF_delay[2]; // rv 0
  assign PIPETX5EQCOEFF_in[3] = (PIPETX5EQCOEFF[3] !== 1'bz) && PIPETX5EQCOEFF_delay[3]; // rv 0
  assign PIPETX5EQCOEFF_in[4] = (PIPETX5EQCOEFF[4] !== 1'bz) && PIPETX5EQCOEFF_delay[4]; // rv 0
  assign PIPETX5EQCOEFF_in[5] = (PIPETX5EQCOEFF[5] !== 1'bz) && PIPETX5EQCOEFF_delay[5]; // rv 0
  assign PIPETX5EQCOEFF_in[6] = (PIPETX5EQCOEFF[6] !== 1'bz) && PIPETX5EQCOEFF_delay[6]; // rv 0
  assign PIPETX5EQCOEFF_in[7] = (PIPETX5EQCOEFF[7] !== 1'bz) && PIPETX5EQCOEFF_delay[7]; // rv 0
  assign PIPETX5EQCOEFF_in[8] = (PIPETX5EQCOEFF[8] !== 1'bz) && PIPETX5EQCOEFF_delay[8]; // rv 0
  assign PIPETX5EQCOEFF_in[9] = (PIPETX5EQCOEFF[9] !== 1'bz) && PIPETX5EQCOEFF_delay[9]; // rv 0
  assign PIPETX5EQDONE_in = (PIPETX5EQDONE !== 1'bz) && PIPETX5EQDONE_delay; // rv 0
  assign PIPETX6EQCOEFF_in[0] = (PIPETX6EQCOEFF[0] !== 1'bz) && PIPETX6EQCOEFF_delay[0]; // rv 0
  assign PIPETX6EQCOEFF_in[10] = (PIPETX6EQCOEFF[10] !== 1'bz) && PIPETX6EQCOEFF_delay[10]; // rv 0
  assign PIPETX6EQCOEFF_in[11] = (PIPETX6EQCOEFF[11] !== 1'bz) && PIPETX6EQCOEFF_delay[11]; // rv 0
  assign PIPETX6EQCOEFF_in[12] = (PIPETX6EQCOEFF[12] !== 1'bz) && PIPETX6EQCOEFF_delay[12]; // rv 0
  assign PIPETX6EQCOEFF_in[13] = (PIPETX6EQCOEFF[13] !== 1'bz) && PIPETX6EQCOEFF_delay[13]; // rv 0
  assign PIPETX6EQCOEFF_in[14] = (PIPETX6EQCOEFF[14] !== 1'bz) && PIPETX6EQCOEFF_delay[14]; // rv 0
  assign PIPETX6EQCOEFF_in[15] = (PIPETX6EQCOEFF[15] !== 1'bz) && PIPETX6EQCOEFF_delay[15]; // rv 0
  assign PIPETX6EQCOEFF_in[16] = (PIPETX6EQCOEFF[16] !== 1'bz) && PIPETX6EQCOEFF_delay[16]; // rv 0
  assign PIPETX6EQCOEFF_in[17] = (PIPETX6EQCOEFF[17] !== 1'bz) && PIPETX6EQCOEFF_delay[17]; // rv 0
  assign PIPETX6EQCOEFF_in[1] = (PIPETX6EQCOEFF[1] !== 1'bz) && PIPETX6EQCOEFF_delay[1]; // rv 0
  assign PIPETX6EQCOEFF_in[2] = (PIPETX6EQCOEFF[2] !== 1'bz) && PIPETX6EQCOEFF_delay[2]; // rv 0
  assign PIPETX6EQCOEFF_in[3] = (PIPETX6EQCOEFF[3] !== 1'bz) && PIPETX6EQCOEFF_delay[3]; // rv 0
  assign PIPETX6EQCOEFF_in[4] = (PIPETX6EQCOEFF[4] !== 1'bz) && PIPETX6EQCOEFF_delay[4]; // rv 0
  assign PIPETX6EQCOEFF_in[5] = (PIPETX6EQCOEFF[5] !== 1'bz) && PIPETX6EQCOEFF_delay[5]; // rv 0
  assign PIPETX6EQCOEFF_in[6] = (PIPETX6EQCOEFF[6] !== 1'bz) && PIPETX6EQCOEFF_delay[6]; // rv 0
  assign PIPETX6EQCOEFF_in[7] = (PIPETX6EQCOEFF[7] !== 1'bz) && PIPETX6EQCOEFF_delay[7]; // rv 0
  assign PIPETX6EQCOEFF_in[8] = (PIPETX6EQCOEFF[8] !== 1'bz) && PIPETX6EQCOEFF_delay[8]; // rv 0
  assign PIPETX6EQCOEFF_in[9] = (PIPETX6EQCOEFF[9] !== 1'bz) && PIPETX6EQCOEFF_delay[9]; // rv 0
  assign PIPETX6EQDONE_in = (PIPETX6EQDONE !== 1'bz) && PIPETX6EQDONE_delay; // rv 0
  assign PIPETX7EQCOEFF_in[0] = (PIPETX7EQCOEFF[0] !== 1'bz) && PIPETX7EQCOEFF_delay[0]; // rv 0
  assign PIPETX7EQCOEFF_in[10] = (PIPETX7EQCOEFF[10] !== 1'bz) && PIPETX7EQCOEFF_delay[10]; // rv 0
  assign PIPETX7EQCOEFF_in[11] = (PIPETX7EQCOEFF[11] !== 1'bz) && PIPETX7EQCOEFF_delay[11]; // rv 0
  assign PIPETX7EQCOEFF_in[12] = (PIPETX7EQCOEFF[12] !== 1'bz) && PIPETX7EQCOEFF_delay[12]; // rv 0
  assign PIPETX7EQCOEFF_in[13] = (PIPETX7EQCOEFF[13] !== 1'bz) && PIPETX7EQCOEFF_delay[13]; // rv 0
  assign PIPETX7EQCOEFF_in[14] = (PIPETX7EQCOEFF[14] !== 1'bz) && PIPETX7EQCOEFF_delay[14]; // rv 0
  assign PIPETX7EQCOEFF_in[15] = (PIPETX7EQCOEFF[15] !== 1'bz) && PIPETX7EQCOEFF_delay[15]; // rv 0
  assign PIPETX7EQCOEFF_in[16] = (PIPETX7EQCOEFF[16] !== 1'bz) && PIPETX7EQCOEFF_delay[16]; // rv 0
  assign PIPETX7EQCOEFF_in[17] = (PIPETX7EQCOEFF[17] !== 1'bz) && PIPETX7EQCOEFF_delay[17]; // rv 0
  assign PIPETX7EQCOEFF_in[1] = (PIPETX7EQCOEFF[1] !== 1'bz) && PIPETX7EQCOEFF_delay[1]; // rv 0
  assign PIPETX7EQCOEFF_in[2] = (PIPETX7EQCOEFF[2] !== 1'bz) && PIPETX7EQCOEFF_delay[2]; // rv 0
  assign PIPETX7EQCOEFF_in[3] = (PIPETX7EQCOEFF[3] !== 1'bz) && PIPETX7EQCOEFF_delay[3]; // rv 0
  assign PIPETX7EQCOEFF_in[4] = (PIPETX7EQCOEFF[4] !== 1'bz) && PIPETX7EQCOEFF_delay[4]; // rv 0
  assign PIPETX7EQCOEFF_in[5] = (PIPETX7EQCOEFF[5] !== 1'bz) && PIPETX7EQCOEFF_delay[5]; // rv 0
  assign PIPETX7EQCOEFF_in[6] = (PIPETX7EQCOEFF[6] !== 1'bz) && PIPETX7EQCOEFF_delay[6]; // rv 0
  assign PIPETX7EQCOEFF_in[7] = (PIPETX7EQCOEFF[7] !== 1'bz) && PIPETX7EQCOEFF_delay[7]; // rv 0
  assign PIPETX7EQCOEFF_in[8] = (PIPETX7EQCOEFF[8] !== 1'bz) && PIPETX7EQCOEFF_delay[8]; // rv 0
  assign PIPETX7EQCOEFF_in[9] = (PIPETX7EQCOEFF[9] !== 1'bz) && PIPETX7EQCOEFF_delay[9]; // rv 0
  assign PIPETX7EQDONE_in = (PIPETX7EQDONE !== 1'bz) && PIPETX7EQDONE_delay; // rv 0
  assign PLEQRESETEIEOSCOUNT_in = (PLEQRESETEIEOSCOUNT !== 1'bz) && PLEQRESETEIEOSCOUNT_delay; // rv 0
  assign PLGEN2UPSTREAMPREFERDEEMPH_in = (PLGEN2UPSTREAMPREFERDEEMPH !== 1'bz) && PLGEN2UPSTREAMPREFERDEEMPH_delay; // rv 0
  assign RESETN_in = (RESETN !== 1'bz) && RESETN_delay; // rv 0
  assign SAXISCCTDATA_in[0] = (SAXISCCTDATA[0] === 1'bz) || SAXISCCTDATA_delay[0]; // rv 1
  assign SAXISCCTDATA_in[100] = (SAXISCCTDATA[100] === 1'bz) || SAXISCCTDATA_delay[100]; // rv 1
  assign SAXISCCTDATA_in[101] = (SAXISCCTDATA[101] === 1'bz) || SAXISCCTDATA_delay[101]; // rv 1
  assign SAXISCCTDATA_in[102] = (SAXISCCTDATA[102] === 1'bz) || SAXISCCTDATA_delay[102]; // rv 1
  assign SAXISCCTDATA_in[103] = (SAXISCCTDATA[103] === 1'bz) || SAXISCCTDATA_delay[103]; // rv 1
  assign SAXISCCTDATA_in[104] = (SAXISCCTDATA[104] === 1'bz) || SAXISCCTDATA_delay[104]; // rv 1
  assign SAXISCCTDATA_in[105] = (SAXISCCTDATA[105] === 1'bz) || SAXISCCTDATA_delay[105]; // rv 1
  assign SAXISCCTDATA_in[106] = (SAXISCCTDATA[106] === 1'bz) || SAXISCCTDATA_delay[106]; // rv 1
  assign SAXISCCTDATA_in[107] = (SAXISCCTDATA[107] === 1'bz) || SAXISCCTDATA_delay[107]; // rv 1
  assign SAXISCCTDATA_in[108] = (SAXISCCTDATA[108] === 1'bz) || SAXISCCTDATA_delay[108]; // rv 1
  assign SAXISCCTDATA_in[109] = (SAXISCCTDATA[109] === 1'bz) || SAXISCCTDATA_delay[109]; // rv 1
  assign SAXISCCTDATA_in[10] = (SAXISCCTDATA[10] === 1'bz) || SAXISCCTDATA_delay[10]; // rv 1
  assign SAXISCCTDATA_in[110] = (SAXISCCTDATA[110] === 1'bz) || SAXISCCTDATA_delay[110]; // rv 1
  assign SAXISCCTDATA_in[111] = (SAXISCCTDATA[111] === 1'bz) || SAXISCCTDATA_delay[111]; // rv 1
  assign SAXISCCTDATA_in[112] = (SAXISCCTDATA[112] === 1'bz) || SAXISCCTDATA_delay[112]; // rv 1
  assign SAXISCCTDATA_in[113] = (SAXISCCTDATA[113] === 1'bz) || SAXISCCTDATA_delay[113]; // rv 1
  assign SAXISCCTDATA_in[114] = (SAXISCCTDATA[114] === 1'bz) || SAXISCCTDATA_delay[114]; // rv 1
  assign SAXISCCTDATA_in[115] = (SAXISCCTDATA[115] === 1'bz) || SAXISCCTDATA_delay[115]; // rv 1
  assign SAXISCCTDATA_in[116] = (SAXISCCTDATA[116] === 1'bz) || SAXISCCTDATA_delay[116]; // rv 1
  assign SAXISCCTDATA_in[117] = (SAXISCCTDATA[117] === 1'bz) || SAXISCCTDATA_delay[117]; // rv 1
  assign SAXISCCTDATA_in[118] = (SAXISCCTDATA[118] === 1'bz) || SAXISCCTDATA_delay[118]; // rv 1
  assign SAXISCCTDATA_in[119] = (SAXISCCTDATA[119] === 1'bz) || SAXISCCTDATA_delay[119]; // rv 1
  assign SAXISCCTDATA_in[11] = (SAXISCCTDATA[11] === 1'bz) || SAXISCCTDATA_delay[11]; // rv 1
  assign SAXISCCTDATA_in[120] = (SAXISCCTDATA[120] === 1'bz) || SAXISCCTDATA_delay[120]; // rv 1
  assign SAXISCCTDATA_in[121] = (SAXISCCTDATA[121] === 1'bz) || SAXISCCTDATA_delay[121]; // rv 1
  assign SAXISCCTDATA_in[122] = (SAXISCCTDATA[122] === 1'bz) || SAXISCCTDATA_delay[122]; // rv 1
  assign SAXISCCTDATA_in[123] = (SAXISCCTDATA[123] === 1'bz) || SAXISCCTDATA_delay[123]; // rv 1
  assign SAXISCCTDATA_in[124] = (SAXISCCTDATA[124] === 1'bz) || SAXISCCTDATA_delay[124]; // rv 1
  assign SAXISCCTDATA_in[125] = (SAXISCCTDATA[125] === 1'bz) || SAXISCCTDATA_delay[125]; // rv 1
  assign SAXISCCTDATA_in[126] = (SAXISCCTDATA[126] === 1'bz) || SAXISCCTDATA_delay[126]; // rv 1
  assign SAXISCCTDATA_in[127] = (SAXISCCTDATA[127] === 1'bz) || SAXISCCTDATA_delay[127]; // rv 1
  assign SAXISCCTDATA_in[128] = (SAXISCCTDATA[128] === 1'bz) || SAXISCCTDATA_delay[128]; // rv 1
  assign SAXISCCTDATA_in[129] = (SAXISCCTDATA[129] === 1'bz) || SAXISCCTDATA_delay[129]; // rv 1
  assign SAXISCCTDATA_in[12] = (SAXISCCTDATA[12] === 1'bz) || SAXISCCTDATA_delay[12]; // rv 1
  assign SAXISCCTDATA_in[130] = (SAXISCCTDATA[130] === 1'bz) || SAXISCCTDATA_delay[130]; // rv 1
  assign SAXISCCTDATA_in[131] = (SAXISCCTDATA[131] === 1'bz) || SAXISCCTDATA_delay[131]; // rv 1
  assign SAXISCCTDATA_in[132] = (SAXISCCTDATA[132] === 1'bz) || SAXISCCTDATA_delay[132]; // rv 1
  assign SAXISCCTDATA_in[133] = (SAXISCCTDATA[133] === 1'bz) || SAXISCCTDATA_delay[133]; // rv 1
  assign SAXISCCTDATA_in[134] = (SAXISCCTDATA[134] === 1'bz) || SAXISCCTDATA_delay[134]; // rv 1
  assign SAXISCCTDATA_in[135] = (SAXISCCTDATA[135] === 1'bz) || SAXISCCTDATA_delay[135]; // rv 1
  assign SAXISCCTDATA_in[136] = (SAXISCCTDATA[136] === 1'bz) || SAXISCCTDATA_delay[136]; // rv 1
  assign SAXISCCTDATA_in[137] = (SAXISCCTDATA[137] === 1'bz) || SAXISCCTDATA_delay[137]; // rv 1
  assign SAXISCCTDATA_in[138] = (SAXISCCTDATA[138] === 1'bz) || SAXISCCTDATA_delay[138]; // rv 1
  assign SAXISCCTDATA_in[139] = (SAXISCCTDATA[139] === 1'bz) || SAXISCCTDATA_delay[139]; // rv 1
  assign SAXISCCTDATA_in[13] = (SAXISCCTDATA[13] === 1'bz) || SAXISCCTDATA_delay[13]; // rv 1
  assign SAXISCCTDATA_in[140] = (SAXISCCTDATA[140] === 1'bz) || SAXISCCTDATA_delay[140]; // rv 1
  assign SAXISCCTDATA_in[141] = (SAXISCCTDATA[141] === 1'bz) || SAXISCCTDATA_delay[141]; // rv 1
  assign SAXISCCTDATA_in[142] = (SAXISCCTDATA[142] === 1'bz) || SAXISCCTDATA_delay[142]; // rv 1
  assign SAXISCCTDATA_in[143] = (SAXISCCTDATA[143] === 1'bz) || SAXISCCTDATA_delay[143]; // rv 1
  assign SAXISCCTDATA_in[144] = (SAXISCCTDATA[144] === 1'bz) || SAXISCCTDATA_delay[144]; // rv 1
  assign SAXISCCTDATA_in[145] = (SAXISCCTDATA[145] === 1'bz) || SAXISCCTDATA_delay[145]; // rv 1
  assign SAXISCCTDATA_in[146] = (SAXISCCTDATA[146] === 1'bz) || SAXISCCTDATA_delay[146]; // rv 1
  assign SAXISCCTDATA_in[147] = (SAXISCCTDATA[147] === 1'bz) || SAXISCCTDATA_delay[147]; // rv 1
  assign SAXISCCTDATA_in[148] = (SAXISCCTDATA[148] === 1'bz) || SAXISCCTDATA_delay[148]; // rv 1
  assign SAXISCCTDATA_in[149] = (SAXISCCTDATA[149] === 1'bz) || SAXISCCTDATA_delay[149]; // rv 1
  assign SAXISCCTDATA_in[14] = (SAXISCCTDATA[14] === 1'bz) || SAXISCCTDATA_delay[14]; // rv 1
  assign SAXISCCTDATA_in[150] = (SAXISCCTDATA[150] === 1'bz) || SAXISCCTDATA_delay[150]; // rv 1
  assign SAXISCCTDATA_in[151] = (SAXISCCTDATA[151] === 1'bz) || SAXISCCTDATA_delay[151]; // rv 1
  assign SAXISCCTDATA_in[152] = (SAXISCCTDATA[152] === 1'bz) || SAXISCCTDATA_delay[152]; // rv 1
  assign SAXISCCTDATA_in[153] = (SAXISCCTDATA[153] === 1'bz) || SAXISCCTDATA_delay[153]; // rv 1
  assign SAXISCCTDATA_in[154] = (SAXISCCTDATA[154] === 1'bz) || SAXISCCTDATA_delay[154]; // rv 1
  assign SAXISCCTDATA_in[155] = (SAXISCCTDATA[155] === 1'bz) || SAXISCCTDATA_delay[155]; // rv 1
  assign SAXISCCTDATA_in[156] = (SAXISCCTDATA[156] === 1'bz) || SAXISCCTDATA_delay[156]; // rv 1
  assign SAXISCCTDATA_in[157] = (SAXISCCTDATA[157] === 1'bz) || SAXISCCTDATA_delay[157]; // rv 1
  assign SAXISCCTDATA_in[158] = (SAXISCCTDATA[158] === 1'bz) || SAXISCCTDATA_delay[158]; // rv 1
  assign SAXISCCTDATA_in[159] = (SAXISCCTDATA[159] === 1'bz) || SAXISCCTDATA_delay[159]; // rv 1
  assign SAXISCCTDATA_in[15] = (SAXISCCTDATA[15] === 1'bz) || SAXISCCTDATA_delay[15]; // rv 1
  assign SAXISCCTDATA_in[160] = (SAXISCCTDATA[160] === 1'bz) || SAXISCCTDATA_delay[160]; // rv 1
  assign SAXISCCTDATA_in[161] = (SAXISCCTDATA[161] === 1'bz) || SAXISCCTDATA_delay[161]; // rv 1
  assign SAXISCCTDATA_in[162] = (SAXISCCTDATA[162] === 1'bz) || SAXISCCTDATA_delay[162]; // rv 1
  assign SAXISCCTDATA_in[163] = (SAXISCCTDATA[163] === 1'bz) || SAXISCCTDATA_delay[163]; // rv 1
  assign SAXISCCTDATA_in[164] = (SAXISCCTDATA[164] === 1'bz) || SAXISCCTDATA_delay[164]; // rv 1
  assign SAXISCCTDATA_in[165] = (SAXISCCTDATA[165] === 1'bz) || SAXISCCTDATA_delay[165]; // rv 1
  assign SAXISCCTDATA_in[166] = (SAXISCCTDATA[166] === 1'bz) || SAXISCCTDATA_delay[166]; // rv 1
  assign SAXISCCTDATA_in[167] = (SAXISCCTDATA[167] === 1'bz) || SAXISCCTDATA_delay[167]; // rv 1
  assign SAXISCCTDATA_in[168] = (SAXISCCTDATA[168] === 1'bz) || SAXISCCTDATA_delay[168]; // rv 1
  assign SAXISCCTDATA_in[169] = (SAXISCCTDATA[169] === 1'bz) || SAXISCCTDATA_delay[169]; // rv 1
  assign SAXISCCTDATA_in[16] = (SAXISCCTDATA[16] === 1'bz) || SAXISCCTDATA_delay[16]; // rv 1
  assign SAXISCCTDATA_in[170] = (SAXISCCTDATA[170] === 1'bz) || SAXISCCTDATA_delay[170]; // rv 1
  assign SAXISCCTDATA_in[171] = (SAXISCCTDATA[171] === 1'bz) || SAXISCCTDATA_delay[171]; // rv 1
  assign SAXISCCTDATA_in[172] = (SAXISCCTDATA[172] === 1'bz) || SAXISCCTDATA_delay[172]; // rv 1
  assign SAXISCCTDATA_in[173] = (SAXISCCTDATA[173] === 1'bz) || SAXISCCTDATA_delay[173]; // rv 1
  assign SAXISCCTDATA_in[174] = (SAXISCCTDATA[174] === 1'bz) || SAXISCCTDATA_delay[174]; // rv 1
  assign SAXISCCTDATA_in[175] = (SAXISCCTDATA[175] === 1'bz) || SAXISCCTDATA_delay[175]; // rv 1
  assign SAXISCCTDATA_in[176] = (SAXISCCTDATA[176] === 1'bz) || SAXISCCTDATA_delay[176]; // rv 1
  assign SAXISCCTDATA_in[177] = (SAXISCCTDATA[177] === 1'bz) || SAXISCCTDATA_delay[177]; // rv 1
  assign SAXISCCTDATA_in[178] = (SAXISCCTDATA[178] === 1'bz) || SAXISCCTDATA_delay[178]; // rv 1
  assign SAXISCCTDATA_in[179] = (SAXISCCTDATA[179] === 1'bz) || SAXISCCTDATA_delay[179]; // rv 1
  assign SAXISCCTDATA_in[17] = (SAXISCCTDATA[17] === 1'bz) || SAXISCCTDATA_delay[17]; // rv 1
  assign SAXISCCTDATA_in[180] = (SAXISCCTDATA[180] === 1'bz) || SAXISCCTDATA_delay[180]; // rv 1
  assign SAXISCCTDATA_in[181] = (SAXISCCTDATA[181] === 1'bz) || SAXISCCTDATA_delay[181]; // rv 1
  assign SAXISCCTDATA_in[182] = (SAXISCCTDATA[182] === 1'bz) || SAXISCCTDATA_delay[182]; // rv 1
  assign SAXISCCTDATA_in[183] = (SAXISCCTDATA[183] === 1'bz) || SAXISCCTDATA_delay[183]; // rv 1
  assign SAXISCCTDATA_in[184] = (SAXISCCTDATA[184] === 1'bz) || SAXISCCTDATA_delay[184]; // rv 1
  assign SAXISCCTDATA_in[185] = (SAXISCCTDATA[185] === 1'bz) || SAXISCCTDATA_delay[185]; // rv 1
  assign SAXISCCTDATA_in[186] = (SAXISCCTDATA[186] === 1'bz) || SAXISCCTDATA_delay[186]; // rv 1
  assign SAXISCCTDATA_in[187] = (SAXISCCTDATA[187] === 1'bz) || SAXISCCTDATA_delay[187]; // rv 1
  assign SAXISCCTDATA_in[188] = (SAXISCCTDATA[188] === 1'bz) || SAXISCCTDATA_delay[188]; // rv 1
  assign SAXISCCTDATA_in[189] = (SAXISCCTDATA[189] === 1'bz) || SAXISCCTDATA_delay[189]; // rv 1
  assign SAXISCCTDATA_in[18] = (SAXISCCTDATA[18] === 1'bz) || SAXISCCTDATA_delay[18]; // rv 1
  assign SAXISCCTDATA_in[190] = (SAXISCCTDATA[190] === 1'bz) || SAXISCCTDATA_delay[190]; // rv 1
  assign SAXISCCTDATA_in[191] = (SAXISCCTDATA[191] === 1'bz) || SAXISCCTDATA_delay[191]; // rv 1
  assign SAXISCCTDATA_in[192] = (SAXISCCTDATA[192] === 1'bz) || SAXISCCTDATA_delay[192]; // rv 1
  assign SAXISCCTDATA_in[193] = (SAXISCCTDATA[193] === 1'bz) || SAXISCCTDATA_delay[193]; // rv 1
  assign SAXISCCTDATA_in[194] = (SAXISCCTDATA[194] === 1'bz) || SAXISCCTDATA_delay[194]; // rv 1
  assign SAXISCCTDATA_in[195] = (SAXISCCTDATA[195] === 1'bz) || SAXISCCTDATA_delay[195]; // rv 1
  assign SAXISCCTDATA_in[196] = (SAXISCCTDATA[196] === 1'bz) || SAXISCCTDATA_delay[196]; // rv 1
  assign SAXISCCTDATA_in[197] = (SAXISCCTDATA[197] === 1'bz) || SAXISCCTDATA_delay[197]; // rv 1
  assign SAXISCCTDATA_in[198] = (SAXISCCTDATA[198] === 1'bz) || SAXISCCTDATA_delay[198]; // rv 1
  assign SAXISCCTDATA_in[199] = (SAXISCCTDATA[199] === 1'bz) || SAXISCCTDATA_delay[199]; // rv 1
  assign SAXISCCTDATA_in[19] = (SAXISCCTDATA[19] === 1'bz) || SAXISCCTDATA_delay[19]; // rv 1
  assign SAXISCCTDATA_in[1] = (SAXISCCTDATA[1] === 1'bz) || SAXISCCTDATA_delay[1]; // rv 1
  assign SAXISCCTDATA_in[200] = (SAXISCCTDATA[200] === 1'bz) || SAXISCCTDATA_delay[200]; // rv 1
  assign SAXISCCTDATA_in[201] = (SAXISCCTDATA[201] === 1'bz) || SAXISCCTDATA_delay[201]; // rv 1
  assign SAXISCCTDATA_in[202] = (SAXISCCTDATA[202] === 1'bz) || SAXISCCTDATA_delay[202]; // rv 1
  assign SAXISCCTDATA_in[203] = (SAXISCCTDATA[203] === 1'bz) || SAXISCCTDATA_delay[203]; // rv 1
  assign SAXISCCTDATA_in[204] = (SAXISCCTDATA[204] === 1'bz) || SAXISCCTDATA_delay[204]; // rv 1
  assign SAXISCCTDATA_in[205] = (SAXISCCTDATA[205] === 1'bz) || SAXISCCTDATA_delay[205]; // rv 1
  assign SAXISCCTDATA_in[206] = (SAXISCCTDATA[206] === 1'bz) || SAXISCCTDATA_delay[206]; // rv 1
  assign SAXISCCTDATA_in[207] = (SAXISCCTDATA[207] === 1'bz) || SAXISCCTDATA_delay[207]; // rv 1
  assign SAXISCCTDATA_in[208] = (SAXISCCTDATA[208] === 1'bz) || SAXISCCTDATA_delay[208]; // rv 1
  assign SAXISCCTDATA_in[209] = (SAXISCCTDATA[209] === 1'bz) || SAXISCCTDATA_delay[209]; // rv 1
  assign SAXISCCTDATA_in[20] = (SAXISCCTDATA[20] === 1'bz) || SAXISCCTDATA_delay[20]; // rv 1
  assign SAXISCCTDATA_in[210] = (SAXISCCTDATA[210] === 1'bz) || SAXISCCTDATA_delay[210]; // rv 1
  assign SAXISCCTDATA_in[211] = (SAXISCCTDATA[211] === 1'bz) || SAXISCCTDATA_delay[211]; // rv 1
  assign SAXISCCTDATA_in[212] = (SAXISCCTDATA[212] === 1'bz) || SAXISCCTDATA_delay[212]; // rv 1
  assign SAXISCCTDATA_in[213] = (SAXISCCTDATA[213] === 1'bz) || SAXISCCTDATA_delay[213]; // rv 1
  assign SAXISCCTDATA_in[214] = (SAXISCCTDATA[214] === 1'bz) || SAXISCCTDATA_delay[214]; // rv 1
  assign SAXISCCTDATA_in[215] = (SAXISCCTDATA[215] === 1'bz) || SAXISCCTDATA_delay[215]; // rv 1
  assign SAXISCCTDATA_in[216] = (SAXISCCTDATA[216] === 1'bz) || SAXISCCTDATA_delay[216]; // rv 1
  assign SAXISCCTDATA_in[217] = (SAXISCCTDATA[217] === 1'bz) || SAXISCCTDATA_delay[217]; // rv 1
  assign SAXISCCTDATA_in[218] = (SAXISCCTDATA[218] === 1'bz) || SAXISCCTDATA_delay[218]; // rv 1
  assign SAXISCCTDATA_in[219] = (SAXISCCTDATA[219] === 1'bz) || SAXISCCTDATA_delay[219]; // rv 1
  assign SAXISCCTDATA_in[21] = (SAXISCCTDATA[21] === 1'bz) || SAXISCCTDATA_delay[21]; // rv 1
  assign SAXISCCTDATA_in[220] = (SAXISCCTDATA[220] === 1'bz) || SAXISCCTDATA_delay[220]; // rv 1
  assign SAXISCCTDATA_in[221] = (SAXISCCTDATA[221] === 1'bz) || SAXISCCTDATA_delay[221]; // rv 1
  assign SAXISCCTDATA_in[222] = (SAXISCCTDATA[222] === 1'bz) || SAXISCCTDATA_delay[222]; // rv 1
  assign SAXISCCTDATA_in[223] = (SAXISCCTDATA[223] === 1'bz) || SAXISCCTDATA_delay[223]; // rv 1
  assign SAXISCCTDATA_in[224] = (SAXISCCTDATA[224] === 1'bz) || SAXISCCTDATA_delay[224]; // rv 1
  assign SAXISCCTDATA_in[225] = (SAXISCCTDATA[225] === 1'bz) || SAXISCCTDATA_delay[225]; // rv 1
  assign SAXISCCTDATA_in[226] = (SAXISCCTDATA[226] === 1'bz) || SAXISCCTDATA_delay[226]; // rv 1
  assign SAXISCCTDATA_in[227] = (SAXISCCTDATA[227] === 1'bz) || SAXISCCTDATA_delay[227]; // rv 1
  assign SAXISCCTDATA_in[228] = (SAXISCCTDATA[228] === 1'bz) || SAXISCCTDATA_delay[228]; // rv 1
  assign SAXISCCTDATA_in[229] = (SAXISCCTDATA[229] === 1'bz) || SAXISCCTDATA_delay[229]; // rv 1
  assign SAXISCCTDATA_in[22] = (SAXISCCTDATA[22] === 1'bz) || SAXISCCTDATA_delay[22]; // rv 1
  assign SAXISCCTDATA_in[230] = (SAXISCCTDATA[230] === 1'bz) || SAXISCCTDATA_delay[230]; // rv 1
  assign SAXISCCTDATA_in[231] = (SAXISCCTDATA[231] === 1'bz) || SAXISCCTDATA_delay[231]; // rv 1
  assign SAXISCCTDATA_in[232] = (SAXISCCTDATA[232] === 1'bz) || SAXISCCTDATA_delay[232]; // rv 1
  assign SAXISCCTDATA_in[233] = (SAXISCCTDATA[233] === 1'bz) || SAXISCCTDATA_delay[233]; // rv 1
  assign SAXISCCTDATA_in[234] = (SAXISCCTDATA[234] === 1'bz) || SAXISCCTDATA_delay[234]; // rv 1
  assign SAXISCCTDATA_in[235] = (SAXISCCTDATA[235] === 1'bz) || SAXISCCTDATA_delay[235]; // rv 1
  assign SAXISCCTDATA_in[236] = (SAXISCCTDATA[236] === 1'bz) || SAXISCCTDATA_delay[236]; // rv 1
  assign SAXISCCTDATA_in[237] = (SAXISCCTDATA[237] === 1'bz) || SAXISCCTDATA_delay[237]; // rv 1
  assign SAXISCCTDATA_in[238] = (SAXISCCTDATA[238] === 1'bz) || SAXISCCTDATA_delay[238]; // rv 1
  assign SAXISCCTDATA_in[239] = (SAXISCCTDATA[239] === 1'bz) || SAXISCCTDATA_delay[239]; // rv 1
  assign SAXISCCTDATA_in[23] = (SAXISCCTDATA[23] === 1'bz) || SAXISCCTDATA_delay[23]; // rv 1
  assign SAXISCCTDATA_in[240] = (SAXISCCTDATA[240] === 1'bz) || SAXISCCTDATA_delay[240]; // rv 1
  assign SAXISCCTDATA_in[241] = (SAXISCCTDATA[241] === 1'bz) || SAXISCCTDATA_delay[241]; // rv 1
  assign SAXISCCTDATA_in[242] = (SAXISCCTDATA[242] === 1'bz) || SAXISCCTDATA_delay[242]; // rv 1
  assign SAXISCCTDATA_in[243] = (SAXISCCTDATA[243] === 1'bz) || SAXISCCTDATA_delay[243]; // rv 1
  assign SAXISCCTDATA_in[244] = (SAXISCCTDATA[244] === 1'bz) || SAXISCCTDATA_delay[244]; // rv 1
  assign SAXISCCTDATA_in[245] = (SAXISCCTDATA[245] === 1'bz) || SAXISCCTDATA_delay[245]; // rv 1
  assign SAXISCCTDATA_in[246] = (SAXISCCTDATA[246] === 1'bz) || SAXISCCTDATA_delay[246]; // rv 1
  assign SAXISCCTDATA_in[247] = (SAXISCCTDATA[247] === 1'bz) || SAXISCCTDATA_delay[247]; // rv 1
  assign SAXISCCTDATA_in[248] = (SAXISCCTDATA[248] === 1'bz) || SAXISCCTDATA_delay[248]; // rv 1
  assign SAXISCCTDATA_in[249] = (SAXISCCTDATA[249] === 1'bz) || SAXISCCTDATA_delay[249]; // rv 1
  assign SAXISCCTDATA_in[24] = (SAXISCCTDATA[24] === 1'bz) || SAXISCCTDATA_delay[24]; // rv 1
  assign SAXISCCTDATA_in[250] = (SAXISCCTDATA[250] === 1'bz) || SAXISCCTDATA_delay[250]; // rv 1
  assign SAXISCCTDATA_in[251] = (SAXISCCTDATA[251] === 1'bz) || SAXISCCTDATA_delay[251]; // rv 1
  assign SAXISCCTDATA_in[252] = (SAXISCCTDATA[252] === 1'bz) || SAXISCCTDATA_delay[252]; // rv 1
  assign SAXISCCTDATA_in[253] = (SAXISCCTDATA[253] === 1'bz) || SAXISCCTDATA_delay[253]; // rv 1
  assign SAXISCCTDATA_in[254] = (SAXISCCTDATA[254] === 1'bz) || SAXISCCTDATA_delay[254]; // rv 1
  assign SAXISCCTDATA_in[255] = (SAXISCCTDATA[255] === 1'bz) || SAXISCCTDATA_delay[255]; // rv 1
  assign SAXISCCTDATA_in[25] = (SAXISCCTDATA[25] === 1'bz) || SAXISCCTDATA_delay[25]; // rv 1
  assign SAXISCCTDATA_in[26] = (SAXISCCTDATA[26] === 1'bz) || SAXISCCTDATA_delay[26]; // rv 1
  assign SAXISCCTDATA_in[27] = (SAXISCCTDATA[27] === 1'bz) || SAXISCCTDATA_delay[27]; // rv 1
  assign SAXISCCTDATA_in[28] = (SAXISCCTDATA[28] === 1'bz) || SAXISCCTDATA_delay[28]; // rv 1
  assign SAXISCCTDATA_in[29] = (SAXISCCTDATA[29] === 1'bz) || SAXISCCTDATA_delay[29]; // rv 1
  assign SAXISCCTDATA_in[2] = (SAXISCCTDATA[2] === 1'bz) || SAXISCCTDATA_delay[2]; // rv 1
  assign SAXISCCTDATA_in[30] = (SAXISCCTDATA[30] === 1'bz) || SAXISCCTDATA_delay[30]; // rv 1
  assign SAXISCCTDATA_in[31] = (SAXISCCTDATA[31] === 1'bz) || SAXISCCTDATA_delay[31]; // rv 1
  assign SAXISCCTDATA_in[32] = (SAXISCCTDATA[32] === 1'bz) || SAXISCCTDATA_delay[32]; // rv 1
  assign SAXISCCTDATA_in[33] = (SAXISCCTDATA[33] === 1'bz) || SAXISCCTDATA_delay[33]; // rv 1
  assign SAXISCCTDATA_in[34] = (SAXISCCTDATA[34] === 1'bz) || SAXISCCTDATA_delay[34]; // rv 1
  assign SAXISCCTDATA_in[35] = (SAXISCCTDATA[35] === 1'bz) || SAXISCCTDATA_delay[35]; // rv 1
  assign SAXISCCTDATA_in[36] = (SAXISCCTDATA[36] === 1'bz) || SAXISCCTDATA_delay[36]; // rv 1
  assign SAXISCCTDATA_in[37] = (SAXISCCTDATA[37] === 1'bz) || SAXISCCTDATA_delay[37]; // rv 1
  assign SAXISCCTDATA_in[38] = (SAXISCCTDATA[38] === 1'bz) || SAXISCCTDATA_delay[38]; // rv 1
  assign SAXISCCTDATA_in[39] = (SAXISCCTDATA[39] === 1'bz) || SAXISCCTDATA_delay[39]; // rv 1
  assign SAXISCCTDATA_in[3] = (SAXISCCTDATA[3] === 1'bz) || SAXISCCTDATA_delay[3]; // rv 1
  assign SAXISCCTDATA_in[40] = (SAXISCCTDATA[40] === 1'bz) || SAXISCCTDATA_delay[40]; // rv 1
  assign SAXISCCTDATA_in[41] = (SAXISCCTDATA[41] === 1'bz) || SAXISCCTDATA_delay[41]; // rv 1
  assign SAXISCCTDATA_in[42] = (SAXISCCTDATA[42] === 1'bz) || SAXISCCTDATA_delay[42]; // rv 1
  assign SAXISCCTDATA_in[43] = (SAXISCCTDATA[43] === 1'bz) || SAXISCCTDATA_delay[43]; // rv 1
  assign SAXISCCTDATA_in[44] = (SAXISCCTDATA[44] === 1'bz) || SAXISCCTDATA_delay[44]; // rv 1
  assign SAXISCCTDATA_in[45] = (SAXISCCTDATA[45] === 1'bz) || SAXISCCTDATA_delay[45]; // rv 1
  assign SAXISCCTDATA_in[46] = (SAXISCCTDATA[46] === 1'bz) || SAXISCCTDATA_delay[46]; // rv 1
  assign SAXISCCTDATA_in[47] = (SAXISCCTDATA[47] === 1'bz) || SAXISCCTDATA_delay[47]; // rv 1
  assign SAXISCCTDATA_in[48] = (SAXISCCTDATA[48] === 1'bz) || SAXISCCTDATA_delay[48]; // rv 1
  assign SAXISCCTDATA_in[49] = (SAXISCCTDATA[49] === 1'bz) || SAXISCCTDATA_delay[49]; // rv 1
  assign SAXISCCTDATA_in[4] = (SAXISCCTDATA[4] === 1'bz) || SAXISCCTDATA_delay[4]; // rv 1
  assign SAXISCCTDATA_in[50] = (SAXISCCTDATA[50] === 1'bz) || SAXISCCTDATA_delay[50]; // rv 1
  assign SAXISCCTDATA_in[51] = (SAXISCCTDATA[51] === 1'bz) || SAXISCCTDATA_delay[51]; // rv 1
  assign SAXISCCTDATA_in[52] = (SAXISCCTDATA[52] === 1'bz) || SAXISCCTDATA_delay[52]; // rv 1
  assign SAXISCCTDATA_in[53] = (SAXISCCTDATA[53] === 1'bz) || SAXISCCTDATA_delay[53]; // rv 1
  assign SAXISCCTDATA_in[54] = (SAXISCCTDATA[54] === 1'bz) || SAXISCCTDATA_delay[54]; // rv 1
  assign SAXISCCTDATA_in[55] = (SAXISCCTDATA[55] === 1'bz) || SAXISCCTDATA_delay[55]; // rv 1
  assign SAXISCCTDATA_in[56] = (SAXISCCTDATA[56] === 1'bz) || SAXISCCTDATA_delay[56]; // rv 1
  assign SAXISCCTDATA_in[57] = (SAXISCCTDATA[57] === 1'bz) || SAXISCCTDATA_delay[57]; // rv 1
  assign SAXISCCTDATA_in[58] = (SAXISCCTDATA[58] === 1'bz) || SAXISCCTDATA_delay[58]; // rv 1
  assign SAXISCCTDATA_in[59] = (SAXISCCTDATA[59] === 1'bz) || SAXISCCTDATA_delay[59]; // rv 1
  assign SAXISCCTDATA_in[5] = (SAXISCCTDATA[5] === 1'bz) || SAXISCCTDATA_delay[5]; // rv 1
  assign SAXISCCTDATA_in[60] = (SAXISCCTDATA[60] === 1'bz) || SAXISCCTDATA_delay[60]; // rv 1
  assign SAXISCCTDATA_in[61] = (SAXISCCTDATA[61] === 1'bz) || SAXISCCTDATA_delay[61]; // rv 1
  assign SAXISCCTDATA_in[62] = (SAXISCCTDATA[62] === 1'bz) || SAXISCCTDATA_delay[62]; // rv 1
  assign SAXISCCTDATA_in[63] = (SAXISCCTDATA[63] === 1'bz) || SAXISCCTDATA_delay[63]; // rv 1
  assign SAXISCCTDATA_in[64] = (SAXISCCTDATA[64] === 1'bz) || SAXISCCTDATA_delay[64]; // rv 1
  assign SAXISCCTDATA_in[65] = (SAXISCCTDATA[65] === 1'bz) || SAXISCCTDATA_delay[65]; // rv 1
  assign SAXISCCTDATA_in[66] = (SAXISCCTDATA[66] === 1'bz) || SAXISCCTDATA_delay[66]; // rv 1
  assign SAXISCCTDATA_in[67] = (SAXISCCTDATA[67] === 1'bz) || SAXISCCTDATA_delay[67]; // rv 1
  assign SAXISCCTDATA_in[68] = (SAXISCCTDATA[68] === 1'bz) || SAXISCCTDATA_delay[68]; // rv 1
  assign SAXISCCTDATA_in[69] = (SAXISCCTDATA[69] === 1'bz) || SAXISCCTDATA_delay[69]; // rv 1
  assign SAXISCCTDATA_in[6] = (SAXISCCTDATA[6] === 1'bz) || SAXISCCTDATA_delay[6]; // rv 1
  assign SAXISCCTDATA_in[70] = (SAXISCCTDATA[70] === 1'bz) || SAXISCCTDATA_delay[70]; // rv 1
  assign SAXISCCTDATA_in[71] = (SAXISCCTDATA[71] === 1'bz) || SAXISCCTDATA_delay[71]; // rv 1
  assign SAXISCCTDATA_in[72] = (SAXISCCTDATA[72] === 1'bz) || SAXISCCTDATA_delay[72]; // rv 1
  assign SAXISCCTDATA_in[73] = (SAXISCCTDATA[73] === 1'bz) || SAXISCCTDATA_delay[73]; // rv 1
  assign SAXISCCTDATA_in[74] = (SAXISCCTDATA[74] === 1'bz) || SAXISCCTDATA_delay[74]; // rv 1
  assign SAXISCCTDATA_in[75] = (SAXISCCTDATA[75] === 1'bz) || SAXISCCTDATA_delay[75]; // rv 1
  assign SAXISCCTDATA_in[76] = (SAXISCCTDATA[76] === 1'bz) || SAXISCCTDATA_delay[76]; // rv 1
  assign SAXISCCTDATA_in[77] = (SAXISCCTDATA[77] === 1'bz) || SAXISCCTDATA_delay[77]; // rv 1
  assign SAXISCCTDATA_in[78] = (SAXISCCTDATA[78] === 1'bz) || SAXISCCTDATA_delay[78]; // rv 1
  assign SAXISCCTDATA_in[79] = (SAXISCCTDATA[79] === 1'bz) || SAXISCCTDATA_delay[79]; // rv 1
  assign SAXISCCTDATA_in[7] = (SAXISCCTDATA[7] === 1'bz) || SAXISCCTDATA_delay[7]; // rv 1
  assign SAXISCCTDATA_in[80] = (SAXISCCTDATA[80] === 1'bz) || SAXISCCTDATA_delay[80]; // rv 1
  assign SAXISCCTDATA_in[81] = (SAXISCCTDATA[81] === 1'bz) || SAXISCCTDATA_delay[81]; // rv 1
  assign SAXISCCTDATA_in[82] = (SAXISCCTDATA[82] === 1'bz) || SAXISCCTDATA_delay[82]; // rv 1
  assign SAXISCCTDATA_in[83] = (SAXISCCTDATA[83] === 1'bz) || SAXISCCTDATA_delay[83]; // rv 1
  assign SAXISCCTDATA_in[84] = (SAXISCCTDATA[84] === 1'bz) || SAXISCCTDATA_delay[84]; // rv 1
  assign SAXISCCTDATA_in[85] = (SAXISCCTDATA[85] === 1'bz) || SAXISCCTDATA_delay[85]; // rv 1
  assign SAXISCCTDATA_in[86] = (SAXISCCTDATA[86] === 1'bz) || SAXISCCTDATA_delay[86]; // rv 1
  assign SAXISCCTDATA_in[87] = (SAXISCCTDATA[87] === 1'bz) || SAXISCCTDATA_delay[87]; // rv 1
  assign SAXISCCTDATA_in[88] = (SAXISCCTDATA[88] === 1'bz) || SAXISCCTDATA_delay[88]; // rv 1
  assign SAXISCCTDATA_in[89] = (SAXISCCTDATA[89] === 1'bz) || SAXISCCTDATA_delay[89]; // rv 1
  assign SAXISCCTDATA_in[8] = (SAXISCCTDATA[8] === 1'bz) || SAXISCCTDATA_delay[8]; // rv 1
  assign SAXISCCTDATA_in[90] = (SAXISCCTDATA[90] === 1'bz) || SAXISCCTDATA_delay[90]; // rv 1
  assign SAXISCCTDATA_in[91] = (SAXISCCTDATA[91] === 1'bz) || SAXISCCTDATA_delay[91]; // rv 1
  assign SAXISCCTDATA_in[92] = (SAXISCCTDATA[92] === 1'bz) || SAXISCCTDATA_delay[92]; // rv 1
  assign SAXISCCTDATA_in[93] = (SAXISCCTDATA[93] === 1'bz) || SAXISCCTDATA_delay[93]; // rv 1
  assign SAXISCCTDATA_in[94] = (SAXISCCTDATA[94] === 1'bz) || SAXISCCTDATA_delay[94]; // rv 1
  assign SAXISCCTDATA_in[95] = (SAXISCCTDATA[95] === 1'bz) || SAXISCCTDATA_delay[95]; // rv 1
  assign SAXISCCTDATA_in[96] = (SAXISCCTDATA[96] === 1'bz) || SAXISCCTDATA_delay[96]; // rv 1
  assign SAXISCCTDATA_in[97] = (SAXISCCTDATA[97] === 1'bz) || SAXISCCTDATA_delay[97]; // rv 1
  assign SAXISCCTDATA_in[98] = (SAXISCCTDATA[98] === 1'bz) || SAXISCCTDATA_delay[98]; // rv 1
  assign SAXISCCTDATA_in[99] = (SAXISCCTDATA[99] === 1'bz) || SAXISCCTDATA_delay[99]; // rv 1
  assign SAXISCCTDATA_in[9] = (SAXISCCTDATA[9] === 1'bz) || SAXISCCTDATA_delay[9]; // rv 1
  assign SAXISCCTKEEP_in[0] = (SAXISCCTKEEP[0] !== 1'bz) && SAXISCCTKEEP_delay[0]; // rv 0
  assign SAXISCCTKEEP_in[1] = (SAXISCCTKEEP[1] !== 1'bz) && SAXISCCTKEEP_delay[1]; // rv 0
  assign SAXISCCTKEEP_in[2] = (SAXISCCTKEEP[2] !== 1'bz) && SAXISCCTKEEP_delay[2]; // rv 0
  assign SAXISCCTKEEP_in[3] = (SAXISCCTKEEP[3] !== 1'bz) && SAXISCCTKEEP_delay[3]; // rv 0
  assign SAXISCCTKEEP_in[4] = (SAXISCCTKEEP[4] !== 1'bz) && SAXISCCTKEEP_delay[4]; // rv 0
  assign SAXISCCTKEEP_in[5] = (SAXISCCTKEEP[5] !== 1'bz) && SAXISCCTKEEP_delay[5]; // rv 0
  assign SAXISCCTKEEP_in[6] = (SAXISCCTKEEP[6] !== 1'bz) && SAXISCCTKEEP_delay[6]; // rv 0
  assign SAXISCCTKEEP_in[7] = (SAXISCCTKEEP[7] !== 1'bz) && SAXISCCTKEEP_delay[7]; // rv 0
  assign SAXISCCTLAST_in = (SAXISCCTLAST === 1'bz) || SAXISCCTLAST_delay; // rv 1
  assign SAXISCCTUSER_in[0] = (SAXISCCTUSER[0] === 1'bz) || SAXISCCTUSER_delay[0]; // rv 1
  assign SAXISCCTUSER_in[10] = (SAXISCCTUSER[10] === 1'bz) || SAXISCCTUSER_delay[10]; // rv 1
  assign SAXISCCTUSER_in[11] = (SAXISCCTUSER[11] === 1'bz) || SAXISCCTUSER_delay[11]; // rv 1
  assign SAXISCCTUSER_in[12] = (SAXISCCTUSER[12] === 1'bz) || SAXISCCTUSER_delay[12]; // rv 1
  assign SAXISCCTUSER_in[13] = (SAXISCCTUSER[13] === 1'bz) || SAXISCCTUSER_delay[13]; // rv 1
  assign SAXISCCTUSER_in[14] = (SAXISCCTUSER[14] === 1'bz) || SAXISCCTUSER_delay[14]; // rv 1
  assign SAXISCCTUSER_in[15] = (SAXISCCTUSER[15] === 1'bz) || SAXISCCTUSER_delay[15]; // rv 1
  assign SAXISCCTUSER_in[16] = (SAXISCCTUSER[16] === 1'bz) || SAXISCCTUSER_delay[16]; // rv 1
  assign SAXISCCTUSER_in[17] = (SAXISCCTUSER[17] === 1'bz) || SAXISCCTUSER_delay[17]; // rv 1
  assign SAXISCCTUSER_in[18] = (SAXISCCTUSER[18] === 1'bz) || SAXISCCTUSER_delay[18]; // rv 1
  assign SAXISCCTUSER_in[19] = (SAXISCCTUSER[19] === 1'bz) || SAXISCCTUSER_delay[19]; // rv 1
  assign SAXISCCTUSER_in[1] = (SAXISCCTUSER[1] === 1'bz) || SAXISCCTUSER_delay[1]; // rv 1
  assign SAXISCCTUSER_in[20] = (SAXISCCTUSER[20] === 1'bz) || SAXISCCTUSER_delay[20]; // rv 1
  assign SAXISCCTUSER_in[21] = (SAXISCCTUSER[21] === 1'bz) || SAXISCCTUSER_delay[21]; // rv 1
  assign SAXISCCTUSER_in[22] = (SAXISCCTUSER[22] === 1'bz) || SAXISCCTUSER_delay[22]; // rv 1
  assign SAXISCCTUSER_in[23] = (SAXISCCTUSER[23] === 1'bz) || SAXISCCTUSER_delay[23]; // rv 1
  assign SAXISCCTUSER_in[24] = (SAXISCCTUSER[24] === 1'bz) || SAXISCCTUSER_delay[24]; // rv 1
  assign SAXISCCTUSER_in[25] = (SAXISCCTUSER[25] === 1'bz) || SAXISCCTUSER_delay[25]; // rv 1
  assign SAXISCCTUSER_in[26] = (SAXISCCTUSER[26] === 1'bz) || SAXISCCTUSER_delay[26]; // rv 1
  assign SAXISCCTUSER_in[27] = (SAXISCCTUSER[27] === 1'bz) || SAXISCCTUSER_delay[27]; // rv 1
  assign SAXISCCTUSER_in[28] = (SAXISCCTUSER[28] === 1'bz) || SAXISCCTUSER_delay[28]; // rv 1
  assign SAXISCCTUSER_in[29] = (SAXISCCTUSER[29] === 1'bz) || SAXISCCTUSER_delay[29]; // rv 1
  assign SAXISCCTUSER_in[2] = (SAXISCCTUSER[2] === 1'bz) || SAXISCCTUSER_delay[2]; // rv 1
  assign SAXISCCTUSER_in[30] = (SAXISCCTUSER[30] === 1'bz) || SAXISCCTUSER_delay[30]; // rv 1
  assign SAXISCCTUSER_in[31] = (SAXISCCTUSER[31] === 1'bz) || SAXISCCTUSER_delay[31]; // rv 1
  assign SAXISCCTUSER_in[32] = (SAXISCCTUSER[32] === 1'bz) || SAXISCCTUSER_delay[32]; // rv 1
  assign SAXISCCTUSER_in[3] = (SAXISCCTUSER[3] === 1'bz) || SAXISCCTUSER_delay[3]; // rv 1
  assign SAXISCCTUSER_in[4] = (SAXISCCTUSER[4] === 1'bz) || SAXISCCTUSER_delay[4]; // rv 1
  assign SAXISCCTUSER_in[5] = (SAXISCCTUSER[5] === 1'bz) || SAXISCCTUSER_delay[5]; // rv 1
  assign SAXISCCTUSER_in[6] = (SAXISCCTUSER[6] === 1'bz) || SAXISCCTUSER_delay[6]; // rv 1
  assign SAXISCCTUSER_in[7] = (SAXISCCTUSER[7] === 1'bz) || SAXISCCTUSER_delay[7]; // rv 1
  assign SAXISCCTUSER_in[8] = (SAXISCCTUSER[8] === 1'bz) || SAXISCCTUSER_delay[8]; // rv 1
  assign SAXISCCTUSER_in[9] = (SAXISCCTUSER[9] === 1'bz) || SAXISCCTUSER_delay[9]; // rv 1
  assign SAXISCCTVALID_in = (SAXISCCTVALID !== 1'bz) && SAXISCCTVALID_delay; // rv 0
  assign SAXISRQTDATA_in[0] = (SAXISRQTDATA[0] === 1'bz) || SAXISRQTDATA_delay[0]; // rv 1
  assign SAXISRQTDATA_in[100] = (SAXISRQTDATA[100] === 1'bz) || SAXISRQTDATA_delay[100]; // rv 1
  assign SAXISRQTDATA_in[101] = (SAXISRQTDATA[101] === 1'bz) || SAXISRQTDATA_delay[101]; // rv 1
  assign SAXISRQTDATA_in[102] = (SAXISRQTDATA[102] === 1'bz) || SAXISRQTDATA_delay[102]; // rv 1
  assign SAXISRQTDATA_in[103] = (SAXISRQTDATA[103] === 1'bz) || SAXISRQTDATA_delay[103]; // rv 1
  assign SAXISRQTDATA_in[104] = (SAXISRQTDATA[104] === 1'bz) || SAXISRQTDATA_delay[104]; // rv 1
  assign SAXISRQTDATA_in[105] = (SAXISRQTDATA[105] === 1'bz) || SAXISRQTDATA_delay[105]; // rv 1
  assign SAXISRQTDATA_in[106] = (SAXISRQTDATA[106] === 1'bz) || SAXISRQTDATA_delay[106]; // rv 1
  assign SAXISRQTDATA_in[107] = (SAXISRQTDATA[107] === 1'bz) || SAXISRQTDATA_delay[107]; // rv 1
  assign SAXISRQTDATA_in[108] = (SAXISRQTDATA[108] === 1'bz) || SAXISRQTDATA_delay[108]; // rv 1
  assign SAXISRQTDATA_in[109] = (SAXISRQTDATA[109] === 1'bz) || SAXISRQTDATA_delay[109]; // rv 1
  assign SAXISRQTDATA_in[10] = (SAXISRQTDATA[10] === 1'bz) || SAXISRQTDATA_delay[10]; // rv 1
  assign SAXISRQTDATA_in[110] = (SAXISRQTDATA[110] === 1'bz) || SAXISRQTDATA_delay[110]; // rv 1
  assign SAXISRQTDATA_in[111] = (SAXISRQTDATA[111] === 1'bz) || SAXISRQTDATA_delay[111]; // rv 1
  assign SAXISRQTDATA_in[112] = (SAXISRQTDATA[112] === 1'bz) || SAXISRQTDATA_delay[112]; // rv 1
  assign SAXISRQTDATA_in[113] = (SAXISRQTDATA[113] === 1'bz) || SAXISRQTDATA_delay[113]; // rv 1
  assign SAXISRQTDATA_in[114] = (SAXISRQTDATA[114] === 1'bz) || SAXISRQTDATA_delay[114]; // rv 1
  assign SAXISRQTDATA_in[115] = (SAXISRQTDATA[115] === 1'bz) || SAXISRQTDATA_delay[115]; // rv 1
  assign SAXISRQTDATA_in[116] = (SAXISRQTDATA[116] === 1'bz) || SAXISRQTDATA_delay[116]; // rv 1
  assign SAXISRQTDATA_in[117] = (SAXISRQTDATA[117] === 1'bz) || SAXISRQTDATA_delay[117]; // rv 1
  assign SAXISRQTDATA_in[118] = (SAXISRQTDATA[118] === 1'bz) || SAXISRQTDATA_delay[118]; // rv 1
  assign SAXISRQTDATA_in[119] = (SAXISRQTDATA[119] === 1'bz) || SAXISRQTDATA_delay[119]; // rv 1
  assign SAXISRQTDATA_in[11] = (SAXISRQTDATA[11] === 1'bz) || SAXISRQTDATA_delay[11]; // rv 1
  assign SAXISRQTDATA_in[120] = (SAXISRQTDATA[120] === 1'bz) || SAXISRQTDATA_delay[120]; // rv 1
  assign SAXISRQTDATA_in[121] = (SAXISRQTDATA[121] === 1'bz) || SAXISRQTDATA_delay[121]; // rv 1
  assign SAXISRQTDATA_in[122] = (SAXISRQTDATA[122] === 1'bz) || SAXISRQTDATA_delay[122]; // rv 1
  assign SAXISRQTDATA_in[123] = (SAXISRQTDATA[123] === 1'bz) || SAXISRQTDATA_delay[123]; // rv 1
  assign SAXISRQTDATA_in[124] = (SAXISRQTDATA[124] === 1'bz) || SAXISRQTDATA_delay[124]; // rv 1
  assign SAXISRQTDATA_in[125] = (SAXISRQTDATA[125] === 1'bz) || SAXISRQTDATA_delay[125]; // rv 1
  assign SAXISRQTDATA_in[126] = (SAXISRQTDATA[126] === 1'bz) || SAXISRQTDATA_delay[126]; // rv 1
  assign SAXISRQTDATA_in[127] = (SAXISRQTDATA[127] === 1'bz) || SAXISRQTDATA_delay[127]; // rv 1
  assign SAXISRQTDATA_in[128] = (SAXISRQTDATA[128] === 1'bz) || SAXISRQTDATA_delay[128]; // rv 1
  assign SAXISRQTDATA_in[129] = (SAXISRQTDATA[129] === 1'bz) || SAXISRQTDATA_delay[129]; // rv 1
  assign SAXISRQTDATA_in[12] = (SAXISRQTDATA[12] === 1'bz) || SAXISRQTDATA_delay[12]; // rv 1
  assign SAXISRQTDATA_in[130] = (SAXISRQTDATA[130] === 1'bz) || SAXISRQTDATA_delay[130]; // rv 1
  assign SAXISRQTDATA_in[131] = (SAXISRQTDATA[131] === 1'bz) || SAXISRQTDATA_delay[131]; // rv 1
  assign SAXISRQTDATA_in[132] = (SAXISRQTDATA[132] === 1'bz) || SAXISRQTDATA_delay[132]; // rv 1
  assign SAXISRQTDATA_in[133] = (SAXISRQTDATA[133] === 1'bz) || SAXISRQTDATA_delay[133]; // rv 1
  assign SAXISRQTDATA_in[134] = (SAXISRQTDATA[134] === 1'bz) || SAXISRQTDATA_delay[134]; // rv 1
  assign SAXISRQTDATA_in[135] = (SAXISRQTDATA[135] === 1'bz) || SAXISRQTDATA_delay[135]; // rv 1
  assign SAXISRQTDATA_in[136] = (SAXISRQTDATA[136] === 1'bz) || SAXISRQTDATA_delay[136]; // rv 1
  assign SAXISRQTDATA_in[137] = (SAXISRQTDATA[137] === 1'bz) || SAXISRQTDATA_delay[137]; // rv 1
  assign SAXISRQTDATA_in[138] = (SAXISRQTDATA[138] === 1'bz) || SAXISRQTDATA_delay[138]; // rv 1
  assign SAXISRQTDATA_in[139] = (SAXISRQTDATA[139] === 1'bz) || SAXISRQTDATA_delay[139]; // rv 1
  assign SAXISRQTDATA_in[13] = (SAXISRQTDATA[13] === 1'bz) || SAXISRQTDATA_delay[13]; // rv 1
  assign SAXISRQTDATA_in[140] = (SAXISRQTDATA[140] === 1'bz) || SAXISRQTDATA_delay[140]; // rv 1
  assign SAXISRQTDATA_in[141] = (SAXISRQTDATA[141] === 1'bz) || SAXISRQTDATA_delay[141]; // rv 1
  assign SAXISRQTDATA_in[142] = (SAXISRQTDATA[142] === 1'bz) || SAXISRQTDATA_delay[142]; // rv 1
  assign SAXISRQTDATA_in[143] = (SAXISRQTDATA[143] === 1'bz) || SAXISRQTDATA_delay[143]; // rv 1
  assign SAXISRQTDATA_in[144] = (SAXISRQTDATA[144] === 1'bz) || SAXISRQTDATA_delay[144]; // rv 1
  assign SAXISRQTDATA_in[145] = (SAXISRQTDATA[145] === 1'bz) || SAXISRQTDATA_delay[145]; // rv 1
  assign SAXISRQTDATA_in[146] = (SAXISRQTDATA[146] === 1'bz) || SAXISRQTDATA_delay[146]; // rv 1
  assign SAXISRQTDATA_in[147] = (SAXISRQTDATA[147] === 1'bz) || SAXISRQTDATA_delay[147]; // rv 1
  assign SAXISRQTDATA_in[148] = (SAXISRQTDATA[148] === 1'bz) || SAXISRQTDATA_delay[148]; // rv 1
  assign SAXISRQTDATA_in[149] = (SAXISRQTDATA[149] === 1'bz) || SAXISRQTDATA_delay[149]; // rv 1
  assign SAXISRQTDATA_in[14] = (SAXISRQTDATA[14] === 1'bz) || SAXISRQTDATA_delay[14]; // rv 1
  assign SAXISRQTDATA_in[150] = (SAXISRQTDATA[150] === 1'bz) || SAXISRQTDATA_delay[150]; // rv 1
  assign SAXISRQTDATA_in[151] = (SAXISRQTDATA[151] === 1'bz) || SAXISRQTDATA_delay[151]; // rv 1
  assign SAXISRQTDATA_in[152] = (SAXISRQTDATA[152] === 1'bz) || SAXISRQTDATA_delay[152]; // rv 1
  assign SAXISRQTDATA_in[153] = (SAXISRQTDATA[153] === 1'bz) || SAXISRQTDATA_delay[153]; // rv 1
  assign SAXISRQTDATA_in[154] = (SAXISRQTDATA[154] === 1'bz) || SAXISRQTDATA_delay[154]; // rv 1
  assign SAXISRQTDATA_in[155] = (SAXISRQTDATA[155] === 1'bz) || SAXISRQTDATA_delay[155]; // rv 1
  assign SAXISRQTDATA_in[156] = (SAXISRQTDATA[156] === 1'bz) || SAXISRQTDATA_delay[156]; // rv 1
  assign SAXISRQTDATA_in[157] = (SAXISRQTDATA[157] === 1'bz) || SAXISRQTDATA_delay[157]; // rv 1
  assign SAXISRQTDATA_in[158] = (SAXISRQTDATA[158] === 1'bz) || SAXISRQTDATA_delay[158]; // rv 1
  assign SAXISRQTDATA_in[159] = (SAXISRQTDATA[159] === 1'bz) || SAXISRQTDATA_delay[159]; // rv 1
  assign SAXISRQTDATA_in[15] = (SAXISRQTDATA[15] === 1'bz) || SAXISRQTDATA_delay[15]; // rv 1
  assign SAXISRQTDATA_in[160] = (SAXISRQTDATA[160] === 1'bz) || SAXISRQTDATA_delay[160]; // rv 1
  assign SAXISRQTDATA_in[161] = (SAXISRQTDATA[161] === 1'bz) || SAXISRQTDATA_delay[161]; // rv 1
  assign SAXISRQTDATA_in[162] = (SAXISRQTDATA[162] === 1'bz) || SAXISRQTDATA_delay[162]; // rv 1
  assign SAXISRQTDATA_in[163] = (SAXISRQTDATA[163] === 1'bz) || SAXISRQTDATA_delay[163]; // rv 1
  assign SAXISRQTDATA_in[164] = (SAXISRQTDATA[164] === 1'bz) || SAXISRQTDATA_delay[164]; // rv 1
  assign SAXISRQTDATA_in[165] = (SAXISRQTDATA[165] === 1'bz) || SAXISRQTDATA_delay[165]; // rv 1
  assign SAXISRQTDATA_in[166] = (SAXISRQTDATA[166] === 1'bz) || SAXISRQTDATA_delay[166]; // rv 1
  assign SAXISRQTDATA_in[167] = (SAXISRQTDATA[167] === 1'bz) || SAXISRQTDATA_delay[167]; // rv 1
  assign SAXISRQTDATA_in[168] = (SAXISRQTDATA[168] === 1'bz) || SAXISRQTDATA_delay[168]; // rv 1
  assign SAXISRQTDATA_in[169] = (SAXISRQTDATA[169] === 1'bz) || SAXISRQTDATA_delay[169]; // rv 1
  assign SAXISRQTDATA_in[16] = (SAXISRQTDATA[16] === 1'bz) || SAXISRQTDATA_delay[16]; // rv 1
  assign SAXISRQTDATA_in[170] = (SAXISRQTDATA[170] === 1'bz) || SAXISRQTDATA_delay[170]; // rv 1
  assign SAXISRQTDATA_in[171] = (SAXISRQTDATA[171] === 1'bz) || SAXISRQTDATA_delay[171]; // rv 1
  assign SAXISRQTDATA_in[172] = (SAXISRQTDATA[172] === 1'bz) || SAXISRQTDATA_delay[172]; // rv 1
  assign SAXISRQTDATA_in[173] = (SAXISRQTDATA[173] === 1'bz) || SAXISRQTDATA_delay[173]; // rv 1
  assign SAXISRQTDATA_in[174] = (SAXISRQTDATA[174] === 1'bz) || SAXISRQTDATA_delay[174]; // rv 1
  assign SAXISRQTDATA_in[175] = (SAXISRQTDATA[175] === 1'bz) || SAXISRQTDATA_delay[175]; // rv 1
  assign SAXISRQTDATA_in[176] = (SAXISRQTDATA[176] === 1'bz) || SAXISRQTDATA_delay[176]; // rv 1
  assign SAXISRQTDATA_in[177] = (SAXISRQTDATA[177] === 1'bz) || SAXISRQTDATA_delay[177]; // rv 1
  assign SAXISRQTDATA_in[178] = (SAXISRQTDATA[178] === 1'bz) || SAXISRQTDATA_delay[178]; // rv 1
  assign SAXISRQTDATA_in[179] = (SAXISRQTDATA[179] === 1'bz) || SAXISRQTDATA_delay[179]; // rv 1
  assign SAXISRQTDATA_in[17] = (SAXISRQTDATA[17] === 1'bz) || SAXISRQTDATA_delay[17]; // rv 1
  assign SAXISRQTDATA_in[180] = (SAXISRQTDATA[180] === 1'bz) || SAXISRQTDATA_delay[180]; // rv 1
  assign SAXISRQTDATA_in[181] = (SAXISRQTDATA[181] === 1'bz) || SAXISRQTDATA_delay[181]; // rv 1
  assign SAXISRQTDATA_in[182] = (SAXISRQTDATA[182] === 1'bz) || SAXISRQTDATA_delay[182]; // rv 1
  assign SAXISRQTDATA_in[183] = (SAXISRQTDATA[183] === 1'bz) || SAXISRQTDATA_delay[183]; // rv 1
  assign SAXISRQTDATA_in[184] = (SAXISRQTDATA[184] === 1'bz) || SAXISRQTDATA_delay[184]; // rv 1
  assign SAXISRQTDATA_in[185] = (SAXISRQTDATA[185] === 1'bz) || SAXISRQTDATA_delay[185]; // rv 1
  assign SAXISRQTDATA_in[186] = (SAXISRQTDATA[186] === 1'bz) || SAXISRQTDATA_delay[186]; // rv 1
  assign SAXISRQTDATA_in[187] = (SAXISRQTDATA[187] === 1'bz) || SAXISRQTDATA_delay[187]; // rv 1
  assign SAXISRQTDATA_in[188] = (SAXISRQTDATA[188] === 1'bz) || SAXISRQTDATA_delay[188]; // rv 1
  assign SAXISRQTDATA_in[189] = (SAXISRQTDATA[189] === 1'bz) || SAXISRQTDATA_delay[189]; // rv 1
  assign SAXISRQTDATA_in[18] = (SAXISRQTDATA[18] === 1'bz) || SAXISRQTDATA_delay[18]; // rv 1
  assign SAXISRQTDATA_in[190] = (SAXISRQTDATA[190] === 1'bz) || SAXISRQTDATA_delay[190]; // rv 1
  assign SAXISRQTDATA_in[191] = (SAXISRQTDATA[191] === 1'bz) || SAXISRQTDATA_delay[191]; // rv 1
  assign SAXISRQTDATA_in[192] = (SAXISRQTDATA[192] === 1'bz) || SAXISRQTDATA_delay[192]; // rv 1
  assign SAXISRQTDATA_in[193] = (SAXISRQTDATA[193] === 1'bz) || SAXISRQTDATA_delay[193]; // rv 1
  assign SAXISRQTDATA_in[194] = (SAXISRQTDATA[194] === 1'bz) || SAXISRQTDATA_delay[194]; // rv 1
  assign SAXISRQTDATA_in[195] = (SAXISRQTDATA[195] === 1'bz) || SAXISRQTDATA_delay[195]; // rv 1
  assign SAXISRQTDATA_in[196] = (SAXISRQTDATA[196] === 1'bz) || SAXISRQTDATA_delay[196]; // rv 1
  assign SAXISRQTDATA_in[197] = (SAXISRQTDATA[197] === 1'bz) || SAXISRQTDATA_delay[197]; // rv 1
  assign SAXISRQTDATA_in[198] = (SAXISRQTDATA[198] === 1'bz) || SAXISRQTDATA_delay[198]; // rv 1
  assign SAXISRQTDATA_in[199] = (SAXISRQTDATA[199] === 1'bz) || SAXISRQTDATA_delay[199]; // rv 1
  assign SAXISRQTDATA_in[19] = (SAXISRQTDATA[19] === 1'bz) || SAXISRQTDATA_delay[19]; // rv 1
  assign SAXISRQTDATA_in[1] = (SAXISRQTDATA[1] === 1'bz) || SAXISRQTDATA_delay[1]; // rv 1
  assign SAXISRQTDATA_in[200] = (SAXISRQTDATA[200] === 1'bz) || SAXISRQTDATA_delay[200]; // rv 1
  assign SAXISRQTDATA_in[201] = (SAXISRQTDATA[201] === 1'bz) || SAXISRQTDATA_delay[201]; // rv 1
  assign SAXISRQTDATA_in[202] = (SAXISRQTDATA[202] === 1'bz) || SAXISRQTDATA_delay[202]; // rv 1
  assign SAXISRQTDATA_in[203] = (SAXISRQTDATA[203] === 1'bz) || SAXISRQTDATA_delay[203]; // rv 1
  assign SAXISRQTDATA_in[204] = (SAXISRQTDATA[204] === 1'bz) || SAXISRQTDATA_delay[204]; // rv 1
  assign SAXISRQTDATA_in[205] = (SAXISRQTDATA[205] === 1'bz) || SAXISRQTDATA_delay[205]; // rv 1
  assign SAXISRQTDATA_in[206] = (SAXISRQTDATA[206] === 1'bz) || SAXISRQTDATA_delay[206]; // rv 1
  assign SAXISRQTDATA_in[207] = (SAXISRQTDATA[207] === 1'bz) || SAXISRQTDATA_delay[207]; // rv 1
  assign SAXISRQTDATA_in[208] = (SAXISRQTDATA[208] === 1'bz) || SAXISRQTDATA_delay[208]; // rv 1
  assign SAXISRQTDATA_in[209] = (SAXISRQTDATA[209] === 1'bz) || SAXISRQTDATA_delay[209]; // rv 1
  assign SAXISRQTDATA_in[20] = (SAXISRQTDATA[20] === 1'bz) || SAXISRQTDATA_delay[20]; // rv 1
  assign SAXISRQTDATA_in[210] = (SAXISRQTDATA[210] === 1'bz) || SAXISRQTDATA_delay[210]; // rv 1
  assign SAXISRQTDATA_in[211] = (SAXISRQTDATA[211] === 1'bz) || SAXISRQTDATA_delay[211]; // rv 1
  assign SAXISRQTDATA_in[212] = (SAXISRQTDATA[212] === 1'bz) || SAXISRQTDATA_delay[212]; // rv 1
  assign SAXISRQTDATA_in[213] = (SAXISRQTDATA[213] === 1'bz) || SAXISRQTDATA_delay[213]; // rv 1
  assign SAXISRQTDATA_in[214] = (SAXISRQTDATA[214] === 1'bz) || SAXISRQTDATA_delay[214]; // rv 1
  assign SAXISRQTDATA_in[215] = (SAXISRQTDATA[215] === 1'bz) || SAXISRQTDATA_delay[215]; // rv 1
  assign SAXISRQTDATA_in[216] = (SAXISRQTDATA[216] === 1'bz) || SAXISRQTDATA_delay[216]; // rv 1
  assign SAXISRQTDATA_in[217] = (SAXISRQTDATA[217] === 1'bz) || SAXISRQTDATA_delay[217]; // rv 1
  assign SAXISRQTDATA_in[218] = (SAXISRQTDATA[218] === 1'bz) || SAXISRQTDATA_delay[218]; // rv 1
  assign SAXISRQTDATA_in[219] = (SAXISRQTDATA[219] === 1'bz) || SAXISRQTDATA_delay[219]; // rv 1
  assign SAXISRQTDATA_in[21] = (SAXISRQTDATA[21] === 1'bz) || SAXISRQTDATA_delay[21]; // rv 1
  assign SAXISRQTDATA_in[220] = (SAXISRQTDATA[220] === 1'bz) || SAXISRQTDATA_delay[220]; // rv 1
  assign SAXISRQTDATA_in[221] = (SAXISRQTDATA[221] === 1'bz) || SAXISRQTDATA_delay[221]; // rv 1
  assign SAXISRQTDATA_in[222] = (SAXISRQTDATA[222] === 1'bz) || SAXISRQTDATA_delay[222]; // rv 1
  assign SAXISRQTDATA_in[223] = (SAXISRQTDATA[223] === 1'bz) || SAXISRQTDATA_delay[223]; // rv 1
  assign SAXISRQTDATA_in[224] = (SAXISRQTDATA[224] === 1'bz) || SAXISRQTDATA_delay[224]; // rv 1
  assign SAXISRQTDATA_in[225] = (SAXISRQTDATA[225] === 1'bz) || SAXISRQTDATA_delay[225]; // rv 1
  assign SAXISRQTDATA_in[226] = (SAXISRQTDATA[226] === 1'bz) || SAXISRQTDATA_delay[226]; // rv 1
  assign SAXISRQTDATA_in[227] = (SAXISRQTDATA[227] === 1'bz) || SAXISRQTDATA_delay[227]; // rv 1
  assign SAXISRQTDATA_in[228] = (SAXISRQTDATA[228] === 1'bz) || SAXISRQTDATA_delay[228]; // rv 1
  assign SAXISRQTDATA_in[229] = (SAXISRQTDATA[229] === 1'bz) || SAXISRQTDATA_delay[229]; // rv 1
  assign SAXISRQTDATA_in[22] = (SAXISRQTDATA[22] === 1'bz) || SAXISRQTDATA_delay[22]; // rv 1
  assign SAXISRQTDATA_in[230] = (SAXISRQTDATA[230] === 1'bz) || SAXISRQTDATA_delay[230]; // rv 1
  assign SAXISRQTDATA_in[231] = (SAXISRQTDATA[231] === 1'bz) || SAXISRQTDATA_delay[231]; // rv 1
  assign SAXISRQTDATA_in[232] = (SAXISRQTDATA[232] === 1'bz) || SAXISRQTDATA_delay[232]; // rv 1
  assign SAXISRQTDATA_in[233] = (SAXISRQTDATA[233] === 1'bz) || SAXISRQTDATA_delay[233]; // rv 1
  assign SAXISRQTDATA_in[234] = (SAXISRQTDATA[234] === 1'bz) || SAXISRQTDATA_delay[234]; // rv 1
  assign SAXISRQTDATA_in[235] = (SAXISRQTDATA[235] === 1'bz) || SAXISRQTDATA_delay[235]; // rv 1
  assign SAXISRQTDATA_in[236] = (SAXISRQTDATA[236] === 1'bz) || SAXISRQTDATA_delay[236]; // rv 1
  assign SAXISRQTDATA_in[237] = (SAXISRQTDATA[237] === 1'bz) || SAXISRQTDATA_delay[237]; // rv 1
  assign SAXISRQTDATA_in[238] = (SAXISRQTDATA[238] === 1'bz) || SAXISRQTDATA_delay[238]; // rv 1
  assign SAXISRQTDATA_in[239] = (SAXISRQTDATA[239] === 1'bz) || SAXISRQTDATA_delay[239]; // rv 1
  assign SAXISRQTDATA_in[23] = (SAXISRQTDATA[23] === 1'bz) || SAXISRQTDATA_delay[23]; // rv 1
  assign SAXISRQTDATA_in[240] = (SAXISRQTDATA[240] === 1'bz) || SAXISRQTDATA_delay[240]; // rv 1
  assign SAXISRQTDATA_in[241] = (SAXISRQTDATA[241] === 1'bz) || SAXISRQTDATA_delay[241]; // rv 1
  assign SAXISRQTDATA_in[242] = (SAXISRQTDATA[242] === 1'bz) || SAXISRQTDATA_delay[242]; // rv 1
  assign SAXISRQTDATA_in[243] = (SAXISRQTDATA[243] === 1'bz) || SAXISRQTDATA_delay[243]; // rv 1
  assign SAXISRQTDATA_in[244] = (SAXISRQTDATA[244] === 1'bz) || SAXISRQTDATA_delay[244]; // rv 1
  assign SAXISRQTDATA_in[245] = (SAXISRQTDATA[245] === 1'bz) || SAXISRQTDATA_delay[245]; // rv 1
  assign SAXISRQTDATA_in[246] = (SAXISRQTDATA[246] === 1'bz) || SAXISRQTDATA_delay[246]; // rv 1
  assign SAXISRQTDATA_in[247] = (SAXISRQTDATA[247] === 1'bz) || SAXISRQTDATA_delay[247]; // rv 1
  assign SAXISRQTDATA_in[248] = (SAXISRQTDATA[248] === 1'bz) || SAXISRQTDATA_delay[248]; // rv 1
  assign SAXISRQTDATA_in[249] = (SAXISRQTDATA[249] === 1'bz) || SAXISRQTDATA_delay[249]; // rv 1
  assign SAXISRQTDATA_in[24] = (SAXISRQTDATA[24] === 1'bz) || SAXISRQTDATA_delay[24]; // rv 1
  assign SAXISRQTDATA_in[250] = (SAXISRQTDATA[250] === 1'bz) || SAXISRQTDATA_delay[250]; // rv 1
  assign SAXISRQTDATA_in[251] = (SAXISRQTDATA[251] === 1'bz) || SAXISRQTDATA_delay[251]; // rv 1
  assign SAXISRQTDATA_in[252] = (SAXISRQTDATA[252] === 1'bz) || SAXISRQTDATA_delay[252]; // rv 1
  assign SAXISRQTDATA_in[253] = (SAXISRQTDATA[253] === 1'bz) || SAXISRQTDATA_delay[253]; // rv 1
  assign SAXISRQTDATA_in[254] = (SAXISRQTDATA[254] === 1'bz) || SAXISRQTDATA_delay[254]; // rv 1
  assign SAXISRQTDATA_in[255] = (SAXISRQTDATA[255] === 1'bz) || SAXISRQTDATA_delay[255]; // rv 1
  assign SAXISRQTDATA_in[25] = (SAXISRQTDATA[25] === 1'bz) || SAXISRQTDATA_delay[25]; // rv 1
  assign SAXISRQTDATA_in[26] = (SAXISRQTDATA[26] === 1'bz) || SAXISRQTDATA_delay[26]; // rv 1
  assign SAXISRQTDATA_in[27] = (SAXISRQTDATA[27] === 1'bz) || SAXISRQTDATA_delay[27]; // rv 1
  assign SAXISRQTDATA_in[28] = (SAXISRQTDATA[28] === 1'bz) || SAXISRQTDATA_delay[28]; // rv 1
  assign SAXISRQTDATA_in[29] = (SAXISRQTDATA[29] === 1'bz) || SAXISRQTDATA_delay[29]; // rv 1
  assign SAXISRQTDATA_in[2] = (SAXISRQTDATA[2] === 1'bz) || SAXISRQTDATA_delay[2]; // rv 1
  assign SAXISRQTDATA_in[30] = (SAXISRQTDATA[30] === 1'bz) || SAXISRQTDATA_delay[30]; // rv 1
  assign SAXISRQTDATA_in[31] = (SAXISRQTDATA[31] === 1'bz) || SAXISRQTDATA_delay[31]; // rv 1
  assign SAXISRQTDATA_in[32] = (SAXISRQTDATA[32] === 1'bz) || SAXISRQTDATA_delay[32]; // rv 1
  assign SAXISRQTDATA_in[33] = (SAXISRQTDATA[33] === 1'bz) || SAXISRQTDATA_delay[33]; // rv 1
  assign SAXISRQTDATA_in[34] = (SAXISRQTDATA[34] === 1'bz) || SAXISRQTDATA_delay[34]; // rv 1
  assign SAXISRQTDATA_in[35] = (SAXISRQTDATA[35] === 1'bz) || SAXISRQTDATA_delay[35]; // rv 1
  assign SAXISRQTDATA_in[36] = (SAXISRQTDATA[36] === 1'bz) || SAXISRQTDATA_delay[36]; // rv 1
  assign SAXISRQTDATA_in[37] = (SAXISRQTDATA[37] === 1'bz) || SAXISRQTDATA_delay[37]; // rv 1
  assign SAXISRQTDATA_in[38] = (SAXISRQTDATA[38] === 1'bz) || SAXISRQTDATA_delay[38]; // rv 1
  assign SAXISRQTDATA_in[39] = (SAXISRQTDATA[39] === 1'bz) || SAXISRQTDATA_delay[39]; // rv 1
  assign SAXISRQTDATA_in[3] = (SAXISRQTDATA[3] === 1'bz) || SAXISRQTDATA_delay[3]; // rv 1
  assign SAXISRQTDATA_in[40] = (SAXISRQTDATA[40] === 1'bz) || SAXISRQTDATA_delay[40]; // rv 1
  assign SAXISRQTDATA_in[41] = (SAXISRQTDATA[41] === 1'bz) || SAXISRQTDATA_delay[41]; // rv 1
  assign SAXISRQTDATA_in[42] = (SAXISRQTDATA[42] === 1'bz) || SAXISRQTDATA_delay[42]; // rv 1
  assign SAXISRQTDATA_in[43] = (SAXISRQTDATA[43] === 1'bz) || SAXISRQTDATA_delay[43]; // rv 1
  assign SAXISRQTDATA_in[44] = (SAXISRQTDATA[44] === 1'bz) || SAXISRQTDATA_delay[44]; // rv 1
  assign SAXISRQTDATA_in[45] = (SAXISRQTDATA[45] === 1'bz) || SAXISRQTDATA_delay[45]; // rv 1
  assign SAXISRQTDATA_in[46] = (SAXISRQTDATA[46] === 1'bz) || SAXISRQTDATA_delay[46]; // rv 1
  assign SAXISRQTDATA_in[47] = (SAXISRQTDATA[47] === 1'bz) || SAXISRQTDATA_delay[47]; // rv 1
  assign SAXISRQTDATA_in[48] = (SAXISRQTDATA[48] === 1'bz) || SAXISRQTDATA_delay[48]; // rv 1
  assign SAXISRQTDATA_in[49] = (SAXISRQTDATA[49] === 1'bz) || SAXISRQTDATA_delay[49]; // rv 1
  assign SAXISRQTDATA_in[4] = (SAXISRQTDATA[4] === 1'bz) || SAXISRQTDATA_delay[4]; // rv 1
  assign SAXISRQTDATA_in[50] = (SAXISRQTDATA[50] === 1'bz) || SAXISRQTDATA_delay[50]; // rv 1
  assign SAXISRQTDATA_in[51] = (SAXISRQTDATA[51] === 1'bz) || SAXISRQTDATA_delay[51]; // rv 1
  assign SAXISRQTDATA_in[52] = (SAXISRQTDATA[52] === 1'bz) || SAXISRQTDATA_delay[52]; // rv 1
  assign SAXISRQTDATA_in[53] = (SAXISRQTDATA[53] === 1'bz) || SAXISRQTDATA_delay[53]; // rv 1
  assign SAXISRQTDATA_in[54] = (SAXISRQTDATA[54] === 1'bz) || SAXISRQTDATA_delay[54]; // rv 1
  assign SAXISRQTDATA_in[55] = (SAXISRQTDATA[55] === 1'bz) || SAXISRQTDATA_delay[55]; // rv 1
  assign SAXISRQTDATA_in[56] = (SAXISRQTDATA[56] === 1'bz) || SAXISRQTDATA_delay[56]; // rv 1
  assign SAXISRQTDATA_in[57] = (SAXISRQTDATA[57] === 1'bz) || SAXISRQTDATA_delay[57]; // rv 1
  assign SAXISRQTDATA_in[58] = (SAXISRQTDATA[58] === 1'bz) || SAXISRQTDATA_delay[58]; // rv 1
  assign SAXISRQTDATA_in[59] = (SAXISRQTDATA[59] === 1'bz) || SAXISRQTDATA_delay[59]; // rv 1
  assign SAXISRQTDATA_in[5] = (SAXISRQTDATA[5] === 1'bz) || SAXISRQTDATA_delay[5]; // rv 1
  assign SAXISRQTDATA_in[60] = (SAXISRQTDATA[60] === 1'bz) || SAXISRQTDATA_delay[60]; // rv 1
  assign SAXISRQTDATA_in[61] = (SAXISRQTDATA[61] === 1'bz) || SAXISRQTDATA_delay[61]; // rv 1
  assign SAXISRQTDATA_in[62] = (SAXISRQTDATA[62] === 1'bz) || SAXISRQTDATA_delay[62]; // rv 1
  assign SAXISRQTDATA_in[63] = (SAXISRQTDATA[63] === 1'bz) || SAXISRQTDATA_delay[63]; // rv 1
  assign SAXISRQTDATA_in[64] = (SAXISRQTDATA[64] === 1'bz) || SAXISRQTDATA_delay[64]; // rv 1
  assign SAXISRQTDATA_in[65] = (SAXISRQTDATA[65] === 1'bz) || SAXISRQTDATA_delay[65]; // rv 1
  assign SAXISRQTDATA_in[66] = (SAXISRQTDATA[66] === 1'bz) || SAXISRQTDATA_delay[66]; // rv 1
  assign SAXISRQTDATA_in[67] = (SAXISRQTDATA[67] === 1'bz) || SAXISRQTDATA_delay[67]; // rv 1
  assign SAXISRQTDATA_in[68] = (SAXISRQTDATA[68] === 1'bz) || SAXISRQTDATA_delay[68]; // rv 1
  assign SAXISRQTDATA_in[69] = (SAXISRQTDATA[69] === 1'bz) || SAXISRQTDATA_delay[69]; // rv 1
  assign SAXISRQTDATA_in[6] = (SAXISRQTDATA[6] === 1'bz) || SAXISRQTDATA_delay[6]; // rv 1
  assign SAXISRQTDATA_in[70] = (SAXISRQTDATA[70] === 1'bz) || SAXISRQTDATA_delay[70]; // rv 1
  assign SAXISRQTDATA_in[71] = (SAXISRQTDATA[71] === 1'bz) || SAXISRQTDATA_delay[71]; // rv 1
  assign SAXISRQTDATA_in[72] = (SAXISRQTDATA[72] === 1'bz) || SAXISRQTDATA_delay[72]; // rv 1
  assign SAXISRQTDATA_in[73] = (SAXISRQTDATA[73] === 1'bz) || SAXISRQTDATA_delay[73]; // rv 1
  assign SAXISRQTDATA_in[74] = (SAXISRQTDATA[74] === 1'bz) || SAXISRQTDATA_delay[74]; // rv 1
  assign SAXISRQTDATA_in[75] = (SAXISRQTDATA[75] === 1'bz) || SAXISRQTDATA_delay[75]; // rv 1
  assign SAXISRQTDATA_in[76] = (SAXISRQTDATA[76] === 1'bz) || SAXISRQTDATA_delay[76]; // rv 1
  assign SAXISRQTDATA_in[77] = (SAXISRQTDATA[77] === 1'bz) || SAXISRQTDATA_delay[77]; // rv 1
  assign SAXISRQTDATA_in[78] = (SAXISRQTDATA[78] === 1'bz) || SAXISRQTDATA_delay[78]; // rv 1
  assign SAXISRQTDATA_in[79] = (SAXISRQTDATA[79] === 1'bz) || SAXISRQTDATA_delay[79]; // rv 1
  assign SAXISRQTDATA_in[7] = (SAXISRQTDATA[7] === 1'bz) || SAXISRQTDATA_delay[7]; // rv 1
  assign SAXISRQTDATA_in[80] = (SAXISRQTDATA[80] === 1'bz) || SAXISRQTDATA_delay[80]; // rv 1
  assign SAXISRQTDATA_in[81] = (SAXISRQTDATA[81] === 1'bz) || SAXISRQTDATA_delay[81]; // rv 1
  assign SAXISRQTDATA_in[82] = (SAXISRQTDATA[82] === 1'bz) || SAXISRQTDATA_delay[82]; // rv 1
  assign SAXISRQTDATA_in[83] = (SAXISRQTDATA[83] === 1'bz) || SAXISRQTDATA_delay[83]; // rv 1
  assign SAXISRQTDATA_in[84] = (SAXISRQTDATA[84] === 1'bz) || SAXISRQTDATA_delay[84]; // rv 1
  assign SAXISRQTDATA_in[85] = (SAXISRQTDATA[85] === 1'bz) || SAXISRQTDATA_delay[85]; // rv 1
  assign SAXISRQTDATA_in[86] = (SAXISRQTDATA[86] === 1'bz) || SAXISRQTDATA_delay[86]; // rv 1
  assign SAXISRQTDATA_in[87] = (SAXISRQTDATA[87] === 1'bz) || SAXISRQTDATA_delay[87]; // rv 1
  assign SAXISRQTDATA_in[88] = (SAXISRQTDATA[88] === 1'bz) || SAXISRQTDATA_delay[88]; // rv 1
  assign SAXISRQTDATA_in[89] = (SAXISRQTDATA[89] === 1'bz) || SAXISRQTDATA_delay[89]; // rv 1
  assign SAXISRQTDATA_in[8] = (SAXISRQTDATA[8] === 1'bz) || SAXISRQTDATA_delay[8]; // rv 1
  assign SAXISRQTDATA_in[90] = (SAXISRQTDATA[90] === 1'bz) || SAXISRQTDATA_delay[90]; // rv 1
  assign SAXISRQTDATA_in[91] = (SAXISRQTDATA[91] === 1'bz) || SAXISRQTDATA_delay[91]; // rv 1
  assign SAXISRQTDATA_in[92] = (SAXISRQTDATA[92] === 1'bz) || SAXISRQTDATA_delay[92]; // rv 1
  assign SAXISRQTDATA_in[93] = (SAXISRQTDATA[93] === 1'bz) || SAXISRQTDATA_delay[93]; // rv 1
  assign SAXISRQTDATA_in[94] = (SAXISRQTDATA[94] === 1'bz) || SAXISRQTDATA_delay[94]; // rv 1
  assign SAXISRQTDATA_in[95] = (SAXISRQTDATA[95] === 1'bz) || SAXISRQTDATA_delay[95]; // rv 1
  assign SAXISRQTDATA_in[96] = (SAXISRQTDATA[96] === 1'bz) || SAXISRQTDATA_delay[96]; // rv 1
  assign SAXISRQTDATA_in[97] = (SAXISRQTDATA[97] === 1'bz) || SAXISRQTDATA_delay[97]; // rv 1
  assign SAXISRQTDATA_in[98] = (SAXISRQTDATA[98] === 1'bz) || SAXISRQTDATA_delay[98]; // rv 1
  assign SAXISRQTDATA_in[99] = (SAXISRQTDATA[99] === 1'bz) || SAXISRQTDATA_delay[99]; // rv 1
  assign SAXISRQTDATA_in[9] = (SAXISRQTDATA[9] === 1'bz) || SAXISRQTDATA_delay[9]; // rv 1
  assign SAXISRQTKEEP_in[0] = (SAXISRQTKEEP[0] !== 1'bz) && SAXISRQTKEEP_delay[0]; // rv 0
  assign SAXISRQTKEEP_in[1] = (SAXISRQTKEEP[1] !== 1'bz) && SAXISRQTKEEP_delay[1]; // rv 0
  assign SAXISRQTKEEP_in[2] = (SAXISRQTKEEP[2] !== 1'bz) && SAXISRQTKEEP_delay[2]; // rv 0
  assign SAXISRQTKEEP_in[3] = (SAXISRQTKEEP[3] !== 1'bz) && SAXISRQTKEEP_delay[3]; // rv 0
  assign SAXISRQTKEEP_in[4] = (SAXISRQTKEEP[4] !== 1'bz) && SAXISRQTKEEP_delay[4]; // rv 0
  assign SAXISRQTKEEP_in[5] = (SAXISRQTKEEP[5] !== 1'bz) && SAXISRQTKEEP_delay[5]; // rv 0
  assign SAXISRQTKEEP_in[6] = (SAXISRQTKEEP[6] !== 1'bz) && SAXISRQTKEEP_delay[6]; // rv 0
  assign SAXISRQTKEEP_in[7] = (SAXISRQTKEEP[7] !== 1'bz) && SAXISRQTKEEP_delay[7]; // rv 0
  assign SAXISRQTLAST_in = (SAXISRQTLAST === 1'bz) || SAXISRQTLAST_delay; // rv 1
  assign SAXISRQTUSER_in[0] = (SAXISRQTUSER[0] === 1'bz) || SAXISRQTUSER_delay[0]; // rv 1
  assign SAXISRQTUSER_in[10] = (SAXISRQTUSER[10] === 1'bz) || SAXISRQTUSER_delay[10]; // rv 1
  assign SAXISRQTUSER_in[11] = (SAXISRQTUSER[11] === 1'bz) || SAXISRQTUSER_delay[11]; // rv 1
  assign SAXISRQTUSER_in[12] = (SAXISRQTUSER[12] === 1'bz) || SAXISRQTUSER_delay[12]; // rv 1
  assign SAXISRQTUSER_in[13] = (SAXISRQTUSER[13] === 1'bz) || SAXISRQTUSER_delay[13]; // rv 1
  assign SAXISRQTUSER_in[14] = (SAXISRQTUSER[14] === 1'bz) || SAXISRQTUSER_delay[14]; // rv 1
  assign SAXISRQTUSER_in[15] = (SAXISRQTUSER[15] === 1'bz) || SAXISRQTUSER_delay[15]; // rv 1
  assign SAXISRQTUSER_in[16] = (SAXISRQTUSER[16] === 1'bz) || SAXISRQTUSER_delay[16]; // rv 1
  assign SAXISRQTUSER_in[17] = (SAXISRQTUSER[17] === 1'bz) || SAXISRQTUSER_delay[17]; // rv 1
  assign SAXISRQTUSER_in[18] = (SAXISRQTUSER[18] === 1'bz) || SAXISRQTUSER_delay[18]; // rv 1
  assign SAXISRQTUSER_in[19] = (SAXISRQTUSER[19] === 1'bz) || SAXISRQTUSER_delay[19]; // rv 1
  assign SAXISRQTUSER_in[1] = (SAXISRQTUSER[1] === 1'bz) || SAXISRQTUSER_delay[1]; // rv 1
  assign SAXISRQTUSER_in[20] = (SAXISRQTUSER[20] === 1'bz) || SAXISRQTUSER_delay[20]; // rv 1
  assign SAXISRQTUSER_in[21] = (SAXISRQTUSER[21] === 1'bz) || SAXISRQTUSER_delay[21]; // rv 1
  assign SAXISRQTUSER_in[22] = (SAXISRQTUSER[22] === 1'bz) || SAXISRQTUSER_delay[22]; // rv 1
  assign SAXISRQTUSER_in[23] = (SAXISRQTUSER[23] === 1'bz) || SAXISRQTUSER_delay[23]; // rv 1
  assign SAXISRQTUSER_in[24] = (SAXISRQTUSER[24] === 1'bz) || SAXISRQTUSER_delay[24]; // rv 1
  assign SAXISRQTUSER_in[25] = (SAXISRQTUSER[25] === 1'bz) || SAXISRQTUSER_delay[25]; // rv 1
  assign SAXISRQTUSER_in[26] = (SAXISRQTUSER[26] === 1'bz) || SAXISRQTUSER_delay[26]; // rv 1
  assign SAXISRQTUSER_in[27] = (SAXISRQTUSER[27] === 1'bz) || SAXISRQTUSER_delay[27]; // rv 1
  assign SAXISRQTUSER_in[28] = (SAXISRQTUSER[28] === 1'bz) || SAXISRQTUSER_delay[28]; // rv 1
  assign SAXISRQTUSER_in[29] = (SAXISRQTUSER[29] === 1'bz) || SAXISRQTUSER_delay[29]; // rv 1
  assign SAXISRQTUSER_in[2] = (SAXISRQTUSER[2] === 1'bz) || SAXISRQTUSER_delay[2]; // rv 1
  assign SAXISRQTUSER_in[30] = (SAXISRQTUSER[30] === 1'bz) || SAXISRQTUSER_delay[30]; // rv 1
  assign SAXISRQTUSER_in[31] = (SAXISRQTUSER[31] === 1'bz) || SAXISRQTUSER_delay[31]; // rv 1
  assign SAXISRQTUSER_in[32] = (SAXISRQTUSER[32] === 1'bz) || SAXISRQTUSER_delay[32]; // rv 1
  assign SAXISRQTUSER_in[33] = (SAXISRQTUSER[33] === 1'bz) || SAXISRQTUSER_delay[33]; // rv 1
  assign SAXISRQTUSER_in[34] = (SAXISRQTUSER[34] === 1'bz) || SAXISRQTUSER_delay[34]; // rv 1
  assign SAXISRQTUSER_in[35] = (SAXISRQTUSER[35] === 1'bz) || SAXISRQTUSER_delay[35]; // rv 1
  assign SAXISRQTUSER_in[36] = (SAXISRQTUSER[36] === 1'bz) || SAXISRQTUSER_delay[36]; // rv 1
  assign SAXISRQTUSER_in[37] = (SAXISRQTUSER[37] === 1'bz) || SAXISRQTUSER_delay[37]; // rv 1
  assign SAXISRQTUSER_in[38] = (SAXISRQTUSER[38] === 1'bz) || SAXISRQTUSER_delay[38]; // rv 1
  assign SAXISRQTUSER_in[39] = (SAXISRQTUSER[39] === 1'bz) || SAXISRQTUSER_delay[39]; // rv 1
  assign SAXISRQTUSER_in[3] = (SAXISRQTUSER[3] === 1'bz) || SAXISRQTUSER_delay[3]; // rv 1
  assign SAXISRQTUSER_in[40] = (SAXISRQTUSER[40] === 1'bz) || SAXISRQTUSER_delay[40]; // rv 1
  assign SAXISRQTUSER_in[41] = (SAXISRQTUSER[41] === 1'bz) || SAXISRQTUSER_delay[41]; // rv 1
  assign SAXISRQTUSER_in[42] = (SAXISRQTUSER[42] === 1'bz) || SAXISRQTUSER_delay[42]; // rv 1
  assign SAXISRQTUSER_in[43] = (SAXISRQTUSER[43] === 1'bz) || SAXISRQTUSER_delay[43]; // rv 1
  assign SAXISRQTUSER_in[44] = (SAXISRQTUSER[44] === 1'bz) || SAXISRQTUSER_delay[44]; // rv 1
  assign SAXISRQTUSER_in[45] = (SAXISRQTUSER[45] === 1'bz) || SAXISRQTUSER_delay[45]; // rv 1
  assign SAXISRQTUSER_in[46] = (SAXISRQTUSER[46] === 1'bz) || SAXISRQTUSER_delay[46]; // rv 1
  assign SAXISRQTUSER_in[47] = (SAXISRQTUSER[47] === 1'bz) || SAXISRQTUSER_delay[47]; // rv 1
  assign SAXISRQTUSER_in[48] = (SAXISRQTUSER[48] === 1'bz) || SAXISRQTUSER_delay[48]; // rv 1
  assign SAXISRQTUSER_in[49] = (SAXISRQTUSER[49] === 1'bz) || SAXISRQTUSER_delay[49]; // rv 1
  assign SAXISRQTUSER_in[4] = (SAXISRQTUSER[4] === 1'bz) || SAXISRQTUSER_delay[4]; // rv 1
  assign SAXISRQTUSER_in[50] = (SAXISRQTUSER[50] === 1'bz) || SAXISRQTUSER_delay[50]; // rv 1
  assign SAXISRQTUSER_in[51] = (SAXISRQTUSER[51] === 1'bz) || SAXISRQTUSER_delay[51]; // rv 1
  assign SAXISRQTUSER_in[52] = (SAXISRQTUSER[52] === 1'bz) || SAXISRQTUSER_delay[52]; // rv 1
  assign SAXISRQTUSER_in[53] = (SAXISRQTUSER[53] === 1'bz) || SAXISRQTUSER_delay[53]; // rv 1
  assign SAXISRQTUSER_in[54] = (SAXISRQTUSER[54] === 1'bz) || SAXISRQTUSER_delay[54]; // rv 1
  assign SAXISRQTUSER_in[55] = (SAXISRQTUSER[55] === 1'bz) || SAXISRQTUSER_delay[55]; // rv 1
  assign SAXISRQTUSER_in[56] = (SAXISRQTUSER[56] === 1'bz) || SAXISRQTUSER_delay[56]; // rv 1
  assign SAXISRQTUSER_in[57] = (SAXISRQTUSER[57] === 1'bz) || SAXISRQTUSER_delay[57]; // rv 1
  assign SAXISRQTUSER_in[58] = (SAXISRQTUSER[58] === 1'bz) || SAXISRQTUSER_delay[58]; // rv 1
  assign SAXISRQTUSER_in[59] = (SAXISRQTUSER[59] === 1'bz) || SAXISRQTUSER_delay[59]; // rv 1
  assign SAXISRQTUSER_in[5] = (SAXISRQTUSER[5] === 1'bz) || SAXISRQTUSER_delay[5]; // rv 1
  assign SAXISRQTUSER_in[6] = (SAXISRQTUSER[6] === 1'bz) || SAXISRQTUSER_delay[6]; // rv 1
  assign SAXISRQTUSER_in[7] = (SAXISRQTUSER[7] === 1'bz) || SAXISRQTUSER_delay[7]; // rv 1
  assign SAXISRQTUSER_in[8] = (SAXISRQTUSER[8] === 1'bz) || SAXISRQTUSER_delay[8]; // rv 1
  assign SAXISRQTUSER_in[9] = (SAXISRQTUSER[9] === 1'bz) || SAXISRQTUSER_delay[9]; // rv 1
  assign SAXISRQTVALID_in = (SAXISRQTVALID !== 1'bz) && SAXISRQTVALID_delay; // rv 0
  assign SPAREIN_in[0] = (SPAREIN[0] === 1'bz) || SPAREIN_delay[0]; // rv 1
  assign SPAREIN_in[10] = (SPAREIN[10] === 1'bz) || SPAREIN_delay[10]; // rv 1
  assign SPAREIN_in[11] = (SPAREIN[11] === 1'bz) || SPAREIN_delay[11]; // rv 1
  assign SPAREIN_in[12] = (SPAREIN[12] === 1'bz) || SPAREIN_delay[12]; // rv 1
  assign SPAREIN_in[13] = (SPAREIN[13] === 1'bz) || SPAREIN_delay[13]; // rv 1
  assign SPAREIN_in[14] = (SPAREIN[14] === 1'bz) || SPAREIN_delay[14]; // rv 1
  assign SPAREIN_in[15] = (SPAREIN[15] === 1'bz) || SPAREIN_delay[15]; // rv 1
  assign SPAREIN_in[16] = (SPAREIN[16] === 1'bz) || SPAREIN_delay[16]; // rv 1
  assign SPAREIN_in[17] = (SPAREIN[17] === 1'bz) || SPAREIN_delay[17]; // rv 1
  assign SPAREIN_in[18] = (SPAREIN[18] === 1'bz) || SPAREIN_delay[18]; // rv 1
  assign SPAREIN_in[19] = (SPAREIN[19] === 1'bz) || SPAREIN_delay[19]; // rv 1
  assign SPAREIN_in[1] = (SPAREIN[1] === 1'bz) || SPAREIN_delay[1]; // rv 1
  assign SPAREIN_in[20] = (SPAREIN[20] === 1'bz) || SPAREIN_delay[20]; // rv 1
  assign SPAREIN_in[21] = (SPAREIN[21] === 1'bz) || SPAREIN_delay[21]; // rv 1
  assign SPAREIN_in[22] = (SPAREIN[22] === 1'bz) || SPAREIN_delay[22]; // rv 1
  assign SPAREIN_in[23] = (SPAREIN[23] === 1'bz) || SPAREIN_delay[23]; // rv 1
  assign SPAREIN_in[24] = (SPAREIN[24] === 1'bz) || SPAREIN_delay[24]; // rv 1
  assign SPAREIN_in[25] = (SPAREIN[25] === 1'bz) || SPAREIN_delay[25]; // rv 1
  assign SPAREIN_in[26] = (SPAREIN[26] === 1'bz) || SPAREIN_delay[26]; // rv 1
  assign SPAREIN_in[27] = (SPAREIN[27] === 1'bz) || SPAREIN_delay[27]; // rv 1
  assign SPAREIN_in[28] = (SPAREIN[28] === 1'bz) || SPAREIN_delay[28]; // rv 1
  assign SPAREIN_in[29] = (SPAREIN[29] === 1'bz) || SPAREIN_delay[29]; // rv 1
  assign SPAREIN_in[2] = (SPAREIN[2] === 1'bz) || SPAREIN_delay[2]; // rv 1
  assign SPAREIN_in[30] = (SPAREIN[30] === 1'bz) || SPAREIN_delay[30]; // rv 1
  assign SPAREIN_in[31] = (SPAREIN[31] === 1'bz) || SPAREIN_delay[31]; // rv 1
  assign SPAREIN_in[3] = (SPAREIN[3] === 1'bz) || SPAREIN_delay[3]; // rv 1
  assign SPAREIN_in[4] = (SPAREIN[4] === 1'bz) || SPAREIN_delay[4]; // rv 1
  assign SPAREIN_in[5] = (SPAREIN[5] === 1'bz) || SPAREIN_delay[5]; // rv 1
  assign SPAREIN_in[6] = (SPAREIN[6] === 1'bz) || SPAREIN_delay[6]; // rv 1
  assign SPAREIN_in[7] = (SPAREIN[7] === 1'bz) || SPAREIN_delay[7]; // rv 1
  assign SPAREIN_in[8] = (SPAREIN[8] === 1'bz) || SPAREIN_delay[8]; // rv 1
  assign SPAREIN_in[9] = (SPAREIN[9] === 1'bz) || SPAREIN_delay[9]; // rv 1
  assign USERCLK_in = (USERCLK !== 1'bz) && USERCLK_delay; // rv 0


  initial begin
  #1;
  trig_attr = ~trig_attr;
  end

  always @ (trig_attr) begin
    #1;
    if ((ARI_CAP_ENABLE_REG != "FALSE") &&
        (ARI_CAP_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute ARI_CAP_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, ARI_CAP_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((AXISTEN_IF_CC_ALIGNMENT_MODE_REG != "FALSE") &&
        (AXISTEN_IF_CC_ALIGNMENT_MODE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute AXISTEN_IF_CC_ALIGNMENT_MODE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, AXISTEN_IF_CC_ALIGNMENT_MODE_REG);
      attr_err = 1'b1;
    end

    if ((AXISTEN_IF_CC_PARITY_CHK_REG != "TRUE") &&
        (AXISTEN_IF_CC_PARITY_CHK_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute AXISTEN_IF_CC_PARITY_CHK on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, AXISTEN_IF_CC_PARITY_CHK_REG);
      attr_err = 1'b1;
    end

    if ((AXISTEN_IF_CQ_ALIGNMENT_MODE_REG != "FALSE") &&
        (AXISTEN_IF_CQ_ALIGNMENT_MODE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute AXISTEN_IF_CQ_ALIGNMENT_MODE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, AXISTEN_IF_CQ_ALIGNMENT_MODE_REG);
      attr_err = 1'b1;
    end

    if ((AXISTEN_IF_ENABLE_CLIENT_TAG_REG != "FALSE") &&
        (AXISTEN_IF_ENABLE_CLIENT_TAG_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute AXISTEN_IF_ENABLE_CLIENT_TAG on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, AXISTEN_IF_ENABLE_CLIENT_TAG_REG);
      attr_err = 1'b1;
    end

    if ((AXISTEN_IF_ENABLE_RX_MSG_INTFC_REG != "FALSE") &&
        (AXISTEN_IF_ENABLE_RX_MSG_INTFC_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute AXISTEN_IF_ENABLE_RX_MSG_INTFC on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, AXISTEN_IF_ENABLE_RX_MSG_INTFC_REG);
      attr_err = 1'b1;
    end

    if ((AXISTEN_IF_RC_ALIGNMENT_MODE_REG != "FALSE") &&
        (AXISTEN_IF_RC_ALIGNMENT_MODE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute AXISTEN_IF_RC_ALIGNMENT_MODE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, AXISTEN_IF_RC_ALIGNMENT_MODE_REG);
      attr_err = 1'b1;
    end

    if ((AXISTEN_IF_RC_STRADDLE_REG != "FALSE") &&
        (AXISTEN_IF_RC_STRADDLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute AXISTEN_IF_RC_STRADDLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, AXISTEN_IF_RC_STRADDLE_REG);
      attr_err = 1'b1;
    end

    if ((AXISTEN_IF_RQ_ALIGNMENT_MODE_REG != "FALSE") &&
        (AXISTEN_IF_RQ_ALIGNMENT_MODE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute AXISTEN_IF_RQ_ALIGNMENT_MODE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, AXISTEN_IF_RQ_ALIGNMENT_MODE_REG);
      attr_err = 1'b1;
    end

    if ((AXISTEN_IF_RQ_PARITY_CHK_REG != "TRUE") &&
        (AXISTEN_IF_RQ_PARITY_CHK_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute AXISTEN_IF_RQ_PARITY_CHK on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, AXISTEN_IF_RQ_PARITY_CHK_REG);
      attr_err = 1'b1;
    end

    if ((CRM_CORE_CLK_FREQ_500_REG != "TRUE") &&
        (CRM_CORE_CLK_FREQ_500_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute CRM_CORE_CLK_FREQ_500 on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, CRM_CORE_CLK_FREQ_500_REG);
      attr_err = 1'b1;
    end

    if ((DEBUG_CFG_LOCAL_MGMT_REG_ACCESS_OVERRIDE_REG != "FALSE") &&
        (DEBUG_CFG_LOCAL_MGMT_REG_ACCESS_OVERRIDE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute DEBUG_CFG_LOCAL_MGMT_REG_ACCESS_OVERRIDE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, DEBUG_CFG_LOCAL_MGMT_REG_ACCESS_OVERRIDE_REG);
      attr_err = 1'b1;
    end

    if ((DEBUG_PL_DISABLE_EI_INFER_IN_L0_REG != "FALSE") &&
        (DEBUG_PL_DISABLE_EI_INFER_IN_L0_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute DEBUG_PL_DISABLE_EI_INFER_IN_L0 on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, DEBUG_PL_DISABLE_EI_INFER_IN_L0_REG);
      attr_err = 1'b1;
    end

    if ((DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS_REG != "FALSE") &&
        (DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS_REG);
      attr_err = 1'b1;
    end

    if ((LL_ACK_TIMEOUT_EN_REG != "FALSE") &&
        (LL_ACK_TIMEOUT_EN_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute LL_ACK_TIMEOUT_EN on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, LL_ACK_TIMEOUT_EN_REG);
      attr_err = 1'b1;
    end

    if ((LL_ACK_TIMEOUT_FUNC_REG != 0) &&
        (LL_ACK_TIMEOUT_FUNC_REG != 1) &&
        (LL_ACK_TIMEOUT_FUNC_REG != 2) &&
        (LL_ACK_TIMEOUT_FUNC_REG != 3)) begin
      $display("Attribute Syntax Error : The attribute LL_ACK_TIMEOUT_FUNC on %s instance %m is set to %d.  Legal values for this attribute are 0 to 3.", MODULE_NAME, LL_ACK_TIMEOUT_FUNC_REG);
      attr_err = 1'b1;
    end

    if ((LL_CPL_FC_UPDATE_TIMER_OVERRIDE_REG != "FALSE") &&
        (LL_CPL_FC_UPDATE_TIMER_OVERRIDE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute LL_CPL_FC_UPDATE_TIMER_OVERRIDE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, LL_CPL_FC_UPDATE_TIMER_OVERRIDE_REG);
      attr_err = 1'b1;
    end

    if ((LL_FC_UPDATE_TIMER_OVERRIDE_REG != "FALSE") &&
        (LL_FC_UPDATE_TIMER_OVERRIDE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute LL_FC_UPDATE_TIMER_OVERRIDE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, LL_FC_UPDATE_TIMER_OVERRIDE_REG);
      attr_err = 1'b1;
    end

    if ((LL_NP_FC_UPDATE_TIMER_OVERRIDE_REG != "FALSE") &&
        (LL_NP_FC_UPDATE_TIMER_OVERRIDE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute LL_NP_FC_UPDATE_TIMER_OVERRIDE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, LL_NP_FC_UPDATE_TIMER_OVERRIDE_REG);
      attr_err = 1'b1;
    end

    if ((LL_P_FC_UPDATE_TIMER_OVERRIDE_REG != "FALSE") &&
        (LL_P_FC_UPDATE_TIMER_OVERRIDE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute LL_P_FC_UPDATE_TIMER_OVERRIDE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, LL_P_FC_UPDATE_TIMER_OVERRIDE_REG);
      attr_err = 1'b1;
    end

    if ((LL_REPLAY_TIMEOUT_EN_REG != "FALSE") &&
        (LL_REPLAY_TIMEOUT_EN_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute LL_REPLAY_TIMEOUT_EN on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, LL_REPLAY_TIMEOUT_EN_REG);
      attr_err = 1'b1;
    end

    if ((LL_REPLAY_TIMEOUT_FUNC_REG != 0) &&
        (LL_REPLAY_TIMEOUT_FUNC_REG != 1) &&
        (LL_REPLAY_TIMEOUT_FUNC_REG != 2) &&
        (LL_REPLAY_TIMEOUT_FUNC_REG != 3)) begin
      $display("Attribute Syntax Error : The attribute LL_REPLAY_TIMEOUT_FUNC on %s instance %m is set to %d.  Legal values for this attribute are 0 to 3.", MODULE_NAME, LL_REPLAY_TIMEOUT_FUNC_REG);
      attr_err = 1'b1;
    end

    if ((LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE_REG != "FALSE") &&
        (LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE_REG);
      attr_err = 1'b1;
    end

    if ((LTR_TX_MESSAGE_ON_LTR_ENABLE_REG != "FALSE") &&
        (LTR_TX_MESSAGE_ON_LTR_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute LTR_TX_MESSAGE_ON_LTR_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, LTR_TX_MESSAGE_ON_LTR_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((MCAP_CONFIGURE_OVERRIDE_REG != "FALSE") &&
        (MCAP_CONFIGURE_OVERRIDE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute MCAP_CONFIGURE_OVERRIDE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, MCAP_CONFIGURE_OVERRIDE_REG);
      attr_err = 1'b1;
    end

    if ((MCAP_ENABLE_REG != "FALSE") &&
        (MCAP_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute MCAP_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, MCAP_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((MCAP_EOS_DESIGN_SWITCH_REG != "FALSE") &&
        (MCAP_EOS_DESIGN_SWITCH_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute MCAP_EOS_DESIGN_SWITCH on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, MCAP_EOS_DESIGN_SWITCH_REG);
      attr_err = 1'b1;
    end

    if ((MCAP_GATE_IO_ENABLE_DESIGN_SWITCH_REG != "FALSE") &&
        (MCAP_GATE_IO_ENABLE_DESIGN_SWITCH_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute MCAP_GATE_IO_ENABLE_DESIGN_SWITCH on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, MCAP_GATE_IO_ENABLE_DESIGN_SWITCH_REG);
      attr_err = 1'b1;
    end

    if ((MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH_REG != "FALSE") &&
        (MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH_REG);
      attr_err = 1'b1;
    end

    if ((MCAP_INPUT_GATE_DESIGN_SWITCH_REG != "FALSE") &&
        (MCAP_INPUT_GATE_DESIGN_SWITCH_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute MCAP_INPUT_GATE_DESIGN_SWITCH on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, MCAP_INPUT_GATE_DESIGN_SWITCH_REG);
      attr_err = 1'b1;
    end

    if ((MCAP_INTERRUPT_ON_MCAP_EOS_REG != "FALSE") &&
        (MCAP_INTERRUPT_ON_MCAP_EOS_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute MCAP_INTERRUPT_ON_MCAP_EOS on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, MCAP_INTERRUPT_ON_MCAP_EOS_REG);
      attr_err = 1'b1;
    end

    if ((MCAP_INTERRUPT_ON_MCAP_ERROR_REG != "FALSE") &&
        (MCAP_INTERRUPT_ON_MCAP_ERROR_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute MCAP_INTERRUPT_ON_MCAP_ERROR on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, MCAP_INTERRUPT_ON_MCAP_ERROR_REG);
      attr_err = 1'b1;
    end

    if ((PF0_AER_CAP_ECRC_CHECK_CAPABLE_REG != "FALSE") &&
        (PF0_AER_CAP_ECRC_CHECK_CAPABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF0_AER_CAP_ECRC_CHECK_CAPABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF0_AER_CAP_ECRC_CHECK_CAPABLE_REG);
      attr_err = 1'b1;
    end

    if ((PF0_AER_CAP_ECRC_GEN_CAPABLE_REG != "FALSE") &&
        (PF0_AER_CAP_ECRC_GEN_CAPABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF0_AER_CAP_ECRC_GEN_CAPABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF0_AER_CAP_ECRC_GEN_CAPABLE_REG);
      attr_err = 1'b1;
    end

    if ((PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT_REG != "TRUE") &&
        (PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT_REG);
      attr_err = 1'b1;
    end

    if ((PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT_REG != "TRUE") &&
        (PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT_REG);
      attr_err = 1'b1;
    end

    if ((PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT_REG != "TRUE") &&
        (PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT_REG);
      attr_err = 1'b1;
    end

    if ((PF0_DEV_CAP2_ARI_FORWARD_ENABLE_REG != "FALSE") &&
        (PF0_DEV_CAP2_ARI_FORWARD_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF0_DEV_CAP2_ARI_FORWARD_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF0_DEV_CAP2_ARI_FORWARD_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE_REG != "TRUE") &&
        (PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE_REG);
      attr_err = 1'b1;
    end

    if ((PF0_DEV_CAP2_LTR_SUPPORT_REG != "TRUE") &&
        (PF0_DEV_CAP2_LTR_SUPPORT_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PF0_DEV_CAP2_LTR_SUPPORT on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PF0_DEV_CAP2_LTR_SUPPORT_REG);
      attr_err = 1'b1;
    end

    if ((PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT_REG != "FALSE") &&
        (PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT_REG);
      attr_err = 1'b1;
    end

    if ((PF0_DEV_CAP_ENDPOINT_L0S_LATENCY_REG != 0) &&
        (PF0_DEV_CAP_ENDPOINT_L0S_LATENCY_REG != 1) &&
        (PF0_DEV_CAP_ENDPOINT_L0S_LATENCY_REG != 2) &&
        (PF0_DEV_CAP_ENDPOINT_L0S_LATENCY_REG != 3) &&
        (PF0_DEV_CAP_ENDPOINT_L0S_LATENCY_REG != 4) &&
        (PF0_DEV_CAP_ENDPOINT_L0S_LATENCY_REG != 5) &&
        (PF0_DEV_CAP_ENDPOINT_L0S_LATENCY_REG != 6) &&
        (PF0_DEV_CAP_ENDPOINT_L0S_LATENCY_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute PF0_DEV_CAP_ENDPOINT_L0S_LATENCY on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, PF0_DEV_CAP_ENDPOINT_L0S_LATENCY_REG);
      attr_err = 1'b1;
    end

    if ((PF0_DEV_CAP_ENDPOINT_L1_LATENCY_REG != 0) &&
        (PF0_DEV_CAP_ENDPOINT_L1_LATENCY_REG != 1) &&
        (PF0_DEV_CAP_ENDPOINT_L1_LATENCY_REG != 2) &&
        (PF0_DEV_CAP_ENDPOINT_L1_LATENCY_REG != 3) &&
        (PF0_DEV_CAP_ENDPOINT_L1_LATENCY_REG != 4) &&
        (PF0_DEV_CAP_ENDPOINT_L1_LATENCY_REG != 5) &&
        (PF0_DEV_CAP_ENDPOINT_L1_LATENCY_REG != 6) &&
        (PF0_DEV_CAP_ENDPOINT_L1_LATENCY_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute PF0_DEV_CAP_ENDPOINT_L1_LATENCY on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, PF0_DEV_CAP_ENDPOINT_L1_LATENCY_REG);
      attr_err = 1'b1;
    end

    if ((PF0_DEV_CAP_EXT_TAG_SUPPORTED_REG != "TRUE") &&
        (PF0_DEV_CAP_EXT_TAG_SUPPORTED_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PF0_DEV_CAP_EXT_TAG_SUPPORTED on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PF0_DEV_CAP_EXT_TAG_SUPPORTED_REG);
      attr_err = 1'b1;
    end

    if ((PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE_REG != "TRUE") &&
        (PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE_REG);
      attr_err = 1'b1;
    end

    if ((PF0_DPA_CAP_SUB_STATE_CONTROL_EN_REG != "TRUE") &&
        (PF0_DPA_CAP_SUB_STATE_CONTROL_EN_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PF0_DPA_CAP_SUB_STATE_CONTROL_EN on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PF0_DPA_CAP_SUB_STATE_CONTROL_EN_REG);
      attr_err = 1'b1;
    end

    if ((PF0_EXPANSION_ROM_ENABLE_REG != "FALSE") &&
        (PF0_EXPANSION_ROM_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF0_EXPANSION_ROM_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF0_EXPANSION_ROM_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((PF0_LINK_CAP_ASPM_SUPPORT_REG != 0) &&
        (PF0_LINK_CAP_ASPM_SUPPORT_REG != 1) &&
        (PF0_LINK_CAP_ASPM_SUPPORT_REG != 2) &&
        (PF0_LINK_CAP_ASPM_SUPPORT_REG != 3)) begin
      $display("Attribute Syntax Error : The attribute PF0_LINK_CAP_ASPM_SUPPORT on %s instance %m is set to %d.  Legal values for this attribute are 0 to 3.", MODULE_NAME, PF0_LINK_CAP_ASPM_SUPPORT_REG);
      attr_err = 1'b1;
    end

    if ((PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1_REG != 7) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1_REG != 0) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1_REG != 1) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1_REG != 2) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1_REG != 3) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1_REG != 4) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1_REG != 5) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1_REG != 6)) begin
      $display("Attribute Syntax Error : The attribute PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1_REG);
      attr_err = 1'b1;
    end

    if ((PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2_REG != 7) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2_REG != 0) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2_REG != 1) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2_REG != 2) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2_REG != 3) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2_REG != 4) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2_REG != 5) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2_REG != 6)) begin
      $display("Attribute Syntax Error : The attribute PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2_REG);
      attr_err = 1'b1;
    end

    if ((PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3_REG != 7) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3_REG != 0) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3_REG != 1) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3_REG != 2) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3_REG != 3) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3_REG != 4) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3_REG != 5) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3_REG != 6)) begin
      $display("Attribute Syntax Error : The attribute PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3 on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3_REG);
      attr_err = 1'b1;
    end

    if ((PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1_REG != 7) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1_REG != 0) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1_REG != 1) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1_REG != 2) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1_REG != 3) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1_REG != 4) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1_REG != 5) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1_REG != 6)) begin
      $display("Attribute Syntax Error : The attribute PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1 on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1_REG);
      attr_err = 1'b1;
    end

    if ((PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2_REG != 7) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2_REG != 0) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2_REG != 1) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2_REG != 2) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2_REG != 3) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2_REG != 4) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2_REG != 5) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2_REG != 6)) begin
      $display("Attribute Syntax Error : The attribute PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2 on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2_REG);
      attr_err = 1'b1;
    end

    if ((PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3_REG != 7) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3_REG != 0) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3_REG != 1) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3_REG != 2) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3_REG != 3) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3_REG != 4) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3_REG != 5) &&
        (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3_REG != 6)) begin
      $display("Attribute Syntax Error : The attribute PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3 on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3_REG);
      attr_err = 1'b1;
    end

    if ((PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1_REG != 7) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1_REG != 0) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1_REG != 1) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1_REG != 2) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1_REG != 3) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1_REG != 4) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1_REG != 5) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1_REG != 6)) begin
      $display("Attribute Syntax Error : The attribute PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1_REG);
      attr_err = 1'b1;
    end

    if ((PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2_REG != 7) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2_REG != 0) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2_REG != 1) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2_REG != 2) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2_REG != 3) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2_REG != 4) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2_REG != 5) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2_REG != 6)) begin
      $display("Attribute Syntax Error : The attribute PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2_REG);
      attr_err = 1'b1;
    end

    if ((PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3_REG != 7) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3_REG != 0) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3_REG != 1) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3_REG != 2) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3_REG != 3) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3_REG != 4) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3_REG != 5) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3_REG != 6)) begin
      $display("Attribute Syntax Error : The attribute PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3 on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3_REG);
      attr_err = 1'b1;
    end

    if ((PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1_REG != 7) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1_REG != 0) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1_REG != 1) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1_REG != 2) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1_REG != 3) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1_REG != 4) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1_REG != 5) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1_REG != 6)) begin
      $display("Attribute Syntax Error : The attribute PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1 on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1_REG);
      attr_err = 1'b1;
    end

    if ((PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2_REG != 7) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2_REG != 0) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2_REG != 1) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2_REG != 2) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2_REG != 3) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2_REG != 4) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2_REG != 5) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2_REG != 6)) begin
      $display("Attribute Syntax Error : The attribute PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2 on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2_REG);
      attr_err = 1'b1;
    end

    if ((PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3_REG != 7) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3_REG != 0) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3_REG != 1) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3_REG != 2) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3_REG != 3) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3_REG != 4) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3_REG != 5) &&
        (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3_REG != 6)) begin
      $display("Attribute Syntax Error : The attribute PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3 on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3_REG);
      attr_err = 1'b1;
    end

    if ((PF0_LINK_STATUS_SLOT_CLOCK_CONFIG_REG != "TRUE") &&
        (PF0_LINK_STATUS_SLOT_CLOCK_CONFIG_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PF0_LINK_STATUS_SLOT_CLOCK_CONFIG on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PF0_LINK_STATUS_SLOT_CLOCK_CONFIG_REG);
      attr_err = 1'b1;
    end

    if ((PF0_MSIX_CAP_PBA_BIR_REG != 0) &&
        (PF0_MSIX_CAP_PBA_BIR_REG != 1) &&
        (PF0_MSIX_CAP_PBA_BIR_REG != 2) &&
        (PF0_MSIX_CAP_PBA_BIR_REG != 3) &&
        (PF0_MSIX_CAP_PBA_BIR_REG != 4) &&
        (PF0_MSIX_CAP_PBA_BIR_REG != 5) &&
        (PF0_MSIX_CAP_PBA_BIR_REG != 6) &&
        (PF0_MSIX_CAP_PBA_BIR_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute PF0_MSIX_CAP_PBA_BIR on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, PF0_MSIX_CAP_PBA_BIR_REG);
      attr_err = 1'b1;
    end

    if ((PF0_MSIX_CAP_TABLE_BIR_REG != 0) &&
        (PF0_MSIX_CAP_TABLE_BIR_REG != 1) &&
        (PF0_MSIX_CAP_TABLE_BIR_REG != 2) &&
        (PF0_MSIX_CAP_TABLE_BIR_REG != 3) &&
        (PF0_MSIX_CAP_TABLE_BIR_REG != 4) &&
        (PF0_MSIX_CAP_TABLE_BIR_REG != 5) &&
        (PF0_MSIX_CAP_TABLE_BIR_REG != 6) &&
        (PF0_MSIX_CAP_TABLE_BIR_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute PF0_MSIX_CAP_TABLE_BIR on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, PF0_MSIX_CAP_TABLE_BIR_REG);
      attr_err = 1'b1;
    end

    if ((PF0_MSI_CAP_MULTIMSGCAP_REG != 0) &&
        (PF0_MSI_CAP_MULTIMSGCAP_REG != 1) &&
        (PF0_MSI_CAP_MULTIMSGCAP_REG != 2) &&
        (PF0_MSI_CAP_MULTIMSGCAP_REG != 3) &&
        (PF0_MSI_CAP_MULTIMSGCAP_REG != 4) &&
        (PF0_MSI_CAP_MULTIMSGCAP_REG != 5) &&
        (PF0_MSI_CAP_MULTIMSGCAP_REG != 6) &&
        (PF0_MSI_CAP_MULTIMSGCAP_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute PF0_MSI_CAP_MULTIMSGCAP on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, PF0_MSI_CAP_MULTIMSGCAP_REG);
      attr_err = 1'b1;
    end

    if ((PF0_MSI_CAP_PERVECMASKCAP_REG != "FALSE") &&
        (PF0_MSI_CAP_PERVECMASKCAP_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF0_MSI_CAP_PERVECMASKCAP on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF0_MSI_CAP_PERVECMASKCAP_REG);
      attr_err = 1'b1;
    end

    if ((PF0_PB_CAP_SYSTEM_ALLOCATED_REG != "FALSE") &&
        (PF0_PB_CAP_SYSTEM_ALLOCATED_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF0_PB_CAP_SYSTEM_ALLOCATED on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF0_PB_CAP_SYSTEM_ALLOCATED_REG);
      attr_err = 1'b1;
    end

    if ((PF0_PM_CAP_PMESUPPORT_D0_REG != "TRUE") &&
        (PF0_PM_CAP_PMESUPPORT_D0_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PF0_PM_CAP_PMESUPPORT_D0 on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PF0_PM_CAP_PMESUPPORT_D0_REG);
      attr_err = 1'b1;
    end

    if ((PF0_PM_CAP_PMESUPPORT_D1_REG != "TRUE") &&
        (PF0_PM_CAP_PMESUPPORT_D1_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PF0_PM_CAP_PMESUPPORT_D1 on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PF0_PM_CAP_PMESUPPORT_D1_REG);
      attr_err = 1'b1;
    end

    if ((PF0_PM_CAP_PMESUPPORT_D3HOT_REG != "TRUE") &&
        (PF0_PM_CAP_PMESUPPORT_D3HOT_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PF0_PM_CAP_PMESUPPORT_D3HOT on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PF0_PM_CAP_PMESUPPORT_D3HOT_REG);
      attr_err = 1'b1;
    end

    if ((PF0_PM_CAP_SUPP_D1_STATE_REG != "TRUE") &&
        (PF0_PM_CAP_SUPP_D1_STATE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PF0_PM_CAP_SUPP_D1_STATE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PF0_PM_CAP_SUPP_D1_STATE_REG);
      attr_err = 1'b1;
    end

    if ((PF0_PM_CSR_NOSOFTRESET_REG != "TRUE") &&
        (PF0_PM_CSR_NOSOFTRESET_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PF0_PM_CSR_NOSOFTRESET on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PF0_PM_CSR_NOSOFTRESET_REG);
      attr_err = 1'b1;
    end

    if ((PF0_RBAR_CAP_ENABLE_REG != "FALSE") &&
        (PF0_RBAR_CAP_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF0_RBAR_CAP_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF0_RBAR_CAP_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((PF0_TPHR_CAP_DEV_SPECIFIC_MODE_REG != "TRUE") &&
        (PF0_TPHR_CAP_DEV_SPECIFIC_MODE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PF0_TPHR_CAP_DEV_SPECIFIC_MODE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PF0_TPHR_CAP_DEV_SPECIFIC_MODE_REG);
      attr_err = 1'b1;
    end

    if ((PF0_TPHR_CAP_ENABLE_REG != "FALSE") &&
        (PF0_TPHR_CAP_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF0_TPHR_CAP_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF0_TPHR_CAP_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((PF0_TPHR_CAP_INT_VEC_MODE_REG != "TRUE") &&
        (PF0_TPHR_CAP_INT_VEC_MODE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PF0_TPHR_CAP_INT_VEC_MODE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PF0_TPHR_CAP_INT_VEC_MODE_REG);
      attr_err = 1'b1;
    end

    if ((PF0_VC_CAP_ENABLE_REG != "FALSE") &&
        (PF0_VC_CAP_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF0_VC_CAP_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF0_VC_CAP_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((PF1_AER_CAP_ECRC_CHECK_CAPABLE_REG != "FALSE") &&
        (PF1_AER_CAP_ECRC_CHECK_CAPABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF1_AER_CAP_ECRC_CHECK_CAPABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF1_AER_CAP_ECRC_CHECK_CAPABLE_REG);
      attr_err = 1'b1;
    end

    if ((PF1_AER_CAP_ECRC_GEN_CAPABLE_REG != "FALSE") &&
        (PF1_AER_CAP_ECRC_GEN_CAPABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF1_AER_CAP_ECRC_GEN_CAPABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF1_AER_CAP_ECRC_GEN_CAPABLE_REG);
      attr_err = 1'b1;
    end

    if ((PF1_DPA_CAP_SUB_STATE_CONTROL_EN_REG != "TRUE") &&
        (PF1_DPA_CAP_SUB_STATE_CONTROL_EN_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PF1_DPA_CAP_SUB_STATE_CONTROL_EN on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PF1_DPA_CAP_SUB_STATE_CONTROL_EN_REG);
      attr_err = 1'b1;
    end

    if ((PF1_EXPANSION_ROM_ENABLE_REG != "FALSE") &&
        (PF1_EXPANSION_ROM_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF1_EXPANSION_ROM_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF1_EXPANSION_ROM_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((PF1_MSIX_CAP_PBA_BIR_REG != 0) &&
        (PF1_MSIX_CAP_PBA_BIR_REG != 1) &&
        (PF1_MSIX_CAP_PBA_BIR_REG != 2) &&
        (PF1_MSIX_CAP_PBA_BIR_REG != 3) &&
        (PF1_MSIX_CAP_PBA_BIR_REG != 4) &&
        (PF1_MSIX_CAP_PBA_BIR_REG != 5) &&
        (PF1_MSIX_CAP_PBA_BIR_REG != 6) &&
        (PF1_MSIX_CAP_PBA_BIR_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute PF1_MSIX_CAP_PBA_BIR on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, PF1_MSIX_CAP_PBA_BIR_REG);
      attr_err = 1'b1;
    end

    if ((PF1_MSIX_CAP_TABLE_BIR_REG != 0) &&
        (PF1_MSIX_CAP_TABLE_BIR_REG != 1) &&
        (PF1_MSIX_CAP_TABLE_BIR_REG != 2) &&
        (PF1_MSIX_CAP_TABLE_BIR_REG != 3) &&
        (PF1_MSIX_CAP_TABLE_BIR_REG != 4) &&
        (PF1_MSIX_CAP_TABLE_BIR_REG != 5) &&
        (PF1_MSIX_CAP_TABLE_BIR_REG != 6) &&
        (PF1_MSIX_CAP_TABLE_BIR_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute PF1_MSIX_CAP_TABLE_BIR on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, PF1_MSIX_CAP_TABLE_BIR_REG);
      attr_err = 1'b1;
    end

    if ((PF1_MSI_CAP_MULTIMSGCAP_REG != 0) &&
        (PF1_MSI_CAP_MULTIMSGCAP_REG != 1) &&
        (PF1_MSI_CAP_MULTIMSGCAP_REG != 2) &&
        (PF1_MSI_CAP_MULTIMSGCAP_REG != 3) &&
        (PF1_MSI_CAP_MULTIMSGCAP_REG != 4) &&
        (PF1_MSI_CAP_MULTIMSGCAP_REG != 5) &&
        (PF1_MSI_CAP_MULTIMSGCAP_REG != 6) &&
        (PF1_MSI_CAP_MULTIMSGCAP_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute PF1_MSI_CAP_MULTIMSGCAP on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, PF1_MSI_CAP_MULTIMSGCAP_REG);
      attr_err = 1'b1;
    end

    if ((PF1_MSI_CAP_PERVECMASKCAP_REG != "FALSE") &&
        (PF1_MSI_CAP_PERVECMASKCAP_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF1_MSI_CAP_PERVECMASKCAP on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF1_MSI_CAP_PERVECMASKCAP_REG);
      attr_err = 1'b1;
    end

    if ((PF1_PB_CAP_SYSTEM_ALLOCATED_REG != "FALSE") &&
        (PF1_PB_CAP_SYSTEM_ALLOCATED_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF1_PB_CAP_SYSTEM_ALLOCATED on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF1_PB_CAP_SYSTEM_ALLOCATED_REG);
      attr_err = 1'b1;
    end

    if ((PF1_RBAR_CAP_ENABLE_REG != "FALSE") &&
        (PF1_RBAR_CAP_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF1_RBAR_CAP_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF1_RBAR_CAP_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((PF1_TPHR_CAP_DEV_SPECIFIC_MODE_REG != "TRUE") &&
        (PF1_TPHR_CAP_DEV_SPECIFIC_MODE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PF1_TPHR_CAP_DEV_SPECIFIC_MODE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PF1_TPHR_CAP_DEV_SPECIFIC_MODE_REG);
      attr_err = 1'b1;
    end

    if ((PF1_TPHR_CAP_ENABLE_REG != "FALSE") &&
        (PF1_TPHR_CAP_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF1_TPHR_CAP_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF1_TPHR_CAP_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((PF1_TPHR_CAP_INT_VEC_MODE_REG != "TRUE") &&
        (PF1_TPHR_CAP_INT_VEC_MODE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PF1_TPHR_CAP_INT_VEC_MODE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PF1_TPHR_CAP_INT_VEC_MODE_REG);
      attr_err = 1'b1;
    end

    if ((PF2_AER_CAP_ECRC_CHECK_CAPABLE_REG != "FALSE") &&
        (PF2_AER_CAP_ECRC_CHECK_CAPABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF2_AER_CAP_ECRC_CHECK_CAPABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF2_AER_CAP_ECRC_CHECK_CAPABLE_REG);
      attr_err = 1'b1;
    end

    if ((PF2_AER_CAP_ECRC_GEN_CAPABLE_REG != "FALSE") &&
        (PF2_AER_CAP_ECRC_GEN_CAPABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF2_AER_CAP_ECRC_GEN_CAPABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF2_AER_CAP_ECRC_GEN_CAPABLE_REG);
      attr_err = 1'b1;
    end

    if ((PF2_DPA_CAP_SUB_STATE_CONTROL_EN_REG != "TRUE") &&
        (PF2_DPA_CAP_SUB_STATE_CONTROL_EN_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PF2_DPA_CAP_SUB_STATE_CONTROL_EN on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PF2_DPA_CAP_SUB_STATE_CONTROL_EN_REG);
      attr_err = 1'b1;
    end

    if ((PF2_EXPANSION_ROM_ENABLE_REG != "FALSE") &&
        (PF2_EXPANSION_ROM_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF2_EXPANSION_ROM_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF2_EXPANSION_ROM_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((PF2_MSIX_CAP_PBA_BIR_REG != 0) &&
        (PF2_MSIX_CAP_PBA_BIR_REG != 1) &&
        (PF2_MSIX_CAP_PBA_BIR_REG != 2) &&
        (PF2_MSIX_CAP_PBA_BIR_REG != 3) &&
        (PF2_MSIX_CAP_PBA_BIR_REG != 4) &&
        (PF2_MSIX_CAP_PBA_BIR_REG != 5) &&
        (PF2_MSIX_CAP_PBA_BIR_REG != 6) &&
        (PF2_MSIX_CAP_PBA_BIR_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute PF2_MSIX_CAP_PBA_BIR on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, PF2_MSIX_CAP_PBA_BIR_REG);
      attr_err = 1'b1;
    end

    if ((PF2_MSIX_CAP_TABLE_BIR_REG != 0) &&
        (PF2_MSIX_CAP_TABLE_BIR_REG != 1) &&
        (PF2_MSIX_CAP_TABLE_BIR_REG != 2) &&
        (PF2_MSIX_CAP_TABLE_BIR_REG != 3) &&
        (PF2_MSIX_CAP_TABLE_BIR_REG != 4) &&
        (PF2_MSIX_CAP_TABLE_BIR_REG != 5) &&
        (PF2_MSIX_CAP_TABLE_BIR_REG != 6) &&
        (PF2_MSIX_CAP_TABLE_BIR_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute PF2_MSIX_CAP_TABLE_BIR on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, PF2_MSIX_CAP_TABLE_BIR_REG);
      attr_err = 1'b1;
    end

    if ((PF2_MSI_CAP_MULTIMSGCAP_REG != 0) &&
        (PF2_MSI_CAP_MULTIMSGCAP_REG != 1) &&
        (PF2_MSI_CAP_MULTIMSGCAP_REG != 2) &&
        (PF2_MSI_CAP_MULTIMSGCAP_REG != 3) &&
        (PF2_MSI_CAP_MULTIMSGCAP_REG != 4) &&
        (PF2_MSI_CAP_MULTIMSGCAP_REG != 5) &&
        (PF2_MSI_CAP_MULTIMSGCAP_REG != 6) &&
        (PF2_MSI_CAP_MULTIMSGCAP_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute PF2_MSI_CAP_MULTIMSGCAP on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, PF2_MSI_CAP_MULTIMSGCAP_REG);
      attr_err = 1'b1;
    end

    if ((PF2_MSI_CAP_PERVECMASKCAP_REG != "FALSE") &&
        (PF2_MSI_CAP_PERVECMASKCAP_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF2_MSI_CAP_PERVECMASKCAP on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF2_MSI_CAP_PERVECMASKCAP_REG);
      attr_err = 1'b1;
    end

    if ((PF2_PB_CAP_SYSTEM_ALLOCATED_REG != "FALSE") &&
        (PF2_PB_CAP_SYSTEM_ALLOCATED_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF2_PB_CAP_SYSTEM_ALLOCATED on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF2_PB_CAP_SYSTEM_ALLOCATED_REG);
      attr_err = 1'b1;
    end

    if ((PF2_RBAR_CAP_ENABLE_REG != "FALSE") &&
        (PF2_RBAR_CAP_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF2_RBAR_CAP_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF2_RBAR_CAP_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((PF2_TPHR_CAP_DEV_SPECIFIC_MODE_REG != "TRUE") &&
        (PF2_TPHR_CAP_DEV_SPECIFIC_MODE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PF2_TPHR_CAP_DEV_SPECIFIC_MODE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PF2_TPHR_CAP_DEV_SPECIFIC_MODE_REG);
      attr_err = 1'b1;
    end

    if ((PF2_TPHR_CAP_ENABLE_REG != "FALSE") &&
        (PF2_TPHR_CAP_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF2_TPHR_CAP_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF2_TPHR_CAP_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((PF2_TPHR_CAP_INT_VEC_MODE_REG != "TRUE") &&
        (PF2_TPHR_CAP_INT_VEC_MODE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PF2_TPHR_CAP_INT_VEC_MODE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PF2_TPHR_CAP_INT_VEC_MODE_REG);
      attr_err = 1'b1;
    end

    if ((PF3_AER_CAP_ECRC_CHECK_CAPABLE_REG != "FALSE") &&
        (PF3_AER_CAP_ECRC_CHECK_CAPABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF3_AER_CAP_ECRC_CHECK_CAPABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF3_AER_CAP_ECRC_CHECK_CAPABLE_REG);
      attr_err = 1'b1;
    end

    if ((PF3_AER_CAP_ECRC_GEN_CAPABLE_REG != "FALSE") &&
        (PF3_AER_CAP_ECRC_GEN_CAPABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF3_AER_CAP_ECRC_GEN_CAPABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF3_AER_CAP_ECRC_GEN_CAPABLE_REG);
      attr_err = 1'b1;
    end

    if ((PF3_DPA_CAP_SUB_STATE_CONTROL_EN_REG != "TRUE") &&
        (PF3_DPA_CAP_SUB_STATE_CONTROL_EN_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PF3_DPA_CAP_SUB_STATE_CONTROL_EN on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PF3_DPA_CAP_SUB_STATE_CONTROL_EN_REG);
      attr_err = 1'b1;
    end

    if ((PF3_EXPANSION_ROM_ENABLE_REG != "FALSE") &&
        (PF3_EXPANSION_ROM_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF3_EXPANSION_ROM_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF3_EXPANSION_ROM_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((PF3_MSIX_CAP_PBA_BIR_REG != 0) &&
        (PF3_MSIX_CAP_PBA_BIR_REG != 1) &&
        (PF3_MSIX_CAP_PBA_BIR_REG != 2) &&
        (PF3_MSIX_CAP_PBA_BIR_REG != 3) &&
        (PF3_MSIX_CAP_PBA_BIR_REG != 4) &&
        (PF3_MSIX_CAP_PBA_BIR_REG != 5) &&
        (PF3_MSIX_CAP_PBA_BIR_REG != 6) &&
        (PF3_MSIX_CAP_PBA_BIR_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute PF3_MSIX_CAP_PBA_BIR on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, PF3_MSIX_CAP_PBA_BIR_REG);
      attr_err = 1'b1;
    end

    if ((PF3_MSIX_CAP_TABLE_BIR_REG != 0) &&
        (PF3_MSIX_CAP_TABLE_BIR_REG != 1) &&
        (PF3_MSIX_CAP_TABLE_BIR_REG != 2) &&
        (PF3_MSIX_CAP_TABLE_BIR_REG != 3) &&
        (PF3_MSIX_CAP_TABLE_BIR_REG != 4) &&
        (PF3_MSIX_CAP_TABLE_BIR_REG != 5) &&
        (PF3_MSIX_CAP_TABLE_BIR_REG != 6) &&
        (PF3_MSIX_CAP_TABLE_BIR_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute PF3_MSIX_CAP_TABLE_BIR on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, PF3_MSIX_CAP_TABLE_BIR_REG);
      attr_err = 1'b1;
    end

    if ((PF3_MSI_CAP_MULTIMSGCAP_REG != 0) &&
        (PF3_MSI_CAP_MULTIMSGCAP_REG != 1) &&
        (PF3_MSI_CAP_MULTIMSGCAP_REG != 2) &&
        (PF3_MSI_CAP_MULTIMSGCAP_REG != 3) &&
        (PF3_MSI_CAP_MULTIMSGCAP_REG != 4) &&
        (PF3_MSI_CAP_MULTIMSGCAP_REG != 5) &&
        (PF3_MSI_CAP_MULTIMSGCAP_REG != 6) &&
        (PF3_MSI_CAP_MULTIMSGCAP_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute PF3_MSI_CAP_MULTIMSGCAP on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, PF3_MSI_CAP_MULTIMSGCAP_REG);
      attr_err = 1'b1;
    end

    if ((PF3_MSI_CAP_PERVECMASKCAP_REG != "FALSE") &&
        (PF3_MSI_CAP_PERVECMASKCAP_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF3_MSI_CAP_PERVECMASKCAP on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF3_MSI_CAP_PERVECMASKCAP_REG);
      attr_err = 1'b1;
    end

    if ((PF3_PB_CAP_SYSTEM_ALLOCATED_REG != "FALSE") &&
        (PF3_PB_CAP_SYSTEM_ALLOCATED_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF3_PB_CAP_SYSTEM_ALLOCATED on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF3_PB_CAP_SYSTEM_ALLOCATED_REG);
      attr_err = 1'b1;
    end

    if ((PF3_RBAR_CAP_ENABLE_REG != "FALSE") &&
        (PF3_RBAR_CAP_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF3_RBAR_CAP_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF3_RBAR_CAP_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((PF3_TPHR_CAP_DEV_SPECIFIC_MODE_REG != "TRUE") &&
        (PF3_TPHR_CAP_DEV_SPECIFIC_MODE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PF3_TPHR_CAP_DEV_SPECIFIC_MODE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PF3_TPHR_CAP_DEV_SPECIFIC_MODE_REG);
      attr_err = 1'b1;
    end

    if ((PF3_TPHR_CAP_ENABLE_REG != "FALSE") &&
        (PF3_TPHR_CAP_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PF3_TPHR_CAP_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PF3_TPHR_CAP_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((PF3_TPHR_CAP_INT_VEC_MODE_REG != "TRUE") &&
        (PF3_TPHR_CAP_INT_VEC_MODE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PF3_TPHR_CAP_INT_VEC_MODE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PF3_TPHR_CAP_INT_VEC_MODE_REG);
      attr_err = 1'b1;
    end

    if ((PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3_REG != "FALSE") &&
        (PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3 on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3_REG);
      attr_err = 1'b1;
    end

    if ((PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2_REG != "FALSE") &&
        (PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2 on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2_REG);
      attr_err = 1'b1;
    end

    if ((PL_DISABLE_EI_INFER_IN_L0_REG != "FALSE") &&
        (PL_DISABLE_EI_INFER_IN_L0_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PL_DISABLE_EI_INFER_IN_L0 on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PL_DISABLE_EI_INFER_IN_L0_REG);
      attr_err = 1'b1;
    end

    if ((PL_DISABLE_GEN3_DC_BALANCE_REG != "FALSE") &&
        (PL_DISABLE_GEN3_DC_BALANCE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PL_DISABLE_GEN3_DC_BALANCE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PL_DISABLE_GEN3_DC_BALANCE_REG);
      attr_err = 1'b1;
    end

    if ((PL_DISABLE_GEN3_LFSR_UPDATE_ON_SKP_REG != "TRUE") &&
        (PL_DISABLE_GEN3_LFSR_UPDATE_ON_SKP_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PL_DISABLE_GEN3_LFSR_UPDATE_ON_SKP on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PL_DISABLE_GEN3_LFSR_UPDATE_ON_SKP_REG);
      attr_err = 1'b1;
    end

    if ((PL_DISABLE_RETRAIN_ON_FRAMING_ERROR_REG != "FALSE") &&
        (PL_DISABLE_RETRAIN_ON_FRAMING_ERROR_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PL_DISABLE_RETRAIN_ON_FRAMING_ERROR on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PL_DISABLE_RETRAIN_ON_FRAMING_ERROR_REG);
      attr_err = 1'b1;
    end

    if ((PL_DISABLE_SCRAMBLING_REG != "FALSE") &&
        (PL_DISABLE_SCRAMBLING_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PL_DISABLE_SCRAMBLING on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PL_DISABLE_SCRAMBLING_REG);
      attr_err = 1'b1;
    end

    if ((PL_DISABLE_SYNC_HEADER_FRAMING_ERROR_REG != "FALSE") &&
        (PL_DISABLE_SYNC_HEADER_FRAMING_ERROR_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PL_DISABLE_SYNC_HEADER_FRAMING_ERROR on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PL_DISABLE_SYNC_HEADER_FRAMING_ERROR_REG);
      attr_err = 1'b1;
    end

    if ((PL_DISABLE_UPCONFIG_CAPABLE_REG != "FALSE") &&
        (PL_DISABLE_UPCONFIG_CAPABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PL_DISABLE_UPCONFIG_CAPABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PL_DISABLE_UPCONFIG_CAPABLE_REG);
      attr_err = 1'b1;
    end

    if ((PL_EQ_ADAPT_DISABLE_COEFF_CHECK_REG != "FALSE") &&
        (PL_EQ_ADAPT_DISABLE_COEFF_CHECK_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PL_EQ_ADAPT_DISABLE_COEFF_CHECK on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PL_EQ_ADAPT_DISABLE_COEFF_CHECK_REG);
      attr_err = 1'b1;
    end

    if ((PL_EQ_ADAPT_DISABLE_PRESET_CHECK_REG != "FALSE") &&
        (PL_EQ_ADAPT_DISABLE_PRESET_CHECK_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PL_EQ_ADAPT_DISABLE_PRESET_CHECK on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PL_EQ_ADAPT_DISABLE_PRESET_CHECK_REG);
      attr_err = 1'b1;
    end

    if ((PL_EQ_BYPASS_PHASE23_REG != "FALSE") &&
        (PL_EQ_BYPASS_PHASE23_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PL_EQ_BYPASS_PHASE23 on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PL_EQ_BYPASS_PHASE23_REG);
      attr_err = 1'b1;
    end

    if ((PL_EQ_PHASE01_RX_ADAPT_REG != "FALSE") &&
        (PL_EQ_PHASE01_RX_ADAPT_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PL_EQ_PHASE01_RX_ADAPT on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PL_EQ_PHASE01_RX_ADAPT_REG);
      attr_err = 1'b1;
    end

    if ((PL_EQ_SHORT_ADAPT_PHASE_REG != "FALSE") &&
        (PL_EQ_SHORT_ADAPT_PHASE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PL_EQ_SHORT_ADAPT_PHASE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PL_EQ_SHORT_ADAPT_PHASE_REG);
      attr_err = 1'b1;
    end

    if ((PL_N_FTS_COMCLK_GEN1_REG < 0) || (PL_N_FTS_COMCLK_GEN1_REG > 255)) begin
      $display("Attribute Syntax Error : The attribute PL_N_FTS_COMCLK_GEN1 on %s instance %m is set to %d.  Legal values for this attribute are  0 to 255.", MODULE_NAME, PL_N_FTS_COMCLK_GEN1_REG);
      attr_err = 1'b1;
    end

    if ((PL_N_FTS_COMCLK_GEN2_REG < 0) || (PL_N_FTS_COMCLK_GEN2_REG > 255)) begin
      $display("Attribute Syntax Error : The attribute PL_N_FTS_COMCLK_GEN2 on %s instance %m is set to %d.  Legal values for this attribute are  0 to 255.", MODULE_NAME, PL_N_FTS_COMCLK_GEN2_REG);
      attr_err = 1'b1;
    end

    if ((PL_N_FTS_COMCLK_GEN3_REG < 0) || (PL_N_FTS_COMCLK_GEN3_REG > 255)) begin
      $display("Attribute Syntax Error : The attribute PL_N_FTS_COMCLK_GEN3 on %s instance %m is set to %d.  Legal values for this attribute are  0 to 255.", MODULE_NAME, PL_N_FTS_COMCLK_GEN3_REG);
      attr_err = 1'b1;
    end

    if ((PL_N_FTS_GEN1_REG < 0) || (PL_N_FTS_GEN1_REG > 255)) begin
      $display("Attribute Syntax Error : The attribute PL_N_FTS_GEN1 on %s instance %m is set to %d.  Legal values for this attribute are  0 to 255.", MODULE_NAME, PL_N_FTS_GEN1_REG);
      attr_err = 1'b1;
    end

    if ((PL_N_FTS_GEN2_REG < 0) || (PL_N_FTS_GEN2_REG > 255)) begin
      $display("Attribute Syntax Error : The attribute PL_N_FTS_GEN2 on %s instance %m is set to %d.  Legal values for this attribute are  0 to 255.", MODULE_NAME, PL_N_FTS_GEN2_REG);
      attr_err = 1'b1;
    end

    if ((PL_N_FTS_GEN3_REG < 0) || (PL_N_FTS_GEN3_REG > 255)) begin
      $display("Attribute Syntax Error : The attribute PL_N_FTS_GEN3 on %s instance %m is set to %d.  Legal values for this attribute are  0 to 255.", MODULE_NAME, PL_N_FTS_GEN3_REG);
      attr_err = 1'b1;
    end

    if ((PL_REPORT_ALL_PHY_ERRORS_REG != "TRUE") &&
        (PL_REPORT_ALL_PHY_ERRORS_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PL_REPORT_ALL_PHY_ERRORS on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PL_REPORT_ALL_PHY_ERRORS_REG);
      attr_err = 1'b1;
    end

    if ((PL_SIM_FAST_LINK_TRAINING_REG != "FALSE") &&
        (PL_SIM_FAST_LINK_TRAINING_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PL_SIM_FAST_LINK_TRAINING on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PL_SIM_FAST_LINK_TRAINING_REG);
      attr_err = 1'b1;
    end

    if ((PL_UPSTREAM_FACING_REG != "TRUE") &&
        (PL_UPSTREAM_FACING_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PL_UPSTREAM_FACING on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PL_UPSTREAM_FACING_REG);
      attr_err = 1'b1;
    end

    if ((PM_ENABLE_L23_ENTRY_REG != "FALSE") &&
        (PM_ENABLE_L23_ENTRY_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute PM_ENABLE_L23_ENTRY on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, PM_ENABLE_L23_ENTRY_REG);
      attr_err = 1'b1;
    end

    if ((PM_ENABLE_SLOT_POWER_CAPTURE_REG != "TRUE") &&
        (PM_ENABLE_SLOT_POWER_CAPTURE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute PM_ENABLE_SLOT_POWER_CAPTURE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, PM_ENABLE_SLOT_POWER_CAPTURE_REG);
      attr_err = 1'b1;
    end

    if ((SIM_VERSION_REG != "1.0") &&
        (SIM_VERSION_REG != "1.1") &&
        (SIM_VERSION_REG != "1.2") &&
        (SIM_VERSION_REG != "1.3") &&
        (SIM_VERSION_REG != "2.0") &&
        (SIM_VERSION_REG != "3.0") &&
        (SIM_VERSION_REG != "4.0")) begin
      $display("Attribute Syntax Error : The attribute SIM_VERSION on %s instance %m is set to %s.  Legal values for this attribute are 1.0, 1.1, 1.2, 1.3, 2.0, 3.0 or 4.0.", MODULE_NAME, SIM_VERSION_REG);
      attr_err = 1'b1;
    end

    if ((SPARE_BIT0_REG != 0) &&
        (SPARE_BIT0_REG != 1)) begin
      $display("Attribute Syntax Error : The attribute SPARE_BIT0 on %s instance %m is set to %d.  Legal values for this attribute are 0 to 1.", MODULE_NAME, SPARE_BIT0_REG);
      attr_err = 1'b1;
    end

    if ((SPARE_BIT1_REG != 0) &&
        (SPARE_BIT1_REG != 1)) begin
      $display("Attribute Syntax Error : The attribute SPARE_BIT1 on %s instance %m is set to %d.  Legal values for this attribute are 0 to 1.", MODULE_NAME, SPARE_BIT1_REG);
      attr_err = 1'b1;
    end

    if ((SPARE_BIT2_REG != 0) &&
        (SPARE_BIT2_REG != 1)) begin
      $display("Attribute Syntax Error : The attribute SPARE_BIT2 on %s instance %m is set to %d.  Legal values for this attribute are 0 to 1.", MODULE_NAME, SPARE_BIT2_REG);
      attr_err = 1'b1;
    end

    if ((SPARE_BIT3_REG != 0) &&
        (SPARE_BIT3_REG != 1)) begin
      $display("Attribute Syntax Error : The attribute SPARE_BIT3 on %s instance %m is set to %d.  Legal values for this attribute are 0 to 1.", MODULE_NAME, SPARE_BIT3_REG);
      attr_err = 1'b1;
    end

    if ((SPARE_BIT4_REG != 0) &&
        (SPARE_BIT4_REG != 1)) begin
      $display("Attribute Syntax Error : The attribute SPARE_BIT4 on %s instance %m is set to %d.  Legal values for this attribute are 0 to 1.", MODULE_NAME, SPARE_BIT4_REG);
      attr_err = 1'b1;
    end

    if ((SPARE_BIT5_REG != 0) &&
        (SPARE_BIT5_REG != 1)) begin
      $display("Attribute Syntax Error : The attribute SPARE_BIT5 on %s instance %m is set to %d.  Legal values for this attribute are 0 to 1.", MODULE_NAME, SPARE_BIT5_REG);
      attr_err = 1'b1;
    end

    if ((SPARE_BIT6_REG != 0) &&
        (SPARE_BIT6_REG != 1)) begin
      $display("Attribute Syntax Error : The attribute SPARE_BIT6 on %s instance %m is set to %d.  Legal values for this attribute are 0 to 1.", MODULE_NAME, SPARE_BIT6_REG);
      attr_err = 1'b1;
    end

    if ((SPARE_BIT7_REG != 0) &&
        (SPARE_BIT7_REG != 1)) begin
      $display("Attribute Syntax Error : The attribute SPARE_BIT7 on %s instance %m is set to %d.  Legal values for this attribute are 0 to 1.", MODULE_NAME, SPARE_BIT7_REG);
      attr_err = 1'b1;
    end

    if ((SPARE_BIT8_REG != 0) &&
        (SPARE_BIT8_REG != 1)) begin
      $display("Attribute Syntax Error : The attribute SPARE_BIT8 on %s instance %m is set to %d.  Legal values for this attribute are 0 to 1.", MODULE_NAME, SPARE_BIT8_REG);
      attr_err = 1'b1;
    end

    if ((SRIOV_CAP_ENABLE_REG != "FALSE") &&
        (SRIOV_CAP_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute SRIOV_CAP_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, SRIOV_CAP_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((TL_COMPLETION_RAM_SIZE_16K_REG != "TRUE") &&
        (TL_COMPLETION_RAM_SIZE_16K_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute TL_COMPLETION_RAM_SIZE_16K on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, TL_COMPLETION_RAM_SIZE_16K_REG);
      attr_err = 1'b1;
    end

    if ((TL_ENABLE_MESSAGE_RID_CHECK_ENABLE_REG != "TRUE") &&
        (TL_ENABLE_MESSAGE_RID_CHECK_ENABLE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute TL_ENABLE_MESSAGE_RID_CHECK_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, TL_ENABLE_MESSAGE_RID_CHECK_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE_REG != "FALSE") &&
        (TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE_REG != "FALSE") &&
        (TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((TL_LEGACY_MODE_ENABLE_REG != "FALSE") &&
        (TL_LEGACY_MODE_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute TL_LEGACY_MODE_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, TL_LEGACY_MODE_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((TL_TX_MUX_STRICT_PRIORITY_REG != "TRUE") &&
        (TL_TX_MUX_STRICT_PRIORITY_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute TL_TX_MUX_STRICT_PRIORITY on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, TL_TX_MUX_STRICT_PRIORITY_REG);
      attr_err = 1'b1;
    end

    if ((TWO_LAYER_MODE_DLCMSM_ENABLE_REG != "TRUE") &&
        (TWO_LAYER_MODE_DLCMSM_ENABLE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute TWO_LAYER_MODE_DLCMSM_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, TWO_LAYER_MODE_DLCMSM_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((TWO_LAYER_MODE_ENABLE_REG != "FALSE") &&
        (TWO_LAYER_MODE_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute TWO_LAYER_MODE_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, TWO_LAYER_MODE_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((TWO_LAYER_MODE_WIDTH_256_REG != "TRUE") &&
        (TWO_LAYER_MODE_WIDTH_256_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute TWO_LAYER_MODE_WIDTH_256 on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, TWO_LAYER_MODE_WIDTH_256_REG);
      attr_err = 1'b1;
    end

    if ((VF0_MSIX_CAP_PBA_BIR_REG != 0) &&
        (VF0_MSIX_CAP_PBA_BIR_REG != 1) &&
        (VF0_MSIX_CAP_PBA_BIR_REG != 2) &&
        (VF0_MSIX_CAP_PBA_BIR_REG != 3) &&
        (VF0_MSIX_CAP_PBA_BIR_REG != 4) &&
        (VF0_MSIX_CAP_PBA_BIR_REG != 5) &&
        (VF0_MSIX_CAP_PBA_BIR_REG != 6) &&
        (VF0_MSIX_CAP_PBA_BIR_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute VF0_MSIX_CAP_PBA_BIR on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, VF0_MSIX_CAP_PBA_BIR_REG);
      attr_err = 1'b1;
    end

    if ((VF0_MSIX_CAP_TABLE_BIR_REG != 0) &&
        (VF0_MSIX_CAP_TABLE_BIR_REG != 1) &&
        (VF0_MSIX_CAP_TABLE_BIR_REG != 2) &&
        (VF0_MSIX_CAP_TABLE_BIR_REG != 3) &&
        (VF0_MSIX_CAP_TABLE_BIR_REG != 4) &&
        (VF0_MSIX_CAP_TABLE_BIR_REG != 5) &&
        (VF0_MSIX_CAP_TABLE_BIR_REG != 6) &&
        (VF0_MSIX_CAP_TABLE_BIR_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute VF0_MSIX_CAP_TABLE_BIR on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, VF0_MSIX_CAP_TABLE_BIR_REG);
      attr_err = 1'b1;
    end

    if ((VF0_MSI_CAP_MULTIMSGCAP_REG != 0) &&
        (VF0_MSI_CAP_MULTIMSGCAP_REG != 1) &&
        (VF0_MSI_CAP_MULTIMSGCAP_REG != 2) &&
        (VF0_MSI_CAP_MULTIMSGCAP_REG != 3) &&
        (VF0_MSI_CAP_MULTIMSGCAP_REG != 4) &&
        (VF0_MSI_CAP_MULTIMSGCAP_REG != 5) &&
        (VF0_MSI_CAP_MULTIMSGCAP_REG != 6) &&
        (VF0_MSI_CAP_MULTIMSGCAP_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute VF0_MSI_CAP_MULTIMSGCAP on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, VF0_MSI_CAP_MULTIMSGCAP_REG);
      attr_err = 1'b1;
    end

    if ((VF0_TPHR_CAP_DEV_SPECIFIC_MODE_REG != "TRUE") &&
        (VF0_TPHR_CAP_DEV_SPECIFIC_MODE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute VF0_TPHR_CAP_DEV_SPECIFIC_MODE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, VF0_TPHR_CAP_DEV_SPECIFIC_MODE_REG);
      attr_err = 1'b1;
    end

    if ((VF0_TPHR_CAP_ENABLE_REG != "FALSE") &&
        (VF0_TPHR_CAP_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute VF0_TPHR_CAP_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, VF0_TPHR_CAP_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((VF0_TPHR_CAP_INT_VEC_MODE_REG != "TRUE") &&
        (VF0_TPHR_CAP_INT_VEC_MODE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute VF0_TPHR_CAP_INT_VEC_MODE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, VF0_TPHR_CAP_INT_VEC_MODE_REG);
      attr_err = 1'b1;
    end

    if ((VF1_MSIX_CAP_PBA_BIR_REG != 0) &&
        (VF1_MSIX_CAP_PBA_BIR_REG != 1) &&
        (VF1_MSIX_CAP_PBA_BIR_REG != 2) &&
        (VF1_MSIX_CAP_PBA_BIR_REG != 3) &&
        (VF1_MSIX_CAP_PBA_BIR_REG != 4) &&
        (VF1_MSIX_CAP_PBA_BIR_REG != 5) &&
        (VF1_MSIX_CAP_PBA_BIR_REG != 6) &&
        (VF1_MSIX_CAP_PBA_BIR_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute VF1_MSIX_CAP_PBA_BIR on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, VF1_MSIX_CAP_PBA_BIR_REG);
      attr_err = 1'b1;
    end

    if ((VF1_MSIX_CAP_TABLE_BIR_REG != 0) &&
        (VF1_MSIX_CAP_TABLE_BIR_REG != 1) &&
        (VF1_MSIX_CAP_TABLE_BIR_REG != 2) &&
        (VF1_MSIX_CAP_TABLE_BIR_REG != 3) &&
        (VF1_MSIX_CAP_TABLE_BIR_REG != 4) &&
        (VF1_MSIX_CAP_TABLE_BIR_REG != 5) &&
        (VF1_MSIX_CAP_TABLE_BIR_REG != 6) &&
        (VF1_MSIX_CAP_TABLE_BIR_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute VF1_MSIX_CAP_TABLE_BIR on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, VF1_MSIX_CAP_TABLE_BIR_REG);
      attr_err = 1'b1;
    end

    if ((VF1_MSI_CAP_MULTIMSGCAP_REG != 0) &&
        (VF1_MSI_CAP_MULTIMSGCAP_REG != 1) &&
        (VF1_MSI_CAP_MULTIMSGCAP_REG != 2) &&
        (VF1_MSI_CAP_MULTIMSGCAP_REG != 3) &&
        (VF1_MSI_CAP_MULTIMSGCAP_REG != 4) &&
        (VF1_MSI_CAP_MULTIMSGCAP_REG != 5) &&
        (VF1_MSI_CAP_MULTIMSGCAP_REG != 6) &&
        (VF1_MSI_CAP_MULTIMSGCAP_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute VF1_MSI_CAP_MULTIMSGCAP on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, VF1_MSI_CAP_MULTIMSGCAP_REG);
      attr_err = 1'b1;
    end

    if ((VF1_TPHR_CAP_DEV_SPECIFIC_MODE_REG != "TRUE") &&
        (VF1_TPHR_CAP_DEV_SPECIFIC_MODE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute VF1_TPHR_CAP_DEV_SPECIFIC_MODE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, VF1_TPHR_CAP_DEV_SPECIFIC_MODE_REG);
      attr_err = 1'b1;
    end

    if ((VF1_TPHR_CAP_ENABLE_REG != "FALSE") &&
        (VF1_TPHR_CAP_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute VF1_TPHR_CAP_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, VF1_TPHR_CAP_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((VF1_TPHR_CAP_INT_VEC_MODE_REG != "TRUE") &&
        (VF1_TPHR_CAP_INT_VEC_MODE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute VF1_TPHR_CAP_INT_VEC_MODE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, VF1_TPHR_CAP_INT_VEC_MODE_REG);
      attr_err = 1'b1;
    end

    if ((VF2_MSIX_CAP_PBA_BIR_REG != 0) &&
        (VF2_MSIX_CAP_PBA_BIR_REG != 1) &&
        (VF2_MSIX_CAP_PBA_BIR_REG != 2) &&
        (VF2_MSIX_CAP_PBA_BIR_REG != 3) &&
        (VF2_MSIX_CAP_PBA_BIR_REG != 4) &&
        (VF2_MSIX_CAP_PBA_BIR_REG != 5) &&
        (VF2_MSIX_CAP_PBA_BIR_REG != 6) &&
        (VF2_MSIX_CAP_PBA_BIR_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute VF2_MSIX_CAP_PBA_BIR on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, VF2_MSIX_CAP_PBA_BIR_REG);
      attr_err = 1'b1;
    end

    if ((VF2_MSIX_CAP_TABLE_BIR_REG != 0) &&
        (VF2_MSIX_CAP_TABLE_BIR_REG != 1) &&
        (VF2_MSIX_CAP_TABLE_BIR_REG != 2) &&
        (VF2_MSIX_CAP_TABLE_BIR_REG != 3) &&
        (VF2_MSIX_CAP_TABLE_BIR_REG != 4) &&
        (VF2_MSIX_CAP_TABLE_BIR_REG != 5) &&
        (VF2_MSIX_CAP_TABLE_BIR_REG != 6) &&
        (VF2_MSIX_CAP_TABLE_BIR_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute VF2_MSIX_CAP_TABLE_BIR on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, VF2_MSIX_CAP_TABLE_BIR_REG);
      attr_err = 1'b1;
    end

    if ((VF2_MSI_CAP_MULTIMSGCAP_REG != 0) &&
        (VF2_MSI_CAP_MULTIMSGCAP_REG != 1) &&
        (VF2_MSI_CAP_MULTIMSGCAP_REG != 2) &&
        (VF2_MSI_CAP_MULTIMSGCAP_REG != 3) &&
        (VF2_MSI_CAP_MULTIMSGCAP_REG != 4) &&
        (VF2_MSI_CAP_MULTIMSGCAP_REG != 5) &&
        (VF2_MSI_CAP_MULTIMSGCAP_REG != 6) &&
        (VF2_MSI_CAP_MULTIMSGCAP_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute VF2_MSI_CAP_MULTIMSGCAP on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, VF2_MSI_CAP_MULTIMSGCAP_REG);
      attr_err = 1'b1;
    end

    if ((VF2_TPHR_CAP_DEV_SPECIFIC_MODE_REG != "TRUE") &&
        (VF2_TPHR_CAP_DEV_SPECIFIC_MODE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute VF2_TPHR_CAP_DEV_SPECIFIC_MODE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, VF2_TPHR_CAP_DEV_SPECIFIC_MODE_REG);
      attr_err = 1'b1;
    end

    if ((VF2_TPHR_CAP_ENABLE_REG != "FALSE") &&
        (VF2_TPHR_CAP_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute VF2_TPHR_CAP_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, VF2_TPHR_CAP_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((VF2_TPHR_CAP_INT_VEC_MODE_REG != "TRUE") &&
        (VF2_TPHR_CAP_INT_VEC_MODE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute VF2_TPHR_CAP_INT_VEC_MODE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, VF2_TPHR_CAP_INT_VEC_MODE_REG);
      attr_err = 1'b1;
    end

    if ((VF3_MSIX_CAP_PBA_BIR_REG != 0) &&
        (VF3_MSIX_CAP_PBA_BIR_REG != 1) &&
        (VF3_MSIX_CAP_PBA_BIR_REG != 2) &&
        (VF3_MSIX_CAP_PBA_BIR_REG != 3) &&
        (VF3_MSIX_CAP_PBA_BIR_REG != 4) &&
        (VF3_MSIX_CAP_PBA_BIR_REG != 5) &&
        (VF3_MSIX_CAP_PBA_BIR_REG != 6) &&
        (VF3_MSIX_CAP_PBA_BIR_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute VF3_MSIX_CAP_PBA_BIR on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, VF3_MSIX_CAP_PBA_BIR_REG);
      attr_err = 1'b1;
    end

    if ((VF3_MSIX_CAP_TABLE_BIR_REG != 0) &&
        (VF3_MSIX_CAP_TABLE_BIR_REG != 1) &&
        (VF3_MSIX_CAP_TABLE_BIR_REG != 2) &&
        (VF3_MSIX_CAP_TABLE_BIR_REG != 3) &&
        (VF3_MSIX_CAP_TABLE_BIR_REG != 4) &&
        (VF3_MSIX_CAP_TABLE_BIR_REG != 5) &&
        (VF3_MSIX_CAP_TABLE_BIR_REG != 6) &&
        (VF3_MSIX_CAP_TABLE_BIR_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute VF3_MSIX_CAP_TABLE_BIR on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, VF3_MSIX_CAP_TABLE_BIR_REG);
      attr_err = 1'b1;
    end

    if ((VF3_MSI_CAP_MULTIMSGCAP_REG != 0) &&
        (VF3_MSI_CAP_MULTIMSGCAP_REG != 1) &&
        (VF3_MSI_CAP_MULTIMSGCAP_REG != 2) &&
        (VF3_MSI_CAP_MULTIMSGCAP_REG != 3) &&
        (VF3_MSI_CAP_MULTIMSGCAP_REG != 4) &&
        (VF3_MSI_CAP_MULTIMSGCAP_REG != 5) &&
        (VF3_MSI_CAP_MULTIMSGCAP_REG != 6) &&
        (VF3_MSI_CAP_MULTIMSGCAP_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute VF3_MSI_CAP_MULTIMSGCAP on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, VF3_MSI_CAP_MULTIMSGCAP_REG);
      attr_err = 1'b1;
    end

    if ((VF3_TPHR_CAP_DEV_SPECIFIC_MODE_REG != "TRUE") &&
        (VF3_TPHR_CAP_DEV_SPECIFIC_MODE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute VF3_TPHR_CAP_DEV_SPECIFIC_MODE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, VF3_TPHR_CAP_DEV_SPECIFIC_MODE_REG);
      attr_err = 1'b1;
    end

    if ((VF3_TPHR_CAP_ENABLE_REG != "FALSE") &&
        (VF3_TPHR_CAP_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute VF3_TPHR_CAP_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, VF3_TPHR_CAP_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((VF3_TPHR_CAP_INT_VEC_MODE_REG != "TRUE") &&
        (VF3_TPHR_CAP_INT_VEC_MODE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute VF3_TPHR_CAP_INT_VEC_MODE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, VF3_TPHR_CAP_INT_VEC_MODE_REG);
      attr_err = 1'b1;
    end

    if ((VF4_MSIX_CAP_PBA_BIR_REG != 0) &&
        (VF4_MSIX_CAP_PBA_BIR_REG != 1) &&
        (VF4_MSIX_CAP_PBA_BIR_REG != 2) &&
        (VF4_MSIX_CAP_PBA_BIR_REG != 3) &&
        (VF4_MSIX_CAP_PBA_BIR_REG != 4) &&
        (VF4_MSIX_CAP_PBA_BIR_REG != 5) &&
        (VF4_MSIX_CAP_PBA_BIR_REG != 6) &&
        (VF4_MSIX_CAP_PBA_BIR_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute VF4_MSIX_CAP_PBA_BIR on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, VF4_MSIX_CAP_PBA_BIR_REG);
      attr_err = 1'b1;
    end

    if ((VF4_MSIX_CAP_TABLE_BIR_REG != 0) &&
        (VF4_MSIX_CAP_TABLE_BIR_REG != 1) &&
        (VF4_MSIX_CAP_TABLE_BIR_REG != 2) &&
        (VF4_MSIX_CAP_TABLE_BIR_REG != 3) &&
        (VF4_MSIX_CAP_TABLE_BIR_REG != 4) &&
        (VF4_MSIX_CAP_TABLE_BIR_REG != 5) &&
        (VF4_MSIX_CAP_TABLE_BIR_REG != 6) &&
        (VF4_MSIX_CAP_TABLE_BIR_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute VF4_MSIX_CAP_TABLE_BIR on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, VF4_MSIX_CAP_TABLE_BIR_REG);
      attr_err = 1'b1;
    end

    if ((VF4_MSI_CAP_MULTIMSGCAP_REG != 0) &&
        (VF4_MSI_CAP_MULTIMSGCAP_REG != 1) &&
        (VF4_MSI_CAP_MULTIMSGCAP_REG != 2) &&
        (VF4_MSI_CAP_MULTIMSGCAP_REG != 3) &&
        (VF4_MSI_CAP_MULTIMSGCAP_REG != 4) &&
        (VF4_MSI_CAP_MULTIMSGCAP_REG != 5) &&
        (VF4_MSI_CAP_MULTIMSGCAP_REG != 6) &&
        (VF4_MSI_CAP_MULTIMSGCAP_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute VF4_MSI_CAP_MULTIMSGCAP on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, VF4_MSI_CAP_MULTIMSGCAP_REG);
      attr_err = 1'b1;
    end

    if ((VF4_TPHR_CAP_DEV_SPECIFIC_MODE_REG != "TRUE") &&
        (VF4_TPHR_CAP_DEV_SPECIFIC_MODE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute VF4_TPHR_CAP_DEV_SPECIFIC_MODE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, VF4_TPHR_CAP_DEV_SPECIFIC_MODE_REG);
      attr_err = 1'b1;
    end

    if ((VF4_TPHR_CAP_ENABLE_REG != "FALSE") &&
        (VF4_TPHR_CAP_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute VF4_TPHR_CAP_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, VF4_TPHR_CAP_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((VF4_TPHR_CAP_INT_VEC_MODE_REG != "TRUE") &&
        (VF4_TPHR_CAP_INT_VEC_MODE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute VF4_TPHR_CAP_INT_VEC_MODE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, VF4_TPHR_CAP_INT_VEC_MODE_REG);
      attr_err = 1'b1;
    end

    if ((VF5_MSIX_CAP_PBA_BIR_REG != 0) &&
        (VF5_MSIX_CAP_PBA_BIR_REG != 1) &&
        (VF5_MSIX_CAP_PBA_BIR_REG != 2) &&
        (VF5_MSIX_CAP_PBA_BIR_REG != 3) &&
        (VF5_MSIX_CAP_PBA_BIR_REG != 4) &&
        (VF5_MSIX_CAP_PBA_BIR_REG != 5) &&
        (VF5_MSIX_CAP_PBA_BIR_REG != 6) &&
        (VF5_MSIX_CAP_PBA_BIR_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute VF5_MSIX_CAP_PBA_BIR on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, VF5_MSIX_CAP_PBA_BIR_REG);
      attr_err = 1'b1;
    end

    if ((VF5_MSIX_CAP_TABLE_BIR_REG != 0) &&
        (VF5_MSIX_CAP_TABLE_BIR_REG != 1) &&
        (VF5_MSIX_CAP_TABLE_BIR_REG != 2) &&
        (VF5_MSIX_CAP_TABLE_BIR_REG != 3) &&
        (VF5_MSIX_CAP_TABLE_BIR_REG != 4) &&
        (VF5_MSIX_CAP_TABLE_BIR_REG != 5) &&
        (VF5_MSIX_CAP_TABLE_BIR_REG != 6) &&
        (VF5_MSIX_CAP_TABLE_BIR_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute VF5_MSIX_CAP_TABLE_BIR on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, VF5_MSIX_CAP_TABLE_BIR_REG);
      attr_err = 1'b1;
    end

    if ((VF5_MSI_CAP_MULTIMSGCAP_REG != 0) &&
        (VF5_MSI_CAP_MULTIMSGCAP_REG != 1) &&
        (VF5_MSI_CAP_MULTIMSGCAP_REG != 2) &&
        (VF5_MSI_CAP_MULTIMSGCAP_REG != 3) &&
        (VF5_MSI_CAP_MULTIMSGCAP_REG != 4) &&
        (VF5_MSI_CAP_MULTIMSGCAP_REG != 5) &&
        (VF5_MSI_CAP_MULTIMSGCAP_REG != 6) &&
        (VF5_MSI_CAP_MULTIMSGCAP_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute VF5_MSI_CAP_MULTIMSGCAP on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, VF5_MSI_CAP_MULTIMSGCAP_REG);
      attr_err = 1'b1;
    end

    if ((VF5_TPHR_CAP_DEV_SPECIFIC_MODE_REG != "TRUE") &&
        (VF5_TPHR_CAP_DEV_SPECIFIC_MODE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute VF5_TPHR_CAP_DEV_SPECIFIC_MODE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, VF5_TPHR_CAP_DEV_SPECIFIC_MODE_REG);
      attr_err = 1'b1;
    end

    if ((VF5_TPHR_CAP_ENABLE_REG != "FALSE") &&
        (VF5_TPHR_CAP_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute VF5_TPHR_CAP_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, VF5_TPHR_CAP_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((VF5_TPHR_CAP_INT_VEC_MODE_REG != "TRUE") &&
        (VF5_TPHR_CAP_INT_VEC_MODE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute VF5_TPHR_CAP_INT_VEC_MODE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, VF5_TPHR_CAP_INT_VEC_MODE_REG);
      attr_err = 1'b1;
    end

    if ((VF6_MSIX_CAP_PBA_BIR_REG != 0) &&
        (VF6_MSIX_CAP_PBA_BIR_REG != 1) &&
        (VF6_MSIX_CAP_PBA_BIR_REG != 2) &&
        (VF6_MSIX_CAP_PBA_BIR_REG != 3) &&
        (VF6_MSIX_CAP_PBA_BIR_REG != 4) &&
        (VF6_MSIX_CAP_PBA_BIR_REG != 5) &&
        (VF6_MSIX_CAP_PBA_BIR_REG != 6) &&
        (VF6_MSIX_CAP_PBA_BIR_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute VF6_MSIX_CAP_PBA_BIR on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, VF6_MSIX_CAP_PBA_BIR_REG);
      attr_err = 1'b1;
    end

    if ((VF6_MSIX_CAP_TABLE_BIR_REG != 0) &&
        (VF6_MSIX_CAP_TABLE_BIR_REG != 1) &&
        (VF6_MSIX_CAP_TABLE_BIR_REG != 2) &&
        (VF6_MSIX_CAP_TABLE_BIR_REG != 3) &&
        (VF6_MSIX_CAP_TABLE_BIR_REG != 4) &&
        (VF6_MSIX_CAP_TABLE_BIR_REG != 5) &&
        (VF6_MSIX_CAP_TABLE_BIR_REG != 6) &&
        (VF6_MSIX_CAP_TABLE_BIR_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute VF6_MSIX_CAP_TABLE_BIR on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, VF6_MSIX_CAP_TABLE_BIR_REG);
      attr_err = 1'b1;
    end

    if ((VF6_MSI_CAP_MULTIMSGCAP_REG != 0) &&
        (VF6_MSI_CAP_MULTIMSGCAP_REG != 1) &&
        (VF6_MSI_CAP_MULTIMSGCAP_REG != 2) &&
        (VF6_MSI_CAP_MULTIMSGCAP_REG != 3) &&
        (VF6_MSI_CAP_MULTIMSGCAP_REG != 4) &&
        (VF6_MSI_CAP_MULTIMSGCAP_REG != 5) &&
        (VF6_MSI_CAP_MULTIMSGCAP_REG != 6) &&
        (VF6_MSI_CAP_MULTIMSGCAP_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute VF6_MSI_CAP_MULTIMSGCAP on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, VF6_MSI_CAP_MULTIMSGCAP_REG);
      attr_err = 1'b1;
    end

    if ((VF6_TPHR_CAP_DEV_SPECIFIC_MODE_REG != "TRUE") &&
        (VF6_TPHR_CAP_DEV_SPECIFIC_MODE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute VF6_TPHR_CAP_DEV_SPECIFIC_MODE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, VF6_TPHR_CAP_DEV_SPECIFIC_MODE_REG);
      attr_err = 1'b1;
    end

    if ((VF6_TPHR_CAP_ENABLE_REG != "FALSE") &&
        (VF6_TPHR_CAP_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute VF6_TPHR_CAP_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, VF6_TPHR_CAP_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((VF6_TPHR_CAP_INT_VEC_MODE_REG != "TRUE") &&
        (VF6_TPHR_CAP_INT_VEC_MODE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute VF6_TPHR_CAP_INT_VEC_MODE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, VF6_TPHR_CAP_INT_VEC_MODE_REG);
      attr_err = 1'b1;
    end

    if ((VF7_MSIX_CAP_PBA_BIR_REG != 0) &&
        (VF7_MSIX_CAP_PBA_BIR_REG != 1) &&
        (VF7_MSIX_CAP_PBA_BIR_REG != 2) &&
        (VF7_MSIX_CAP_PBA_BIR_REG != 3) &&
        (VF7_MSIX_CAP_PBA_BIR_REG != 4) &&
        (VF7_MSIX_CAP_PBA_BIR_REG != 5) &&
        (VF7_MSIX_CAP_PBA_BIR_REG != 6) &&
        (VF7_MSIX_CAP_PBA_BIR_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute VF7_MSIX_CAP_PBA_BIR on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, VF7_MSIX_CAP_PBA_BIR_REG);
      attr_err = 1'b1;
    end

    if ((VF7_MSIX_CAP_TABLE_BIR_REG != 0) &&
        (VF7_MSIX_CAP_TABLE_BIR_REG != 1) &&
        (VF7_MSIX_CAP_TABLE_BIR_REG != 2) &&
        (VF7_MSIX_CAP_TABLE_BIR_REG != 3) &&
        (VF7_MSIX_CAP_TABLE_BIR_REG != 4) &&
        (VF7_MSIX_CAP_TABLE_BIR_REG != 5) &&
        (VF7_MSIX_CAP_TABLE_BIR_REG != 6) &&
        (VF7_MSIX_CAP_TABLE_BIR_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute VF7_MSIX_CAP_TABLE_BIR on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, VF7_MSIX_CAP_TABLE_BIR_REG);
      attr_err = 1'b1;
    end

    if ((VF7_MSI_CAP_MULTIMSGCAP_REG != 0) &&
        (VF7_MSI_CAP_MULTIMSGCAP_REG != 1) &&
        (VF7_MSI_CAP_MULTIMSGCAP_REG != 2) &&
        (VF7_MSI_CAP_MULTIMSGCAP_REG != 3) &&
        (VF7_MSI_CAP_MULTIMSGCAP_REG != 4) &&
        (VF7_MSI_CAP_MULTIMSGCAP_REG != 5) &&
        (VF7_MSI_CAP_MULTIMSGCAP_REG != 6) &&
        (VF7_MSI_CAP_MULTIMSGCAP_REG != 7)) begin
      $display("Attribute Syntax Error : The attribute VF7_MSI_CAP_MULTIMSGCAP on %s instance %m is set to %d.  Legal values for this attribute are 0 to 7.", MODULE_NAME, VF7_MSI_CAP_MULTIMSGCAP_REG);
      attr_err = 1'b1;
    end

    if ((VF7_TPHR_CAP_DEV_SPECIFIC_MODE_REG != "TRUE") &&
        (VF7_TPHR_CAP_DEV_SPECIFIC_MODE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute VF7_TPHR_CAP_DEV_SPECIFIC_MODE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, VF7_TPHR_CAP_DEV_SPECIFIC_MODE_REG);
      attr_err = 1'b1;
    end

    if ((VF7_TPHR_CAP_ENABLE_REG != "FALSE") &&
        (VF7_TPHR_CAP_ENABLE_REG != "TRUE")) begin
      $display("Attribute Syntax Error : The attribute VF7_TPHR_CAP_ENABLE on %s instance %m is set to %s.  Legal values for this attribute are FALSE or TRUE.", MODULE_NAME, VF7_TPHR_CAP_ENABLE_REG);
      attr_err = 1'b1;
    end

    if ((VF7_TPHR_CAP_INT_VEC_MODE_REG != "TRUE") &&
        (VF7_TPHR_CAP_INT_VEC_MODE_REG != "FALSE")) begin
      $display("Attribute Syntax Error : The attribute VF7_TPHR_CAP_INT_VEC_MODE on %s instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", MODULE_NAME, VF7_TPHR_CAP_INT_VEC_MODE_REG);
      attr_err = 1'b1;
    end

  if (attr_err == 1'b1) $finish;
  end

  assign XILUNCONNCLK_in = 951'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111; // tie off

  assign PMVDIVIDE_in = 2'b11; // tie off
  assign PMVENABLEN_in = 1'b1; // tie off
  assign PMVSELECT_in = 3'b111; // tie off
  assign SCANENABLEN_in = 1'b1; // tie off
  assign SCANIN_in = 96'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111; // tie off
  assign SCANMODEN_in = 1'b1; // tie off
  assign XILUNCONNBYP_in = 1920'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111; // tie off
  assign XILUNCONNIN_in = 3189'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111; // tie off

  SIP_PCIE_3_1 # (
.MCAP_ENABLE_PAR (MCAP_ENABLE),
.SIM_JTAG_IDCODE (SIM_JTAG_IDCODE)
)  SIP_PCIE_3_1_INST (
     
    .ARI_CAP_ENABLE (ARI_CAP_ENABLE_REG),
    .AXISTEN_IF_CC_ALIGNMENT_MODE (AXISTEN_IF_CC_ALIGNMENT_MODE_REG),
    .AXISTEN_IF_CC_PARITY_CHK (AXISTEN_IF_CC_PARITY_CHK_REG),
    .AXISTEN_IF_CQ_ALIGNMENT_MODE (AXISTEN_IF_CQ_ALIGNMENT_MODE_REG),
    .AXISTEN_IF_ENABLE_CLIENT_TAG (AXISTEN_IF_ENABLE_CLIENT_TAG_REG),
    .AXISTEN_IF_ENABLE_MSG_ROUTE (AXISTEN_IF_ENABLE_MSG_ROUTE_REG),
    .AXISTEN_IF_ENABLE_RX_MSG_INTFC (AXISTEN_IF_ENABLE_RX_MSG_INTFC_REG),
    .AXISTEN_IF_RC_ALIGNMENT_MODE (AXISTEN_IF_RC_ALIGNMENT_MODE_REG),
    .AXISTEN_IF_RC_STRADDLE (AXISTEN_IF_RC_STRADDLE_REG),
    .AXISTEN_IF_RQ_ALIGNMENT_MODE (AXISTEN_IF_RQ_ALIGNMENT_MODE_REG),
    .AXISTEN_IF_RQ_PARITY_CHK (AXISTEN_IF_RQ_PARITY_CHK_REG),
    .AXISTEN_IF_WIDTH (AXISTEN_IF_WIDTH_REG),
    .CRM_CORE_CLK_FREQ_500 (CRM_CORE_CLK_FREQ_500_REG),
    .CRM_USER_CLK_FREQ (CRM_USER_CLK_FREQ_REG),
    .DEBUG_CFG_LOCAL_MGMT_REG_ACCESS_OVERRIDE (DEBUG_CFG_LOCAL_MGMT_REG_ACCESS_OVERRIDE_REG),
    .DEBUG_PL_DISABLE_EI_INFER_IN_L0 (DEBUG_PL_DISABLE_EI_INFER_IN_L0_REG),
    .DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS (DEBUG_TL_DISABLE_RX_TLP_ORDER_CHECKS_REG),
    .DNSTREAM_LINK_NUM (DNSTREAM_LINK_NUM_REG),
    .LL_ACK_TIMEOUT (LL_ACK_TIMEOUT_REG),
    .LL_ACK_TIMEOUT_EN (LL_ACK_TIMEOUT_EN_REG),
    .LL_ACK_TIMEOUT_FUNC (LL_ACK_TIMEOUT_FUNC_REG),
    .LL_CPL_FC_UPDATE_TIMER (LL_CPL_FC_UPDATE_TIMER_REG),
    .LL_CPL_FC_UPDATE_TIMER_OVERRIDE (LL_CPL_FC_UPDATE_TIMER_OVERRIDE_REG),
    .LL_FC_UPDATE_TIMER (LL_FC_UPDATE_TIMER_REG),
    .LL_FC_UPDATE_TIMER_OVERRIDE (LL_FC_UPDATE_TIMER_OVERRIDE_REG),
    .LL_NP_FC_UPDATE_TIMER (LL_NP_FC_UPDATE_TIMER_REG),
    .LL_NP_FC_UPDATE_TIMER_OVERRIDE (LL_NP_FC_UPDATE_TIMER_OVERRIDE_REG),
    .LL_P_FC_UPDATE_TIMER (LL_P_FC_UPDATE_TIMER_REG),
    .LL_P_FC_UPDATE_TIMER_OVERRIDE (LL_P_FC_UPDATE_TIMER_OVERRIDE_REG),
    .LL_REPLAY_TIMEOUT (LL_REPLAY_TIMEOUT_REG),
    .LL_REPLAY_TIMEOUT_EN (LL_REPLAY_TIMEOUT_EN_REG),
    .LL_REPLAY_TIMEOUT_FUNC (LL_REPLAY_TIMEOUT_FUNC_REG),
    .LTR_TX_MESSAGE_MINIMUM_INTERVAL (LTR_TX_MESSAGE_MINIMUM_INTERVAL_REG),
    .LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE (LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE_REG),
    .LTR_TX_MESSAGE_ON_LTR_ENABLE (LTR_TX_MESSAGE_ON_LTR_ENABLE_REG),
    .MCAP_CAP_NEXTPTR (MCAP_CAP_NEXTPTR_REG),
    .MCAP_CONFIGURE_OVERRIDE (MCAP_CONFIGURE_OVERRIDE_REG),
    .MCAP_ENABLE (MCAP_ENABLE_REG),
    .MCAP_EOS_DESIGN_SWITCH (MCAP_EOS_DESIGN_SWITCH_REG),
    .MCAP_FPGA_BITSTREAM_VERSION (MCAP_FPGA_BITSTREAM_VERSION_REG),
    .MCAP_GATE_IO_ENABLE_DESIGN_SWITCH (MCAP_GATE_IO_ENABLE_DESIGN_SWITCH_REG),
    .MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH (MCAP_GATE_MEM_ENABLE_DESIGN_SWITCH_REG),
    .MCAP_INPUT_GATE_DESIGN_SWITCH (MCAP_INPUT_GATE_DESIGN_SWITCH_REG),
    .MCAP_INTERRUPT_ON_MCAP_EOS (MCAP_INTERRUPT_ON_MCAP_EOS_REG),
    .MCAP_INTERRUPT_ON_MCAP_ERROR (MCAP_INTERRUPT_ON_MCAP_ERROR_REG),
    .MCAP_VSEC_ID (MCAP_VSEC_ID_REG),
    .MCAP_VSEC_LEN (MCAP_VSEC_LEN_REG),
    .MCAP_VSEC_REV (MCAP_VSEC_REV_REG),
    .PF0_AER_CAP_ECRC_CHECK_CAPABLE (PF0_AER_CAP_ECRC_CHECK_CAPABLE_REG),
    .PF0_AER_CAP_ECRC_GEN_CAPABLE (PF0_AER_CAP_ECRC_GEN_CAPABLE_REG),
    .PF0_AER_CAP_NEXTPTR (PF0_AER_CAP_NEXTPTR_REG),
    .PF0_ARI_CAP_NEXTPTR (PF0_ARI_CAP_NEXTPTR_REG),
    .PF0_ARI_CAP_NEXT_FUNC (PF0_ARI_CAP_NEXT_FUNC_REG),
    .PF0_ARI_CAP_VER (PF0_ARI_CAP_VER_REG),
    .PF0_BAR0_APERTURE_SIZE (PF0_BAR0_APERTURE_SIZE_REG),
    .PF0_BAR0_CONTROL (PF0_BAR0_CONTROL_REG),
    .PF0_BAR1_APERTURE_SIZE (PF0_BAR1_APERTURE_SIZE_REG),
    .PF0_BAR1_CONTROL (PF0_BAR1_CONTROL_REG),
    .PF0_BAR2_APERTURE_SIZE (PF0_BAR2_APERTURE_SIZE_REG),
    .PF0_BAR2_CONTROL (PF0_BAR2_CONTROL_REG),
    .PF0_BAR3_APERTURE_SIZE (PF0_BAR3_APERTURE_SIZE_REG),
    .PF0_BAR3_CONTROL (PF0_BAR3_CONTROL_REG),
    .PF0_BAR4_APERTURE_SIZE (PF0_BAR4_APERTURE_SIZE_REG),
    .PF0_BAR4_CONTROL (PF0_BAR4_CONTROL_REG),
    .PF0_BAR5_APERTURE_SIZE (PF0_BAR5_APERTURE_SIZE_REG),
    .PF0_BAR5_CONTROL (PF0_BAR5_CONTROL_REG),
    .PF0_BIST_REGISTER (PF0_BIST_REGISTER_REG),
    .PF0_CAPABILITY_POINTER (PF0_CAPABILITY_POINTER_REG),
    .PF0_CLASS_CODE (PF0_CLASS_CODE_REG),
    .PF0_DEVICE_ID (PF0_DEVICE_ID_REG),
    .PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT (PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT_REG),
    .PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT (PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT_REG),
    .PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT (PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT_REG),
    .PF0_DEV_CAP2_ARI_FORWARD_ENABLE (PF0_DEV_CAP2_ARI_FORWARD_ENABLE_REG),
    .PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE (PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE_REG),
    .PF0_DEV_CAP2_LTR_SUPPORT (PF0_DEV_CAP2_LTR_SUPPORT_REG),
    .PF0_DEV_CAP2_OBFF_SUPPORT (PF0_DEV_CAP2_OBFF_SUPPORT_REG),
    .PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT (PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT_REG),
    .PF0_DEV_CAP_ENDPOINT_L0S_LATENCY (PF0_DEV_CAP_ENDPOINT_L0S_LATENCY_REG),
    .PF0_DEV_CAP_ENDPOINT_L1_LATENCY (PF0_DEV_CAP_ENDPOINT_L1_LATENCY_REG),
    .PF0_DEV_CAP_EXT_TAG_SUPPORTED (PF0_DEV_CAP_EXT_TAG_SUPPORTED_REG),
    .PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE (PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE_REG),
    .PF0_DEV_CAP_MAX_PAYLOAD_SIZE (PF0_DEV_CAP_MAX_PAYLOAD_SIZE_REG),
    .PF0_DPA_CAP_NEXTPTR (PF0_DPA_CAP_NEXTPTR_REG),
    .PF0_DPA_CAP_SUB_STATE_CONTROL (PF0_DPA_CAP_SUB_STATE_CONTROL_REG),
    .PF0_DPA_CAP_SUB_STATE_CONTROL_EN (PF0_DPA_CAP_SUB_STATE_CONTROL_EN_REG),
    .PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 (PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION0_REG),
    .PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 (PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION1_REG),
    .PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 (PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION2_REG),
    .PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 (PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION3_REG),
    .PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 (PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION4_REG),
    .PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 (PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION5_REG),
    .PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 (PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION6_REG),
    .PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 (PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION7_REG),
    .PF0_DPA_CAP_VER (PF0_DPA_CAP_VER_REG),
    .PF0_DSN_CAP_NEXTPTR (PF0_DSN_CAP_NEXTPTR_REG),
    .PF0_EXPANSION_ROM_APERTURE_SIZE (PF0_EXPANSION_ROM_APERTURE_SIZE_REG),
    .PF0_EXPANSION_ROM_ENABLE (PF0_EXPANSION_ROM_ENABLE_REG),
    .PF0_INTERRUPT_LINE (PF0_INTERRUPT_LINE_REG),
    .PF0_INTERRUPT_PIN (PF0_INTERRUPT_PIN_REG),
    .PF0_LINK_CAP_ASPM_SUPPORT (PF0_LINK_CAP_ASPM_SUPPORT_REG),
    .PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1_REG),
    .PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2_REG),
    .PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3 (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3_REG),
    .PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1 (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1_REG),
    .PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2 (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2_REG),
    .PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3 (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3_REG),
    .PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1_REG),
    .PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2_REG),
    .PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3 (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3_REG),
    .PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1 (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1_REG),
    .PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2 (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2_REG),
    .PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3 (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3_REG),
    .PF0_LINK_STATUS_SLOT_CLOCK_CONFIG (PF0_LINK_STATUS_SLOT_CLOCK_CONFIG_REG),
    .PF0_LTR_CAP_MAX_NOSNOOP_LAT (PF0_LTR_CAP_MAX_NOSNOOP_LAT_REG),
    .PF0_LTR_CAP_MAX_SNOOP_LAT (PF0_LTR_CAP_MAX_SNOOP_LAT_REG),
    .PF0_LTR_CAP_NEXTPTR (PF0_LTR_CAP_NEXTPTR_REG),
    .PF0_LTR_CAP_VER (PF0_LTR_CAP_VER_REG),
    .PF0_MSIX_CAP_NEXTPTR (PF0_MSIX_CAP_NEXTPTR_REG),
    .PF0_MSIX_CAP_PBA_BIR (PF0_MSIX_CAP_PBA_BIR_REG),
    .PF0_MSIX_CAP_PBA_OFFSET (PF0_MSIX_CAP_PBA_OFFSET_REG),
    .PF0_MSIX_CAP_TABLE_BIR (PF0_MSIX_CAP_TABLE_BIR_REG),
    .PF0_MSIX_CAP_TABLE_OFFSET (PF0_MSIX_CAP_TABLE_OFFSET_REG),
    .PF0_MSIX_CAP_TABLE_SIZE (PF0_MSIX_CAP_TABLE_SIZE_REG),
    .PF0_MSI_CAP_MULTIMSGCAP (PF0_MSI_CAP_MULTIMSGCAP_REG),
    .PF0_MSI_CAP_NEXTPTR (PF0_MSI_CAP_NEXTPTR_REG),
    .PF0_MSI_CAP_PERVECMASKCAP (PF0_MSI_CAP_PERVECMASKCAP_REG),
    .PF0_PB_CAP_DATA_REG_D0 (PF0_PB_CAP_DATA_REG_D0_REG),
    .PF0_PB_CAP_DATA_REG_D0_SUSTAINED (PF0_PB_CAP_DATA_REG_D0_SUSTAINED_REG),
    .PF0_PB_CAP_DATA_REG_D1 (PF0_PB_CAP_DATA_REG_D1_REG),
    .PF0_PB_CAP_DATA_REG_D3HOT (PF0_PB_CAP_DATA_REG_D3HOT_REG),
    .PF0_PB_CAP_NEXTPTR (PF0_PB_CAP_NEXTPTR_REG),
    .PF0_PB_CAP_SYSTEM_ALLOCATED (PF0_PB_CAP_SYSTEM_ALLOCATED_REG),
    .PF0_PB_CAP_VER (PF0_PB_CAP_VER_REG),
    .PF0_PM_CAP_ID (PF0_PM_CAP_ID_REG),
    .PF0_PM_CAP_NEXTPTR (PF0_PM_CAP_NEXTPTR_REG),
    .PF0_PM_CAP_PMESUPPORT_D0 (PF0_PM_CAP_PMESUPPORT_D0_REG),
    .PF0_PM_CAP_PMESUPPORT_D1 (PF0_PM_CAP_PMESUPPORT_D1_REG),
    .PF0_PM_CAP_PMESUPPORT_D3HOT (PF0_PM_CAP_PMESUPPORT_D3HOT_REG),
    .PF0_PM_CAP_SUPP_D1_STATE (PF0_PM_CAP_SUPP_D1_STATE_REG),
    .PF0_PM_CAP_VER_ID (PF0_PM_CAP_VER_ID_REG),
    .PF0_PM_CSR_NOSOFTRESET (PF0_PM_CSR_NOSOFTRESET_REG),
    .PF0_RBAR_CAP_ENABLE (PF0_RBAR_CAP_ENABLE_REG),
    .PF0_RBAR_CAP_NEXTPTR (PF0_RBAR_CAP_NEXTPTR_REG),
    .PF0_RBAR_CAP_SIZE0 (PF0_RBAR_CAP_SIZE0_REG),
    .PF0_RBAR_CAP_SIZE1 (PF0_RBAR_CAP_SIZE1_REG),
    .PF0_RBAR_CAP_SIZE2 (PF0_RBAR_CAP_SIZE2_REG),
    .PF0_RBAR_CAP_VER (PF0_RBAR_CAP_VER_REG),
    .PF0_RBAR_CONTROL_INDEX0 (PF0_RBAR_CONTROL_INDEX0_REG),
    .PF0_RBAR_CONTROL_INDEX1 (PF0_RBAR_CONTROL_INDEX1_REG),
    .PF0_RBAR_CONTROL_INDEX2 (PF0_RBAR_CONTROL_INDEX2_REG),
    .PF0_RBAR_CONTROL_SIZE0 (PF0_RBAR_CONTROL_SIZE0_REG),
    .PF0_RBAR_CONTROL_SIZE1 (PF0_RBAR_CONTROL_SIZE1_REG),
    .PF0_RBAR_CONTROL_SIZE2 (PF0_RBAR_CONTROL_SIZE2_REG),
    .PF0_RBAR_NUM (PF0_RBAR_NUM_REG),
    .PF0_REVISION_ID (PF0_REVISION_ID_REG),
    .PF0_SECONDARY_PCIE_CAP_NEXTPTR (PF0_SECONDARY_PCIE_CAP_NEXTPTR_REG),
    .PF0_SRIOV_BAR0_APERTURE_SIZE (PF0_SRIOV_BAR0_APERTURE_SIZE_REG),
    .PF0_SRIOV_BAR0_CONTROL (PF0_SRIOV_BAR0_CONTROL_REG),
    .PF0_SRIOV_BAR1_APERTURE_SIZE (PF0_SRIOV_BAR1_APERTURE_SIZE_REG),
    .PF0_SRIOV_BAR1_CONTROL (PF0_SRIOV_BAR1_CONTROL_REG),
    .PF0_SRIOV_BAR2_APERTURE_SIZE (PF0_SRIOV_BAR2_APERTURE_SIZE_REG),
    .PF0_SRIOV_BAR2_CONTROL (PF0_SRIOV_BAR2_CONTROL_REG),
    .PF0_SRIOV_BAR3_APERTURE_SIZE (PF0_SRIOV_BAR3_APERTURE_SIZE_REG),
    .PF0_SRIOV_BAR3_CONTROL (PF0_SRIOV_BAR3_CONTROL_REG),
    .PF0_SRIOV_BAR4_APERTURE_SIZE (PF0_SRIOV_BAR4_APERTURE_SIZE_REG),
    .PF0_SRIOV_BAR4_CONTROL (PF0_SRIOV_BAR4_CONTROL_REG),
    .PF0_SRIOV_BAR5_APERTURE_SIZE (PF0_SRIOV_BAR5_APERTURE_SIZE_REG),
    .PF0_SRIOV_BAR5_CONTROL (PF0_SRIOV_BAR5_CONTROL_REG),
    .PF0_SRIOV_CAP_INITIAL_VF (PF0_SRIOV_CAP_INITIAL_VF_REG),
    .PF0_SRIOV_CAP_NEXTPTR (PF0_SRIOV_CAP_NEXTPTR_REG),
    .PF0_SRIOV_CAP_TOTAL_VF (PF0_SRIOV_CAP_TOTAL_VF_REG),
    .PF0_SRIOV_CAP_VER (PF0_SRIOV_CAP_VER_REG),
    .PF0_SRIOV_FIRST_VF_OFFSET (PF0_SRIOV_FIRST_VF_OFFSET_REG),
    .PF0_SRIOV_FUNC_DEP_LINK (PF0_SRIOV_FUNC_DEP_LINK_REG),
    .PF0_SRIOV_SUPPORTED_PAGE_SIZE (PF0_SRIOV_SUPPORTED_PAGE_SIZE_REG),
    .PF0_SRIOV_VF_DEVICE_ID (PF0_SRIOV_VF_DEVICE_ID_REG),
    .PF0_SUBSYSTEM_ID (PF0_SUBSYSTEM_ID_REG),
    .PF0_TPHR_CAP_DEV_SPECIFIC_MODE (PF0_TPHR_CAP_DEV_SPECIFIC_MODE_REG),
    .PF0_TPHR_CAP_ENABLE (PF0_TPHR_CAP_ENABLE_REG),
    .PF0_TPHR_CAP_INT_VEC_MODE (PF0_TPHR_CAP_INT_VEC_MODE_REG),
    .PF0_TPHR_CAP_NEXTPTR (PF0_TPHR_CAP_NEXTPTR_REG),
    .PF0_TPHR_CAP_ST_MODE_SEL (PF0_TPHR_CAP_ST_MODE_SEL_REG),
    .PF0_TPHR_CAP_ST_TABLE_LOC (PF0_TPHR_CAP_ST_TABLE_LOC_REG),
    .PF0_TPHR_CAP_ST_TABLE_SIZE (PF0_TPHR_CAP_ST_TABLE_SIZE_REG),
    .PF0_TPHR_CAP_VER (PF0_TPHR_CAP_VER_REG),
    .PF0_VC_CAP_ENABLE (PF0_VC_CAP_ENABLE_REG),
    .PF0_VC_CAP_NEXTPTR (PF0_VC_CAP_NEXTPTR_REG),
    .PF0_VC_CAP_VER (PF0_VC_CAP_VER_REG),
    .PF1_AER_CAP_ECRC_CHECK_CAPABLE (PF1_AER_CAP_ECRC_CHECK_CAPABLE_REG),
    .PF1_AER_CAP_ECRC_GEN_CAPABLE (PF1_AER_CAP_ECRC_GEN_CAPABLE_REG),
    .PF1_AER_CAP_NEXTPTR (PF1_AER_CAP_NEXTPTR_REG),
    .PF1_ARI_CAP_NEXTPTR (PF1_ARI_CAP_NEXTPTR_REG),
    .PF1_ARI_CAP_NEXT_FUNC (PF1_ARI_CAP_NEXT_FUNC_REG),
    .PF1_BAR0_APERTURE_SIZE (PF1_BAR0_APERTURE_SIZE_REG),
    .PF1_BAR0_CONTROL (PF1_BAR0_CONTROL_REG),
    .PF1_BAR1_APERTURE_SIZE (PF1_BAR1_APERTURE_SIZE_REG),
    .PF1_BAR1_CONTROL (PF1_BAR1_CONTROL_REG),
    .PF1_BAR2_APERTURE_SIZE (PF1_BAR2_APERTURE_SIZE_REG),
    .PF1_BAR2_CONTROL (PF1_BAR2_CONTROL_REG),
    .PF1_BAR3_APERTURE_SIZE (PF1_BAR3_APERTURE_SIZE_REG),
    .PF1_BAR3_CONTROL (PF1_BAR3_CONTROL_REG),
    .PF1_BAR4_APERTURE_SIZE (PF1_BAR4_APERTURE_SIZE_REG),
    .PF1_BAR4_CONTROL (PF1_BAR4_CONTROL_REG),
    .PF1_BAR5_APERTURE_SIZE (PF1_BAR5_APERTURE_SIZE_REG),
    .PF1_BAR5_CONTROL (PF1_BAR5_CONTROL_REG),
    .PF1_BIST_REGISTER (PF1_BIST_REGISTER_REG),
    .PF1_CAPABILITY_POINTER (PF1_CAPABILITY_POINTER_REG),
    .PF1_CLASS_CODE (PF1_CLASS_CODE_REG),
    .PF1_DEVICE_ID (PF1_DEVICE_ID_REG),
    .PF1_DEV_CAP_MAX_PAYLOAD_SIZE (PF1_DEV_CAP_MAX_PAYLOAD_SIZE_REG),
    .PF1_DPA_CAP_NEXTPTR (PF1_DPA_CAP_NEXTPTR_REG),
    .PF1_DPA_CAP_SUB_STATE_CONTROL (PF1_DPA_CAP_SUB_STATE_CONTROL_REG),
    .PF1_DPA_CAP_SUB_STATE_CONTROL_EN (PF1_DPA_CAP_SUB_STATE_CONTROL_EN_REG),
    .PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 (PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION0_REG),
    .PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 (PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION1_REG),
    .PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 (PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION2_REG),
    .PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 (PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION3_REG),
    .PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 (PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION4_REG),
    .PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 (PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION5_REG),
    .PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 (PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION6_REG),
    .PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 (PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION7_REG),
    .PF1_DPA_CAP_VER (PF1_DPA_CAP_VER_REG),
    .PF1_DSN_CAP_NEXTPTR (PF1_DSN_CAP_NEXTPTR_REG),
    .PF1_EXPANSION_ROM_APERTURE_SIZE (PF1_EXPANSION_ROM_APERTURE_SIZE_REG),
    .PF1_EXPANSION_ROM_ENABLE (PF1_EXPANSION_ROM_ENABLE_REG),
    .PF1_INTERRUPT_LINE (PF1_INTERRUPT_LINE_REG),
    .PF1_INTERRUPT_PIN (PF1_INTERRUPT_PIN_REG),
    .PF1_MSIX_CAP_NEXTPTR (PF1_MSIX_CAP_NEXTPTR_REG),
    .PF1_MSIX_CAP_PBA_BIR (PF1_MSIX_CAP_PBA_BIR_REG),
    .PF1_MSIX_CAP_PBA_OFFSET (PF1_MSIX_CAP_PBA_OFFSET_REG),
    .PF1_MSIX_CAP_TABLE_BIR (PF1_MSIX_CAP_TABLE_BIR_REG),
    .PF1_MSIX_CAP_TABLE_OFFSET (PF1_MSIX_CAP_TABLE_OFFSET_REG),
    .PF1_MSIX_CAP_TABLE_SIZE (PF1_MSIX_CAP_TABLE_SIZE_REG),
    .PF1_MSI_CAP_MULTIMSGCAP (PF1_MSI_CAP_MULTIMSGCAP_REG),
    .PF1_MSI_CAP_NEXTPTR (PF1_MSI_CAP_NEXTPTR_REG),
    .PF1_MSI_CAP_PERVECMASKCAP (PF1_MSI_CAP_PERVECMASKCAP_REG),
    .PF1_PB_CAP_DATA_REG_D0 (PF1_PB_CAP_DATA_REG_D0_REG),
    .PF1_PB_CAP_DATA_REG_D0_SUSTAINED (PF1_PB_CAP_DATA_REG_D0_SUSTAINED_REG),
    .PF1_PB_CAP_DATA_REG_D1 (PF1_PB_CAP_DATA_REG_D1_REG),
    .PF1_PB_CAP_DATA_REG_D3HOT (PF1_PB_CAP_DATA_REG_D3HOT_REG),
    .PF1_PB_CAP_NEXTPTR (PF1_PB_CAP_NEXTPTR_REG),
    .PF1_PB_CAP_SYSTEM_ALLOCATED (PF1_PB_CAP_SYSTEM_ALLOCATED_REG),
    .PF1_PB_CAP_VER (PF1_PB_CAP_VER_REG),
    .PF1_PM_CAP_ID (PF1_PM_CAP_ID_REG),
    .PF1_PM_CAP_NEXTPTR (PF1_PM_CAP_NEXTPTR_REG),
    .PF1_PM_CAP_VER_ID (PF1_PM_CAP_VER_ID_REG),
    .PF1_RBAR_CAP_ENABLE (PF1_RBAR_CAP_ENABLE_REG),
    .PF1_RBAR_CAP_NEXTPTR (PF1_RBAR_CAP_NEXTPTR_REG),
    .PF1_RBAR_CAP_SIZE0 (PF1_RBAR_CAP_SIZE0_REG),
    .PF1_RBAR_CAP_SIZE1 (PF1_RBAR_CAP_SIZE1_REG),
    .PF1_RBAR_CAP_SIZE2 (PF1_RBAR_CAP_SIZE2_REG),
    .PF1_RBAR_CAP_VER (PF1_RBAR_CAP_VER_REG),
    .PF1_RBAR_CONTROL_INDEX0 (PF1_RBAR_CONTROL_INDEX0_REG),
    .PF1_RBAR_CONTROL_INDEX1 (PF1_RBAR_CONTROL_INDEX1_REG),
    .PF1_RBAR_CONTROL_INDEX2 (PF1_RBAR_CONTROL_INDEX2_REG),
    .PF1_RBAR_CONTROL_SIZE0 (PF1_RBAR_CONTROL_SIZE0_REG),
    .PF1_RBAR_CONTROL_SIZE1 (PF1_RBAR_CONTROL_SIZE1_REG),
    .PF1_RBAR_CONTROL_SIZE2 (PF1_RBAR_CONTROL_SIZE2_REG),
    .PF1_RBAR_NUM (PF1_RBAR_NUM_REG),
    .PF1_REVISION_ID (PF1_REVISION_ID_REG),
    .PF1_SRIOV_BAR0_APERTURE_SIZE (PF1_SRIOV_BAR0_APERTURE_SIZE_REG),
    .PF1_SRIOV_BAR0_CONTROL (PF1_SRIOV_BAR0_CONTROL_REG),
    .PF1_SRIOV_BAR1_APERTURE_SIZE (PF1_SRIOV_BAR1_APERTURE_SIZE_REG),
    .PF1_SRIOV_BAR1_CONTROL (PF1_SRIOV_BAR1_CONTROL_REG),
    .PF1_SRIOV_BAR2_APERTURE_SIZE (PF1_SRIOV_BAR2_APERTURE_SIZE_REG),
    .PF1_SRIOV_BAR2_CONTROL (PF1_SRIOV_BAR2_CONTROL_REG),
    .PF1_SRIOV_BAR3_APERTURE_SIZE (PF1_SRIOV_BAR3_APERTURE_SIZE_REG),
    .PF1_SRIOV_BAR3_CONTROL (PF1_SRIOV_BAR3_CONTROL_REG),
    .PF1_SRIOV_BAR4_APERTURE_SIZE (PF1_SRIOV_BAR4_APERTURE_SIZE_REG),
    .PF1_SRIOV_BAR4_CONTROL (PF1_SRIOV_BAR4_CONTROL_REG),
    .PF1_SRIOV_BAR5_APERTURE_SIZE (PF1_SRIOV_BAR5_APERTURE_SIZE_REG),
    .PF1_SRIOV_BAR5_CONTROL (PF1_SRIOV_BAR5_CONTROL_REG),
    .PF1_SRIOV_CAP_INITIAL_VF (PF1_SRIOV_CAP_INITIAL_VF_REG),
    .PF1_SRIOV_CAP_NEXTPTR (PF1_SRIOV_CAP_NEXTPTR_REG),
    .PF1_SRIOV_CAP_TOTAL_VF (PF1_SRIOV_CAP_TOTAL_VF_REG),
    .PF1_SRIOV_CAP_VER (PF1_SRIOV_CAP_VER_REG),
    .PF1_SRIOV_FIRST_VF_OFFSET (PF1_SRIOV_FIRST_VF_OFFSET_REG),
    .PF1_SRIOV_FUNC_DEP_LINK (PF1_SRIOV_FUNC_DEP_LINK_REG),
    .PF1_SRIOV_SUPPORTED_PAGE_SIZE (PF1_SRIOV_SUPPORTED_PAGE_SIZE_REG),
    .PF1_SRIOV_VF_DEVICE_ID (PF1_SRIOV_VF_DEVICE_ID_REG),
    .PF1_SUBSYSTEM_ID (PF1_SUBSYSTEM_ID_REG),
    .PF1_TPHR_CAP_DEV_SPECIFIC_MODE (PF1_TPHR_CAP_DEV_SPECIFIC_MODE_REG),
    .PF1_TPHR_CAP_ENABLE (PF1_TPHR_CAP_ENABLE_REG),
    .PF1_TPHR_CAP_INT_VEC_MODE (PF1_TPHR_CAP_INT_VEC_MODE_REG),
    .PF1_TPHR_CAP_NEXTPTR (PF1_TPHR_CAP_NEXTPTR_REG),
    .PF1_TPHR_CAP_ST_MODE_SEL (PF1_TPHR_CAP_ST_MODE_SEL_REG),
    .PF1_TPHR_CAP_ST_TABLE_LOC (PF1_TPHR_CAP_ST_TABLE_LOC_REG),
    .PF1_TPHR_CAP_ST_TABLE_SIZE (PF1_TPHR_CAP_ST_TABLE_SIZE_REG),
    .PF1_TPHR_CAP_VER (PF1_TPHR_CAP_VER_REG),
    .PF2_AER_CAP_ECRC_CHECK_CAPABLE (PF2_AER_CAP_ECRC_CHECK_CAPABLE_REG),
    .PF2_AER_CAP_ECRC_GEN_CAPABLE (PF2_AER_CAP_ECRC_GEN_CAPABLE_REG),
    .PF2_AER_CAP_NEXTPTR (PF2_AER_CAP_NEXTPTR_REG),
    .PF2_ARI_CAP_NEXTPTR (PF2_ARI_CAP_NEXTPTR_REG),
    .PF2_ARI_CAP_NEXT_FUNC (PF2_ARI_CAP_NEXT_FUNC_REG),
    .PF2_BAR0_APERTURE_SIZE (PF2_BAR0_APERTURE_SIZE_REG),
    .PF2_BAR0_CONTROL (PF2_BAR0_CONTROL_REG),
    .PF2_BAR1_APERTURE_SIZE (PF2_BAR1_APERTURE_SIZE_REG),
    .PF2_BAR1_CONTROL (PF2_BAR1_CONTROL_REG),
    .PF2_BAR2_APERTURE_SIZE (PF2_BAR2_APERTURE_SIZE_REG),
    .PF2_BAR2_CONTROL (PF2_BAR2_CONTROL_REG),
    .PF2_BAR3_APERTURE_SIZE (PF2_BAR3_APERTURE_SIZE_REG),
    .PF2_BAR3_CONTROL (PF2_BAR3_CONTROL_REG),
    .PF2_BAR4_APERTURE_SIZE (PF2_BAR4_APERTURE_SIZE_REG),
    .PF2_BAR4_CONTROL (PF2_BAR4_CONTROL_REG),
    .PF2_BAR5_APERTURE_SIZE (PF2_BAR5_APERTURE_SIZE_REG),
    .PF2_BAR5_CONTROL (PF2_BAR5_CONTROL_REG),
    .PF2_BIST_REGISTER (PF2_BIST_REGISTER_REG),
    .PF2_CAPABILITY_POINTER (PF2_CAPABILITY_POINTER_REG),
    .PF2_CLASS_CODE (PF2_CLASS_CODE_REG),
    .PF2_DEVICE_ID (PF2_DEVICE_ID_REG),
    .PF2_DEV_CAP_MAX_PAYLOAD_SIZE (PF2_DEV_CAP_MAX_PAYLOAD_SIZE_REG),
    .PF2_DPA_CAP_NEXTPTR (PF2_DPA_CAP_NEXTPTR_REG),
    .PF2_DPA_CAP_SUB_STATE_CONTROL (PF2_DPA_CAP_SUB_STATE_CONTROL_REG),
    .PF2_DPA_CAP_SUB_STATE_CONTROL_EN (PF2_DPA_CAP_SUB_STATE_CONTROL_EN_REG),
    .PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 (PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION0_REG),
    .PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 (PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION1_REG),
    .PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 (PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION2_REG),
    .PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 (PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION3_REG),
    .PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 (PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION4_REG),
    .PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 (PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION5_REG),
    .PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 (PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION6_REG),
    .PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 (PF2_DPA_CAP_SUB_STATE_POWER_ALLOCATION7_REG),
    .PF2_DPA_CAP_VER (PF2_DPA_CAP_VER_REG),
    .PF2_DSN_CAP_NEXTPTR (PF2_DSN_CAP_NEXTPTR_REG),
    .PF2_EXPANSION_ROM_APERTURE_SIZE (PF2_EXPANSION_ROM_APERTURE_SIZE_REG),
    .PF2_EXPANSION_ROM_ENABLE (PF2_EXPANSION_ROM_ENABLE_REG),
    .PF2_INTERRUPT_LINE (PF2_INTERRUPT_LINE_REG),
    .PF2_INTERRUPT_PIN (PF2_INTERRUPT_PIN_REG),
    .PF2_MSIX_CAP_NEXTPTR (PF2_MSIX_CAP_NEXTPTR_REG),
    .PF2_MSIX_CAP_PBA_BIR (PF2_MSIX_CAP_PBA_BIR_REG),
    .PF2_MSIX_CAP_PBA_OFFSET (PF2_MSIX_CAP_PBA_OFFSET_REG),
    .PF2_MSIX_CAP_TABLE_BIR (PF2_MSIX_CAP_TABLE_BIR_REG),
    .PF2_MSIX_CAP_TABLE_OFFSET (PF2_MSIX_CAP_TABLE_OFFSET_REG),
    .PF2_MSIX_CAP_TABLE_SIZE (PF2_MSIX_CAP_TABLE_SIZE_REG),
    .PF2_MSI_CAP_MULTIMSGCAP (PF2_MSI_CAP_MULTIMSGCAP_REG),
    .PF2_MSI_CAP_NEXTPTR (PF2_MSI_CAP_NEXTPTR_REG),
    .PF2_MSI_CAP_PERVECMASKCAP (PF2_MSI_CAP_PERVECMASKCAP_REG),
    .PF2_PB_CAP_DATA_REG_D0 (PF2_PB_CAP_DATA_REG_D0_REG),
    .PF2_PB_CAP_DATA_REG_D0_SUSTAINED (PF2_PB_CAP_DATA_REG_D0_SUSTAINED_REG),
    .PF2_PB_CAP_DATA_REG_D1 (PF2_PB_CAP_DATA_REG_D1_REG),
    .PF2_PB_CAP_DATA_REG_D3HOT (PF2_PB_CAP_DATA_REG_D3HOT_REG),
    .PF2_PB_CAP_NEXTPTR (PF2_PB_CAP_NEXTPTR_REG),
    .PF2_PB_CAP_SYSTEM_ALLOCATED (PF2_PB_CAP_SYSTEM_ALLOCATED_REG),
    .PF2_PB_CAP_VER (PF2_PB_CAP_VER_REG),
    .PF2_PM_CAP_ID (PF2_PM_CAP_ID_REG),
    .PF2_PM_CAP_NEXTPTR (PF2_PM_CAP_NEXTPTR_REG),
    .PF2_PM_CAP_VER_ID (PF2_PM_CAP_VER_ID_REG),
    .PF2_RBAR_CAP_ENABLE (PF2_RBAR_CAP_ENABLE_REG),
    .PF2_RBAR_CAP_NEXTPTR (PF2_RBAR_CAP_NEXTPTR_REG),
    .PF2_RBAR_CAP_SIZE0 (PF2_RBAR_CAP_SIZE0_REG),
    .PF2_RBAR_CAP_SIZE1 (PF2_RBAR_CAP_SIZE1_REG),
    .PF2_RBAR_CAP_SIZE2 (PF2_RBAR_CAP_SIZE2_REG),
    .PF2_RBAR_CAP_VER (PF2_RBAR_CAP_VER_REG),
    .PF2_RBAR_CONTROL_INDEX0 (PF2_RBAR_CONTROL_INDEX0_REG),
    .PF2_RBAR_CONTROL_INDEX1 (PF2_RBAR_CONTROL_INDEX1_REG),
    .PF2_RBAR_CONTROL_INDEX2 (PF2_RBAR_CONTROL_INDEX2_REG),
    .PF2_RBAR_CONTROL_SIZE0 (PF2_RBAR_CONTROL_SIZE0_REG),
    .PF2_RBAR_CONTROL_SIZE1 (PF2_RBAR_CONTROL_SIZE1_REG),
    .PF2_RBAR_CONTROL_SIZE2 (PF2_RBAR_CONTROL_SIZE2_REG),
    .PF2_RBAR_NUM (PF2_RBAR_NUM_REG),
    .PF2_REVISION_ID (PF2_REVISION_ID_REG),
    .PF2_SRIOV_BAR0_APERTURE_SIZE (PF2_SRIOV_BAR0_APERTURE_SIZE_REG),
    .PF2_SRIOV_BAR0_CONTROL (PF2_SRIOV_BAR0_CONTROL_REG),
    .PF2_SRIOV_BAR1_APERTURE_SIZE (PF2_SRIOV_BAR1_APERTURE_SIZE_REG),
    .PF2_SRIOV_BAR1_CONTROL (PF2_SRIOV_BAR1_CONTROL_REG),
    .PF2_SRIOV_BAR2_APERTURE_SIZE (PF2_SRIOV_BAR2_APERTURE_SIZE_REG),
    .PF2_SRIOV_BAR2_CONTROL (PF2_SRIOV_BAR2_CONTROL_REG),
    .PF2_SRIOV_BAR3_APERTURE_SIZE (PF2_SRIOV_BAR3_APERTURE_SIZE_REG),
    .PF2_SRIOV_BAR3_CONTROL (PF2_SRIOV_BAR3_CONTROL_REG),
    .PF2_SRIOV_BAR4_APERTURE_SIZE (PF2_SRIOV_BAR4_APERTURE_SIZE_REG),
    .PF2_SRIOV_BAR4_CONTROL (PF2_SRIOV_BAR4_CONTROL_REG),
    .PF2_SRIOV_BAR5_APERTURE_SIZE (PF2_SRIOV_BAR5_APERTURE_SIZE_REG),
    .PF2_SRIOV_BAR5_CONTROL (PF2_SRIOV_BAR5_CONTROL_REG),
    .PF2_SRIOV_CAP_INITIAL_VF (PF2_SRIOV_CAP_INITIAL_VF_REG),
    .PF2_SRIOV_CAP_NEXTPTR (PF2_SRIOV_CAP_NEXTPTR_REG),
    .PF2_SRIOV_CAP_TOTAL_VF (PF2_SRIOV_CAP_TOTAL_VF_REG),
    .PF2_SRIOV_CAP_VER (PF2_SRIOV_CAP_VER_REG),
    .PF2_SRIOV_FIRST_VF_OFFSET (PF2_SRIOV_FIRST_VF_OFFSET_REG),
    .PF2_SRIOV_FUNC_DEP_LINK (PF2_SRIOV_FUNC_DEP_LINK_REG),
    .PF2_SRIOV_SUPPORTED_PAGE_SIZE (PF2_SRIOV_SUPPORTED_PAGE_SIZE_REG),
    .PF2_SRIOV_VF_DEVICE_ID (PF2_SRIOV_VF_DEVICE_ID_REG),
    .PF2_SUBSYSTEM_ID (PF2_SUBSYSTEM_ID_REG),
    .PF2_TPHR_CAP_DEV_SPECIFIC_MODE (PF2_TPHR_CAP_DEV_SPECIFIC_MODE_REG),
    .PF2_TPHR_CAP_ENABLE (PF2_TPHR_CAP_ENABLE_REG),
    .PF2_TPHR_CAP_INT_VEC_MODE (PF2_TPHR_CAP_INT_VEC_MODE_REG),
    .PF2_TPHR_CAP_NEXTPTR (PF2_TPHR_CAP_NEXTPTR_REG),
    .PF2_TPHR_CAP_ST_MODE_SEL (PF2_TPHR_CAP_ST_MODE_SEL_REG),
    .PF2_TPHR_CAP_ST_TABLE_LOC (PF2_TPHR_CAP_ST_TABLE_LOC_REG),
    .PF2_TPHR_CAP_ST_TABLE_SIZE (PF2_TPHR_CAP_ST_TABLE_SIZE_REG),
    .PF2_TPHR_CAP_VER (PF2_TPHR_CAP_VER_REG),
    .PF3_AER_CAP_ECRC_CHECK_CAPABLE (PF3_AER_CAP_ECRC_CHECK_CAPABLE_REG),
    .PF3_AER_CAP_ECRC_GEN_CAPABLE (PF3_AER_CAP_ECRC_GEN_CAPABLE_REG),
    .PF3_AER_CAP_NEXTPTR (PF3_AER_CAP_NEXTPTR_REG),
    .PF3_ARI_CAP_NEXTPTR (PF3_ARI_CAP_NEXTPTR_REG),
    .PF3_ARI_CAP_NEXT_FUNC (PF3_ARI_CAP_NEXT_FUNC_REG),
    .PF3_BAR0_APERTURE_SIZE (PF3_BAR0_APERTURE_SIZE_REG),
    .PF3_BAR0_CONTROL (PF3_BAR0_CONTROL_REG),
    .PF3_BAR1_APERTURE_SIZE (PF3_BAR1_APERTURE_SIZE_REG),
    .PF3_BAR1_CONTROL (PF3_BAR1_CONTROL_REG),
    .PF3_BAR2_APERTURE_SIZE (PF3_BAR2_APERTURE_SIZE_REG),
    .PF3_BAR2_CONTROL (PF3_BAR2_CONTROL_REG),
    .PF3_BAR3_APERTURE_SIZE (PF3_BAR3_APERTURE_SIZE_REG),
    .PF3_BAR3_CONTROL (PF3_BAR3_CONTROL_REG),
    .PF3_BAR4_APERTURE_SIZE (PF3_BAR4_APERTURE_SIZE_REG),
    .PF3_BAR4_CONTROL (PF3_BAR4_CONTROL_REG),
    .PF3_BAR5_APERTURE_SIZE (PF3_BAR5_APERTURE_SIZE_REG),
    .PF3_BAR5_CONTROL (PF3_BAR5_CONTROL_REG),
    .PF3_BIST_REGISTER (PF3_BIST_REGISTER_REG),
    .PF3_CAPABILITY_POINTER (PF3_CAPABILITY_POINTER_REG),
    .PF3_CLASS_CODE (PF3_CLASS_CODE_REG),
    .PF3_DEVICE_ID (PF3_DEVICE_ID_REG),
    .PF3_DEV_CAP_MAX_PAYLOAD_SIZE (PF3_DEV_CAP_MAX_PAYLOAD_SIZE_REG),
    .PF3_DPA_CAP_NEXTPTR (PF3_DPA_CAP_NEXTPTR_REG),
    .PF3_DPA_CAP_SUB_STATE_CONTROL (PF3_DPA_CAP_SUB_STATE_CONTROL_REG),
    .PF3_DPA_CAP_SUB_STATE_CONTROL_EN (PF3_DPA_CAP_SUB_STATE_CONTROL_EN_REG),
    .PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 (PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION0_REG),
    .PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 (PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION1_REG),
    .PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 (PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION2_REG),
    .PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 (PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION3_REG),
    .PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 (PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION4_REG),
    .PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 (PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION5_REG),
    .PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 (PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION6_REG),
    .PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 (PF3_DPA_CAP_SUB_STATE_POWER_ALLOCATION7_REG),
    .PF3_DPA_CAP_VER (PF3_DPA_CAP_VER_REG),
    .PF3_DSN_CAP_NEXTPTR (PF3_DSN_CAP_NEXTPTR_REG),
    .PF3_EXPANSION_ROM_APERTURE_SIZE (PF3_EXPANSION_ROM_APERTURE_SIZE_REG),
    .PF3_EXPANSION_ROM_ENABLE (PF3_EXPANSION_ROM_ENABLE_REG),
    .PF3_INTERRUPT_LINE (PF3_INTERRUPT_LINE_REG),
    .PF3_INTERRUPT_PIN (PF3_INTERRUPT_PIN_REG),
    .PF3_MSIX_CAP_NEXTPTR (PF3_MSIX_CAP_NEXTPTR_REG),
    .PF3_MSIX_CAP_PBA_BIR (PF3_MSIX_CAP_PBA_BIR_REG),
    .PF3_MSIX_CAP_PBA_OFFSET (PF3_MSIX_CAP_PBA_OFFSET_REG),
    .PF3_MSIX_CAP_TABLE_BIR (PF3_MSIX_CAP_TABLE_BIR_REG),
    .PF3_MSIX_CAP_TABLE_OFFSET (PF3_MSIX_CAP_TABLE_OFFSET_REG),
    .PF3_MSIX_CAP_TABLE_SIZE (PF3_MSIX_CAP_TABLE_SIZE_REG),
    .PF3_MSI_CAP_MULTIMSGCAP (PF3_MSI_CAP_MULTIMSGCAP_REG),
    .PF3_MSI_CAP_NEXTPTR (PF3_MSI_CAP_NEXTPTR_REG),
    .PF3_MSI_CAP_PERVECMASKCAP (PF3_MSI_CAP_PERVECMASKCAP_REG),
    .PF3_PB_CAP_DATA_REG_D0 (PF3_PB_CAP_DATA_REG_D0_REG),
    .PF3_PB_CAP_DATA_REG_D0_SUSTAINED (PF3_PB_CAP_DATA_REG_D0_SUSTAINED_REG),
    .PF3_PB_CAP_DATA_REG_D1 (PF3_PB_CAP_DATA_REG_D1_REG),
    .PF3_PB_CAP_DATA_REG_D3HOT (PF3_PB_CAP_DATA_REG_D3HOT_REG),
    .PF3_PB_CAP_NEXTPTR (PF3_PB_CAP_NEXTPTR_REG),
    .PF3_PB_CAP_SYSTEM_ALLOCATED (PF3_PB_CAP_SYSTEM_ALLOCATED_REG),
    .PF3_PB_CAP_VER (PF3_PB_CAP_VER_REG),
    .PF3_PM_CAP_ID (PF3_PM_CAP_ID_REG),
    .PF3_PM_CAP_NEXTPTR (PF3_PM_CAP_NEXTPTR_REG),
    .PF3_PM_CAP_VER_ID (PF3_PM_CAP_VER_ID_REG),
    .PF3_RBAR_CAP_ENABLE (PF3_RBAR_CAP_ENABLE_REG),
    .PF3_RBAR_CAP_NEXTPTR (PF3_RBAR_CAP_NEXTPTR_REG),
    .PF3_RBAR_CAP_SIZE0 (PF3_RBAR_CAP_SIZE0_REG),
    .PF3_RBAR_CAP_SIZE1 (PF3_RBAR_CAP_SIZE1_REG),
    .PF3_RBAR_CAP_SIZE2 (PF3_RBAR_CAP_SIZE2_REG),
    .PF3_RBAR_CAP_VER (PF3_RBAR_CAP_VER_REG),
    .PF3_RBAR_CONTROL_INDEX0 (PF3_RBAR_CONTROL_INDEX0_REG),
    .PF3_RBAR_CONTROL_INDEX1 (PF3_RBAR_CONTROL_INDEX1_REG),
    .PF3_RBAR_CONTROL_INDEX2 (PF3_RBAR_CONTROL_INDEX2_REG),
    .PF3_RBAR_CONTROL_SIZE0 (PF3_RBAR_CONTROL_SIZE0_REG),
    .PF3_RBAR_CONTROL_SIZE1 (PF3_RBAR_CONTROL_SIZE1_REG),
    .PF3_RBAR_CONTROL_SIZE2 (PF3_RBAR_CONTROL_SIZE2_REG),
    .PF3_RBAR_NUM (PF3_RBAR_NUM_REG),
    .PF3_REVISION_ID (PF3_REVISION_ID_REG),
    .PF3_SRIOV_BAR0_APERTURE_SIZE (PF3_SRIOV_BAR0_APERTURE_SIZE_REG),
    .PF3_SRIOV_BAR0_CONTROL (PF3_SRIOV_BAR0_CONTROL_REG),
    .PF3_SRIOV_BAR1_APERTURE_SIZE (PF3_SRIOV_BAR1_APERTURE_SIZE_REG),
    .PF3_SRIOV_BAR1_CONTROL (PF3_SRIOV_BAR1_CONTROL_REG),
    .PF3_SRIOV_BAR2_APERTURE_SIZE (PF3_SRIOV_BAR2_APERTURE_SIZE_REG),
    .PF3_SRIOV_BAR2_CONTROL (PF3_SRIOV_BAR2_CONTROL_REG),
    .PF3_SRIOV_BAR3_APERTURE_SIZE (PF3_SRIOV_BAR3_APERTURE_SIZE_REG),
    .PF3_SRIOV_BAR3_CONTROL (PF3_SRIOV_BAR3_CONTROL_REG),
    .PF3_SRIOV_BAR4_APERTURE_SIZE (PF3_SRIOV_BAR4_APERTURE_SIZE_REG),
    .PF3_SRIOV_BAR4_CONTROL (PF3_SRIOV_BAR4_CONTROL_REG),
    .PF3_SRIOV_BAR5_APERTURE_SIZE (PF3_SRIOV_BAR5_APERTURE_SIZE_REG),
    .PF3_SRIOV_BAR5_CONTROL (PF3_SRIOV_BAR5_CONTROL_REG),
    .PF3_SRIOV_CAP_INITIAL_VF (PF3_SRIOV_CAP_INITIAL_VF_REG),
    .PF3_SRIOV_CAP_NEXTPTR (PF3_SRIOV_CAP_NEXTPTR_REG),
    .PF3_SRIOV_CAP_TOTAL_VF (PF3_SRIOV_CAP_TOTAL_VF_REG),
    .PF3_SRIOV_CAP_VER (PF3_SRIOV_CAP_VER_REG),
    .PF3_SRIOV_FIRST_VF_OFFSET (PF3_SRIOV_FIRST_VF_OFFSET_REG),
    .PF3_SRIOV_FUNC_DEP_LINK (PF3_SRIOV_FUNC_DEP_LINK_REG),
    .PF3_SRIOV_SUPPORTED_PAGE_SIZE (PF3_SRIOV_SUPPORTED_PAGE_SIZE_REG),
    .PF3_SRIOV_VF_DEVICE_ID (PF3_SRIOV_VF_DEVICE_ID_REG),
    .PF3_SUBSYSTEM_ID (PF3_SUBSYSTEM_ID_REG),
    .PF3_TPHR_CAP_DEV_SPECIFIC_MODE (PF3_TPHR_CAP_DEV_SPECIFIC_MODE_REG),
    .PF3_TPHR_CAP_ENABLE (PF3_TPHR_CAP_ENABLE_REG),
    .PF3_TPHR_CAP_INT_VEC_MODE (PF3_TPHR_CAP_INT_VEC_MODE_REG),
    .PF3_TPHR_CAP_NEXTPTR (PF3_TPHR_CAP_NEXTPTR_REG),
    .PF3_TPHR_CAP_ST_MODE_SEL (PF3_TPHR_CAP_ST_MODE_SEL_REG),
    .PF3_TPHR_CAP_ST_TABLE_LOC (PF3_TPHR_CAP_ST_TABLE_LOC_REG),
    .PF3_TPHR_CAP_ST_TABLE_SIZE (PF3_TPHR_CAP_ST_TABLE_SIZE_REG),
    .PF3_TPHR_CAP_VER (PF3_TPHR_CAP_VER_REG),
    .PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3 (PL_DISABLE_AUTO_EQ_SPEED_CHANGE_TO_GEN3_REG),
    .PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2 (PL_DISABLE_AUTO_SPEED_CHANGE_TO_GEN2_REG),
    .PL_DISABLE_EI_INFER_IN_L0 (PL_DISABLE_EI_INFER_IN_L0_REG),
    .PL_DISABLE_GEN3_DC_BALANCE (PL_DISABLE_GEN3_DC_BALANCE_REG),
    .PL_DISABLE_GEN3_LFSR_UPDATE_ON_SKP (PL_DISABLE_GEN3_LFSR_UPDATE_ON_SKP_REG),
    .PL_DISABLE_RETRAIN_ON_FRAMING_ERROR (PL_DISABLE_RETRAIN_ON_FRAMING_ERROR_REG),
    .PL_DISABLE_SCRAMBLING (PL_DISABLE_SCRAMBLING_REG),
    .PL_DISABLE_SYNC_HEADER_FRAMING_ERROR (PL_DISABLE_SYNC_HEADER_FRAMING_ERROR_REG),
    .PL_DISABLE_UPCONFIG_CAPABLE (PL_DISABLE_UPCONFIG_CAPABLE_REG),
    .PL_EQ_ADAPT_DISABLE_COEFF_CHECK (PL_EQ_ADAPT_DISABLE_COEFF_CHECK_REG),
    .PL_EQ_ADAPT_DISABLE_PRESET_CHECK (PL_EQ_ADAPT_DISABLE_PRESET_CHECK_REG),
    .PL_EQ_ADAPT_ITER_COUNT (PL_EQ_ADAPT_ITER_COUNT_REG),
    .PL_EQ_ADAPT_REJECT_RETRY_COUNT (PL_EQ_ADAPT_REJECT_RETRY_COUNT_REG),
    .PL_EQ_BYPASS_PHASE23 (PL_EQ_BYPASS_PHASE23_REG),
    .PL_EQ_DEFAULT_GEN3_RX_PRESET_HINT (PL_EQ_DEFAULT_GEN3_RX_PRESET_HINT_REG),
    .PL_EQ_DEFAULT_GEN3_TX_PRESET (PL_EQ_DEFAULT_GEN3_TX_PRESET_REG),
    .PL_EQ_PHASE01_RX_ADAPT (PL_EQ_PHASE01_RX_ADAPT_REG),
    .PL_EQ_SHORT_ADAPT_PHASE (PL_EQ_SHORT_ADAPT_PHASE_REG),
    .PL_LANE0_EQ_CONTROL (PL_LANE0_EQ_CONTROL_REG),
    .PL_LANE1_EQ_CONTROL (PL_LANE1_EQ_CONTROL_REG),
    .PL_LANE2_EQ_CONTROL (PL_LANE2_EQ_CONTROL_REG),
    .PL_LANE3_EQ_CONTROL (PL_LANE3_EQ_CONTROL_REG),
    .PL_LANE4_EQ_CONTROL (PL_LANE4_EQ_CONTROL_REG),
    .PL_LANE5_EQ_CONTROL (PL_LANE5_EQ_CONTROL_REG),
    .PL_LANE6_EQ_CONTROL (PL_LANE6_EQ_CONTROL_REG),
    .PL_LANE7_EQ_CONTROL (PL_LANE7_EQ_CONTROL_REG),
    .PL_LINK_CAP_MAX_LINK_SPEED (PL_LINK_CAP_MAX_LINK_SPEED_REG),
    .PL_LINK_CAP_MAX_LINK_WIDTH (PL_LINK_CAP_MAX_LINK_WIDTH_REG),
    .PL_N_FTS_COMCLK_GEN1 (PL_N_FTS_COMCLK_GEN1_REG),
    .PL_N_FTS_COMCLK_GEN2 (PL_N_FTS_COMCLK_GEN2_REG),
    .PL_N_FTS_COMCLK_GEN3 (PL_N_FTS_COMCLK_GEN3_REG),
    .PL_N_FTS_GEN1 (PL_N_FTS_GEN1_REG),
    .PL_N_FTS_GEN2 (PL_N_FTS_GEN2_REG),
    .PL_N_FTS_GEN3 (PL_N_FTS_GEN3_REG),
    .PL_REPORT_ALL_PHY_ERRORS (PL_REPORT_ALL_PHY_ERRORS_REG),
    .PL_SIM_FAST_LINK_TRAINING (PL_SIM_FAST_LINK_TRAINING_REG),
    .PL_UPSTREAM_FACING (PL_UPSTREAM_FACING_REG),
    .PM_ASPML0S_TIMEOUT (PM_ASPML0S_TIMEOUT_REG),
    .PM_ASPML1_ENTRY_DELAY (PM_ASPML1_ENTRY_DELAY_REG),
    .PM_ENABLE_L23_ENTRY (PM_ENABLE_L23_ENTRY_REG),
    .PM_ENABLE_SLOT_POWER_CAPTURE (PM_ENABLE_SLOT_POWER_CAPTURE_REG),
    .PM_L1_REENTRY_DELAY (PM_L1_REENTRY_DELAY_REG),
    .PM_PME_SERVICE_TIMEOUT_DELAY (PM_PME_SERVICE_TIMEOUT_DELAY_REG),
    .PM_PME_TURNOFF_ACK_DELAY (PM_PME_TURNOFF_ACK_DELAY_REG),
    .SPARE_BIT0 (SPARE_BIT0_REG),
    .SPARE_BIT1 (SPARE_BIT1_REG),
    .SPARE_BIT2 (SPARE_BIT2_REG),
    .SPARE_BIT3 (SPARE_BIT3_REG),
    .SPARE_BIT4 (SPARE_BIT4_REG),
    .SPARE_BIT5 (SPARE_BIT5_REG),
    .SPARE_BIT6 (SPARE_BIT6_REG),
    .SPARE_BIT7 (SPARE_BIT7_REG),
    .SPARE_BIT8 (SPARE_BIT8_REG),
    .SPARE_BYTE0 (SPARE_BYTE0_REG),
    .SPARE_BYTE1 (SPARE_BYTE1_REG),
    .SPARE_BYTE2 (SPARE_BYTE2_REG),
    .SPARE_BYTE3 (SPARE_BYTE3_REG),
    .SPARE_WORD0 (SPARE_WORD0_REG),
    .SPARE_WORD1 (SPARE_WORD1_REG),
    .SPARE_WORD2 (SPARE_WORD2_REG),
    .SPARE_WORD3 (SPARE_WORD3_REG),
    .SRIOV_CAP_ENABLE (SRIOV_CAP_ENABLE_REG),
    .TEST_MODE_PIN_CHAR (TEST_MODE_PIN_CHAR_REG),
    .TL_COMPLETION_RAM_SIZE_16K (TL_COMPLETION_RAM_SIZE_16K_REG),
    .TL_COMPL_TIMEOUT_REG0 (TL_COMPL_TIMEOUT_REG0_REG),
    .TL_COMPL_TIMEOUT_REG1 (TL_COMPL_TIMEOUT_REG1_REG),
    .TL_CREDITS_CD (TL_CREDITS_CD_REG),
    .TL_CREDITS_CH (TL_CREDITS_CH_REG),
    .TL_CREDITS_NPD (TL_CREDITS_NPD_REG),
    .TL_CREDITS_NPH (TL_CREDITS_NPH_REG),
    .TL_CREDITS_PD (TL_CREDITS_PD_REG),
    .TL_CREDITS_PH (TL_CREDITS_PH_REG),
    .TL_ENABLE_MESSAGE_RID_CHECK_ENABLE (TL_ENABLE_MESSAGE_RID_CHECK_ENABLE_REG),
    .TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE (TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE_REG),
    .TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE (TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE_REG),
    .TL_LEGACY_MODE_ENABLE (TL_LEGACY_MODE_ENABLE_REG),
    .TL_PF_ENABLE_REG (TL_PF_ENABLE_REG_REG),
    .TL_TX_MUX_STRICT_PRIORITY (TL_TX_MUX_STRICT_PRIORITY_REG),
    .TWO_LAYER_MODE_DLCMSM_ENABLE (TWO_LAYER_MODE_DLCMSM_ENABLE_REG),
    .TWO_LAYER_MODE_ENABLE (TWO_LAYER_MODE_ENABLE_REG),
    .TWO_LAYER_MODE_WIDTH_256 (TWO_LAYER_MODE_WIDTH_256_REG),
    .VF0_ARI_CAP_NEXTPTR (VF0_ARI_CAP_NEXTPTR_REG),
    .VF0_CAPABILITY_POINTER (VF0_CAPABILITY_POINTER_REG),
    .VF0_MSIX_CAP_PBA_BIR (VF0_MSIX_CAP_PBA_BIR_REG),
    .VF0_MSIX_CAP_PBA_OFFSET (VF0_MSIX_CAP_PBA_OFFSET_REG),
    .VF0_MSIX_CAP_TABLE_BIR (VF0_MSIX_CAP_TABLE_BIR_REG),
    .VF0_MSIX_CAP_TABLE_OFFSET (VF0_MSIX_CAP_TABLE_OFFSET_REG),
    .VF0_MSIX_CAP_TABLE_SIZE (VF0_MSIX_CAP_TABLE_SIZE_REG),
    .VF0_MSI_CAP_MULTIMSGCAP (VF0_MSI_CAP_MULTIMSGCAP_REG),
    .VF0_PM_CAP_ID (VF0_PM_CAP_ID_REG),
    .VF0_PM_CAP_NEXTPTR (VF0_PM_CAP_NEXTPTR_REG),
    .VF0_PM_CAP_VER_ID (VF0_PM_CAP_VER_ID_REG),
    .VF0_TPHR_CAP_DEV_SPECIFIC_MODE (VF0_TPHR_CAP_DEV_SPECIFIC_MODE_REG),
    .VF0_TPHR_CAP_ENABLE (VF0_TPHR_CAP_ENABLE_REG),
    .VF0_TPHR_CAP_INT_VEC_MODE (VF0_TPHR_CAP_INT_VEC_MODE_REG),
    .VF0_TPHR_CAP_NEXTPTR (VF0_TPHR_CAP_NEXTPTR_REG),
    .VF0_TPHR_CAP_ST_MODE_SEL (VF0_TPHR_CAP_ST_MODE_SEL_REG),
    .VF0_TPHR_CAP_ST_TABLE_LOC (VF0_TPHR_CAP_ST_TABLE_LOC_REG),
    .VF0_TPHR_CAP_ST_TABLE_SIZE (VF0_TPHR_CAP_ST_TABLE_SIZE_REG),
    .VF0_TPHR_CAP_VER (VF0_TPHR_CAP_VER_REG),
    .VF1_ARI_CAP_NEXTPTR (VF1_ARI_CAP_NEXTPTR_REG),
    .VF1_MSIX_CAP_PBA_BIR (VF1_MSIX_CAP_PBA_BIR_REG),
    .VF1_MSIX_CAP_PBA_OFFSET (VF1_MSIX_CAP_PBA_OFFSET_REG),
    .VF1_MSIX_CAP_TABLE_BIR (VF1_MSIX_CAP_TABLE_BIR_REG),
    .VF1_MSIX_CAP_TABLE_OFFSET (VF1_MSIX_CAP_TABLE_OFFSET_REG),
    .VF1_MSIX_CAP_TABLE_SIZE (VF1_MSIX_CAP_TABLE_SIZE_REG),
    .VF1_MSI_CAP_MULTIMSGCAP (VF1_MSI_CAP_MULTIMSGCAP_REG),
    .VF1_PM_CAP_ID (VF1_PM_CAP_ID_REG),
    .VF1_PM_CAP_NEXTPTR (VF1_PM_CAP_NEXTPTR_REG),
    .VF1_PM_CAP_VER_ID (VF1_PM_CAP_VER_ID_REG),
    .VF1_TPHR_CAP_DEV_SPECIFIC_MODE (VF1_TPHR_CAP_DEV_SPECIFIC_MODE_REG),
    .VF1_TPHR_CAP_ENABLE (VF1_TPHR_CAP_ENABLE_REG),
    .VF1_TPHR_CAP_INT_VEC_MODE (VF1_TPHR_CAP_INT_VEC_MODE_REG),
    .VF1_TPHR_CAP_NEXTPTR (VF1_TPHR_CAP_NEXTPTR_REG),
    .VF1_TPHR_CAP_ST_MODE_SEL (VF1_TPHR_CAP_ST_MODE_SEL_REG),
    .VF1_TPHR_CAP_ST_TABLE_LOC (VF1_TPHR_CAP_ST_TABLE_LOC_REG),
    .VF1_TPHR_CAP_ST_TABLE_SIZE (VF1_TPHR_CAP_ST_TABLE_SIZE_REG),
    .VF1_TPHR_CAP_VER (VF1_TPHR_CAP_VER_REG),
    .VF2_ARI_CAP_NEXTPTR (VF2_ARI_CAP_NEXTPTR_REG),
    .VF2_MSIX_CAP_PBA_BIR (VF2_MSIX_CAP_PBA_BIR_REG),
    .VF2_MSIX_CAP_PBA_OFFSET (VF2_MSIX_CAP_PBA_OFFSET_REG),
    .VF2_MSIX_CAP_TABLE_BIR (VF2_MSIX_CAP_TABLE_BIR_REG),
    .VF2_MSIX_CAP_TABLE_OFFSET (VF2_MSIX_CAP_TABLE_OFFSET_REG),
    .VF2_MSIX_CAP_TABLE_SIZE (VF2_MSIX_CAP_TABLE_SIZE_REG),
    .VF2_MSI_CAP_MULTIMSGCAP (VF2_MSI_CAP_MULTIMSGCAP_REG),
    .VF2_PM_CAP_ID (VF2_PM_CAP_ID_REG),
    .VF2_PM_CAP_NEXTPTR (VF2_PM_CAP_NEXTPTR_REG),
    .VF2_PM_CAP_VER_ID (VF2_PM_CAP_VER_ID_REG),
    .VF2_TPHR_CAP_DEV_SPECIFIC_MODE (VF2_TPHR_CAP_DEV_SPECIFIC_MODE_REG),
    .VF2_TPHR_CAP_ENABLE (VF2_TPHR_CAP_ENABLE_REG),
    .VF2_TPHR_CAP_INT_VEC_MODE (VF2_TPHR_CAP_INT_VEC_MODE_REG),
    .VF2_TPHR_CAP_NEXTPTR (VF2_TPHR_CAP_NEXTPTR_REG),
    .VF2_TPHR_CAP_ST_MODE_SEL (VF2_TPHR_CAP_ST_MODE_SEL_REG),
    .VF2_TPHR_CAP_ST_TABLE_LOC (VF2_TPHR_CAP_ST_TABLE_LOC_REG),
    .VF2_TPHR_CAP_ST_TABLE_SIZE (VF2_TPHR_CAP_ST_TABLE_SIZE_REG),
    .VF2_TPHR_CAP_VER (VF2_TPHR_CAP_VER_REG),
    .VF3_ARI_CAP_NEXTPTR (VF3_ARI_CAP_NEXTPTR_REG),
    .VF3_MSIX_CAP_PBA_BIR (VF3_MSIX_CAP_PBA_BIR_REG),
    .VF3_MSIX_CAP_PBA_OFFSET (VF3_MSIX_CAP_PBA_OFFSET_REG),
    .VF3_MSIX_CAP_TABLE_BIR (VF3_MSIX_CAP_TABLE_BIR_REG),
    .VF3_MSIX_CAP_TABLE_OFFSET (VF3_MSIX_CAP_TABLE_OFFSET_REG),
    .VF3_MSIX_CAP_TABLE_SIZE (VF3_MSIX_CAP_TABLE_SIZE_REG),
    .VF3_MSI_CAP_MULTIMSGCAP (VF3_MSI_CAP_MULTIMSGCAP_REG),
    .VF3_PM_CAP_ID (VF3_PM_CAP_ID_REG),
    .VF3_PM_CAP_NEXTPTR (VF3_PM_CAP_NEXTPTR_REG),
    .VF3_PM_CAP_VER_ID (VF3_PM_CAP_VER_ID_REG),
    .VF3_TPHR_CAP_DEV_SPECIFIC_MODE (VF3_TPHR_CAP_DEV_SPECIFIC_MODE_REG),
    .VF3_TPHR_CAP_ENABLE (VF3_TPHR_CAP_ENABLE_REG),
    .VF3_TPHR_CAP_INT_VEC_MODE (VF3_TPHR_CAP_INT_VEC_MODE_REG),
    .VF3_TPHR_CAP_NEXTPTR (VF3_TPHR_CAP_NEXTPTR_REG),
    .VF3_TPHR_CAP_ST_MODE_SEL (VF3_TPHR_CAP_ST_MODE_SEL_REG),
    .VF3_TPHR_CAP_ST_TABLE_LOC (VF3_TPHR_CAP_ST_TABLE_LOC_REG),
    .VF3_TPHR_CAP_ST_TABLE_SIZE (VF3_TPHR_CAP_ST_TABLE_SIZE_REG),
    .VF3_TPHR_CAP_VER (VF3_TPHR_CAP_VER_REG),
    .VF4_ARI_CAP_NEXTPTR (VF4_ARI_CAP_NEXTPTR_REG),
    .VF4_MSIX_CAP_PBA_BIR (VF4_MSIX_CAP_PBA_BIR_REG),
    .VF4_MSIX_CAP_PBA_OFFSET (VF4_MSIX_CAP_PBA_OFFSET_REG),
    .VF4_MSIX_CAP_TABLE_BIR (VF4_MSIX_CAP_TABLE_BIR_REG),
    .VF4_MSIX_CAP_TABLE_OFFSET (VF4_MSIX_CAP_TABLE_OFFSET_REG),
    .VF4_MSIX_CAP_TABLE_SIZE (VF4_MSIX_CAP_TABLE_SIZE_REG),
    .VF4_MSI_CAP_MULTIMSGCAP (VF4_MSI_CAP_MULTIMSGCAP_REG),
    .VF4_PM_CAP_ID (VF4_PM_CAP_ID_REG),
    .VF4_PM_CAP_NEXTPTR (VF4_PM_CAP_NEXTPTR_REG),
    .VF4_PM_CAP_VER_ID (VF4_PM_CAP_VER_ID_REG),
    .VF4_TPHR_CAP_DEV_SPECIFIC_MODE (VF4_TPHR_CAP_DEV_SPECIFIC_MODE_REG),
    .VF4_TPHR_CAP_ENABLE (VF4_TPHR_CAP_ENABLE_REG),
    .VF4_TPHR_CAP_INT_VEC_MODE (VF4_TPHR_CAP_INT_VEC_MODE_REG),
    .VF4_TPHR_CAP_NEXTPTR (VF4_TPHR_CAP_NEXTPTR_REG),
    .VF4_TPHR_CAP_ST_MODE_SEL (VF4_TPHR_CAP_ST_MODE_SEL_REG),
    .VF4_TPHR_CAP_ST_TABLE_LOC (VF4_TPHR_CAP_ST_TABLE_LOC_REG),
    .VF4_TPHR_CAP_ST_TABLE_SIZE (VF4_TPHR_CAP_ST_TABLE_SIZE_REG),
    .VF4_TPHR_CAP_VER (VF4_TPHR_CAP_VER_REG),
    .VF5_ARI_CAP_NEXTPTR (VF5_ARI_CAP_NEXTPTR_REG),
    .VF5_MSIX_CAP_PBA_BIR (VF5_MSIX_CAP_PBA_BIR_REG),
    .VF5_MSIX_CAP_PBA_OFFSET (VF5_MSIX_CAP_PBA_OFFSET_REG),
    .VF5_MSIX_CAP_TABLE_BIR (VF5_MSIX_CAP_TABLE_BIR_REG),
    .VF5_MSIX_CAP_TABLE_OFFSET (VF5_MSIX_CAP_TABLE_OFFSET_REG),
    .VF5_MSIX_CAP_TABLE_SIZE (VF5_MSIX_CAP_TABLE_SIZE_REG),
    .VF5_MSI_CAP_MULTIMSGCAP (VF5_MSI_CAP_MULTIMSGCAP_REG),
    .VF5_PM_CAP_ID (VF5_PM_CAP_ID_REG),
    .VF5_PM_CAP_NEXTPTR (VF5_PM_CAP_NEXTPTR_REG),
    .VF5_PM_CAP_VER_ID (VF5_PM_CAP_VER_ID_REG),
    .VF5_TPHR_CAP_DEV_SPECIFIC_MODE (VF5_TPHR_CAP_DEV_SPECIFIC_MODE_REG),
    .VF5_TPHR_CAP_ENABLE (VF5_TPHR_CAP_ENABLE_REG),
    .VF5_TPHR_CAP_INT_VEC_MODE (VF5_TPHR_CAP_INT_VEC_MODE_REG),
    .VF5_TPHR_CAP_NEXTPTR (VF5_TPHR_CAP_NEXTPTR_REG),
    .VF5_TPHR_CAP_ST_MODE_SEL (VF5_TPHR_CAP_ST_MODE_SEL_REG),
    .VF5_TPHR_CAP_ST_TABLE_LOC (VF5_TPHR_CAP_ST_TABLE_LOC_REG),
    .VF5_TPHR_CAP_ST_TABLE_SIZE (VF5_TPHR_CAP_ST_TABLE_SIZE_REG),
    .VF5_TPHR_CAP_VER (VF5_TPHR_CAP_VER_REG),
    .VF6_ARI_CAP_NEXTPTR (VF6_ARI_CAP_NEXTPTR_REG),
    .VF6_MSIX_CAP_PBA_BIR (VF6_MSIX_CAP_PBA_BIR_REG),
    .VF6_MSIX_CAP_PBA_OFFSET (VF6_MSIX_CAP_PBA_OFFSET_REG),
    .VF6_MSIX_CAP_TABLE_BIR (VF6_MSIX_CAP_TABLE_BIR_REG),
    .VF6_MSIX_CAP_TABLE_OFFSET (VF6_MSIX_CAP_TABLE_OFFSET_REG),
    .VF6_MSIX_CAP_TABLE_SIZE (VF6_MSIX_CAP_TABLE_SIZE_REG),
    .VF6_MSI_CAP_MULTIMSGCAP (VF6_MSI_CAP_MULTIMSGCAP_REG),
    .VF6_PM_CAP_ID (VF6_PM_CAP_ID_REG),
    .VF6_PM_CAP_NEXTPTR (VF6_PM_CAP_NEXTPTR_REG),
    .VF6_PM_CAP_VER_ID (VF6_PM_CAP_VER_ID_REG),
    .VF6_TPHR_CAP_DEV_SPECIFIC_MODE (VF6_TPHR_CAP_DEV_SPECIFIC_MODE_REG),
    .VF6_TPHR_CAP_ENABLE (VF6_TPHR_CAP_ENABLE_REG),
    .VF6_TPHR_CAP_INT_VEC_MODE (VF6_TPHR_CAP_INT_VEC_MODE_REG),
    .VF6_TPHR_CAP_NEXTPTR (VF6_TPHR_CAP_NEXTPTR_REG),
    .VF6_TPHR_CAP_ST_MODE_SEL (VF6_TPHR_CAP_ST_MODE_SEL_REG),
    .VF6_TPHR_CAP_ST_TABLE_LOC (VF6_TPHR_CAP_ST_TABLE_LOC_REG),
    .VF6_TPHR_CAP_ST_TABLE_SIZE (VF6_TPHR_CAP_ST_TABLE_SIZE_REG),
    .VF6_TPHR_CAP_VER (VF6_TPHR_CAP_VER_REG),
    .VF7_ARI_CAP_NEXTPTR (VF7_ARI_CAP_NEXTPTR_REG),
    .VF7_MSIX_CAP_PBA_BIR (VF7_MSIX_CAP_PBA_BIR_REG),
    .VF7_MSIX_CAP_PBA_OFFSET (VF7_MSIX_CAP_PBA_OFFSET_REG),
    .VF7_MSIX_CAP_TABLE_BIR (VF7_MSIX_CAP_TABLE_BIR_REG),
    .VF7_MSIX_CAP_TABLE_OFFSET (VF7_MSIX_CAP_TABLE_OFFSET_REG),
    .VF7_MSIX_CAP_TABLE_SIZE (VF7_MSIX_CAP_TABLE_SIZE_REG),
    .VF7_MSI_CAP_MULTIMSGCAP (VF7_MSI_CAP_MULTIMSGCAP_REG),
    .VF7_PM_CAP_ID (VF7_PM_CAP_ID_REG),
    .VF7_PM_CAP_NEXTPTR (VF7_PM_CAP_NEXTPTR_REG),
    .VF7_PM_CAP_VER_ID (VF7_PM_CAP_VER_ID_REG),
    .VF7_TPHR_CAP_DEV_SPECIFIC_MODE (VF7_TPHR_CAP_DEV_SPECIFIC_MODE_REG),
    .VF7_TPHR_CAP_ENABLE (VF7_TPHR_CAP_ENABLE_REG),
    .VF7_TPHR_CAP_INT_VEC_MODE (VF7_TPHR_CAP_INT_VEC_MODE_REG),
    .VF7_TPHR_CAP_NEXTPTR (VF7_TPHR_CAP_NEXTPTR_REG),
    .VF7_TPHR_CAP_ST_MODE_SEL (VF7_TPHR_CAP_ST_MODE_SEL_REG),
    .VF7_TPHR_CAP_ST_TABLE_LOC (VF7_TPHR_CAP_ST_TABLE_LOC_REG),
    .VF7_TPHR_CAP_ST_TABLE_SIZE (VF7_TPHR_CAP_ST_TABLE_SIZE_REG),
    .VF7_TPHR_CAP_VER (VF7_TPHR_CAP_VER_REG),
    .CFGCURRENTSPEED (CFGCURRENTSPEED_out),
    .CFGDPASUBSTATECHANGE (CFGDPASUBSTATECHANGE_out),
    .CFGERRCOROUT (CFGERRCOROUT_out),
    .CFGERRFATALOUT (CFGERRFATALOUT_out),
    .CFGERRNONFATALOUT (CFGERRNONFATALOUT_out),
    .CFGEXTFUNCTIONNUMBER (CFGEXTFUNCTIONNUMBER_out),
    .CFGEXTREADRECEIVED (CFGEXTREADRECEIVED_out),
    .CFGEXTREGISTERNUMBER (CFGEXTREGISTERNUMBER_out),
    .CFGEXTWRITEBYTEENABLE (CFGEXTWRITEBYTEENABLE_out),
    .CFGEXTWRITEDATA (CFGEXTWRITEDATA_out),
    .CFGEXTWRITERECEIVED (CFGEXTWRITERECEIVED_out),
    .CFGFCCPLD (CFGFCCPLD_out),
    .CFGFCCPLH (CFGFCCPLH_out),
    .CFGFCNPD (CFGFCNPD_out),
    .CFGFCNPH (CFGFCNPH_out),
    .CFGFCPD (CFGFCPD_out),
    .CFGFCPH (CFGFCPH_out),
    .CFGFLRINPROCESS (CFGFLRINPROCESS_out),
    .CFGFUNCTIONPOWERSTATE (CFGFUNCTIONPOWERSTATE_out),
    .CFGFUNCTIONSTATUS (CFGFUNCTIONSTATUS_out),
    .CFGHOTRESETOUT (CFGHOTRESETOUT_out),
    .CFGINTERRUPTMSIDATA (CFGINTERRUPTMSIDATA_out),
    .CFGINTERRUPTMSIENABLE (CFGINTERRUPTMSIENABLE_out),
    .CFGINTERRUPTMSIFAIL (CFGINTERRUPTMSIFAIL_out),
    .CFGINTERRUPTMSIMASKUPDATE (CFGINTERRUPTMSIMASKUPDATE_out),
    .CFGINTERRUPTMSIMMENABLE (CFGINTERRUPTMSIMMENABLE_out),
    .CFGINTERRUPTMSISENT (CFGINTERRUPTMSISENT_out),
    .CFGINTERRUPTMSIVFENABLE (CFGINTERRUPTMSIVFENABLE_out),
    .CFGINTERRUPTMSIXENABLE (CFGINTERRUPTMSIXENABLE_out),
    .CFGINTERRUPTMSIXFAIL (CFGINTERRUPTMSIXFAIL_out),
    .CFGINTERRUPTMSIXMASK (CFGINTERRUPTMSIXMASK_out),
    .CFGINTERRUPTMSIXSENT (CFGINTERRUPTMSIXSENT_out),
    .CFGINTERRUPTMSIXVFENABLE (CFGINTERRUPTMSIXVFENABLE_out),
    .CFGINTERRUPTMSIXVFMASK (CFGINTERRUPTMSIXVFMASK_out),
    .CFGINTERRUPTSENT (CFGINTERRUPTSENT_out),
    .CFGLINKPOWERSTATE (CFGLINKPOWERSTATE_out),
    .CFGLOCALERROR (CFGLOCALERROR_out),
    .CFGLTRENABLE (CFGLTRENABLE_out),
    .CFGLTSSMSTATE (CFGLTSSMSTATE_out),
    .CFGMAXPAYLOAD (CFGMAXPAYLOAD_out),
    .CFGMAXREADREQ (CFGMAXREADREQ_out),
    .CFGMGMTREADDATA (CFGMGMTREADDATA_out),
    .CFGMGMTREADWRITEDONE (CFGMGMTREADWRITEDONE_out),
    .CFGMSGRECEIVED (CFGMSGRECEIVED_out),
    .CFGMSGRECEIVEDDATA (CFGMSGRECEIVEDDATA_out),
    .CFGMSGRECEIVEDTYPE (CFGMSGRECEIVEDTYPE_out),
    .CFGMSGTRANSMITDONE (CFGMSGTRANSMITDONE_out),
    .CFGNEGOTIATEDWIDTH (CFGNEGOTIATEDWIDTH_out),
    .CFGOBFFENABLE (CFGOBFFENABLE_out),
    .CFGPERFUNCSTATUSDATA (CFGPERFUNCSTATUSDATA_out),
    .CFGPERFUNCTIONUPDATEDONE (CFGPERFUNCTIONUPDATEDONE_out),
    .CFGPHYLINKDOWN (CFGPHYLINKDOWN_out),
    .CFGPHYLINKSTATUS (CFGPHYLINKSTATUS_out),
    .CFGPLSTATUSCHANGE (CFGPLSTATUSCHANGE_out),
    .CFGPOWERSTATECHANGEINTERRUPT (CFGPOWERSTATECHANGEINTERRUPT_out),
    .CFGRCBSTATUS (CFGRCBSTATUS_out),
    .CFGTPHFUNCTIONNUM (CFGTPHFUNCTIONNUM_out),
    .CFGTPHREQUESTERENABLE (CFGTPHREQUESTERENABLE_out),
    .CFGTPHSTMODE (CFGTPHSTMODE_out),
    .CFGTPHSTTADDRESS (CFGTPHSTTADDRESS_out),
    .CFGTPHSTTREADENABLE (CFGTPHSTTREADENABLE_out),
    .CFGTPHSTTWRITEBYTEVALID (CFGTPHSTTWRITEBYTEVALID_out),
    .CFGTPHSTTWRITEDATA (CFGTPHSTTWRITEDATA_out),
    .CFGTPHSTTWRITEENABLE (CFGTPHSTTWRITEENABLE_out),
    .CFGVFFLRINPROCESS (CFGVFFLRINPROCESS_out),
    .CFGVFPOWERSTATE (CFGVFPOWERSTATE_out),
    .CFGVFSTATUS (CFGVFSTATUS_out),
    .CFGVFTPHREQUESTERENABLE (CFGVFTPHREQUESTERENABLE_out),
    .CFGVFTPHSTMODE (CFGVFTPHSTMODE_out),
    .CONFMCAPDESIGNSWITCH (CONFMCAPDESIGNSWITCH_out),
    .CONFMCAPEOS (CONFMCAPEOS_out),
    .CONFMCAPINUSEBYPCIE (CONFMCAPINUSEBYPCIE_out),
    .CONFREQREADY (CONFREQREADY_out),
    .CONFRESPRDATA (CONFRESPRDATA_out),
    .CONFRESPVALID (CONFRESPVALID_out),
    .DBGDATAOUT (DBGDATAOUT_out),
    .DBGMCAPCSB (DBGMCAPCSB_out),
    .DBGMCAPDATA (DBGMCAPDATA_out),
    .DBGMCAPEOS (DBGMCAPEOS_out),
    .DBGMCAPERROR (DBGMCAPERROR_out),
    .DBGMCAPMODE (DBGMCAPMODE_out),
    .DBGMCAPRDATAVALID (DBGMCAPRDATAVALID_out),
    .DBGMCAPRDWRB (DBGMCAPRDWRB_out),
    .DBGMCAPRESET (DBGMCAPRESET_out),
    .DBGPLDATABLOCKRECEIVEDAFTEREDS (DBGPLDATABLOCKRECEIVEDAFTEREDS_out),
    .DBGPLGEN3FRAMINGERRORDETECTED (DBGPLGEN3FRAMINGERRORDETECTED_out),
    .DBGPLGEN3SYNCHEADERERRORDETECTED (DBGPLGEN3SYNCHEADERERRORDETECTED_out),
    .DBGPLINFERREDRXELECTRICALIDLE (DBGPLINFERREDRXELECTRICALIDLE_out),
    .DRPDO (DRPDO_out),
    .DRPRDY (DRPRDY_out),
    .LL2LMMASTERTLPSENT0 (LL2LMMASTERTLPSENT0_out),
    .LL2LMMASTERTLPSENT1 (LL2LMMASTERTLPSENT1_out),
    .LL2LMMASTERTLPSENTTLPID0 (LL2LMMASTERTLPSENTTLPID0_out),
    .LL2LMMASTERTLPSENTTLPID1 (LL2LMMASTERTLPSENTTLPID1_out),
    .LL2LMMAXISRXTDATA (LL2LMMAXISRXTDATA_out),
    .LL2LMMAXISRXTUSER (LL2LMMAXISRXTUSER_out),
    .LL2LMMAXISRXTVALID (LL2LMMAXISRXTVALID_out),
    .LL2LMSAXISTXTREADY (LL2LMSAXISTXTREADY_out),
    .MAXISCQTDATA (MAXISCQTDATA_out),
    .MAXISCQTKEEP (MAXISCQTKEEP_out),
    .MAXISCQTLAST (MAXISCQTLAST_out),
    .MAXISCQTUSER (MAXISCQTUSER_out),
    .MAXISCQTVALID (MAXISCQTVALID_out),
    .MAXISRCTDATA (MAXISRCTDATA_out),
    .MAXISRCTKEEP (MAXISRCTKEEP_out),
    .MAXISRCTLAST (MAXISRCTLAST_out),
    .MAXISRCTUSER (MAXISRCTUSER_out),
    .MAXISRCTVALID (MAXISRCTVALID_out),
    .MICOMPLETIONRAMREADADDRESSAL (MICOMPLETIONRAMREADADDRESSAL_out),
    .MICOMPLETIONRAMREADADDRESSAU (MICOMPLETIONRAMREADADDRESSAU_out),
    .MICOMPLETIONRAMREADADDRESSBL (MICOMPLETIONRAMREADADDRESSBL_out),
    .MICOMPLETIONRAMREADADDRESSBU (MICOMPLETIONRAMREADADDRESSBU_out),
    .MICOMPLETIONRAMREADENABLEL (MICOMPLETIONRAMREADENABLEL_out),
    .MICOMPLETIONRAMREADENABLEU (MICOMPLETIONRAMREADENABLEU_out),
    .MICOMPLETIONRAMWRITEADDRESSAL (MICOMPLETIONRAMWRITEADDRESSAL_out),
    .MICOMPLETIONRAMWRITEADDRESSAU (MICOMPLETIONRAMWRITEADDRESSAU_out),
    .MICOMPLETIONRAMWRITEADDRESSBL (MICOMPLETIONRAMWRITEADDRESSBL_out),
    .MICOMPLETIONRAMWRITEADDRESSBU (MICOMPLETIONRAMWRITEADDRESSBU_out),
    .MICOMPLETIONRAMWRITEDATAL (MICOMPLETIONRAMWRITEDATAL_out),
    .MICOMPLETIONRAMWRITEDATAU (MICOMPLETIONRAMWRITEDATAU_out),
    .MICOMPLETIONRAMWRITEENABLEL (MICOMPLETIONRAMWRITEENABLEL_out),
    .MICOMPLETIONRAMWRITEENABLEU (MICOMPLETIONRAMWRITEENABLEU_out),
    .MIREPLAYRAMADDRESS (MIREPLAYRAMADDRESS_out),
    .MIREPLAYRAMREADENABLE (MIREPLAYRAMREADENABLE_out),
    .MIREPLAYRAMWRITEDATA (MIREPLAYRAMWRITEDATA_out),
    .MIREPLAYRAMWRITEENABLE (MIREPLAYRAMWRITEENABLE_out),
    .MIREQUESTRAMREADADDRESSA (MIREQUESTRAMREADADDRESSA_out),
    .MIREQUESTRAMREADADDRESSB (MIREQUESTRAMREADADDRESSB_out),
    .MIREQUESTRAMREADENABLE (MIREQUESTRAMREADENABLE_out),
    .MIREQUESTRAMWRITEADDRESSA (MIREQUESTRAMWRITEADDRESSA_out),
    .MIREQUESTRAMWRITEADDRESSB (MIREQUESTRAMWRITEADDRESSB_out),
    .MIREQUESTRAMWRITEDATA (MIREQUESTRAMWRITEDATA_out),
    .MIREQUESTRAMWRITEENABLE (MIREQUESTRAMWRITEENABLE_out),
    .PCIECQNPREQCOUNT (PCIECQNPREQCOUNT_out),
    .PCIEPERST0B (PCIEPERST0B_out),
    .PCIEPERST1B (PCIEPERST1B_out),
    .PCIERQSEQNUM (PCIERQSEQNUM_out),
    .PCIERQSEQNUMVLD (PCIERQSEQNUMVLD_out),
    .PCIERQTAG (PCIERQTAG_out),
    .PCIERQTAGAV (PCIERQTAGAV_out),
    .PCIERQTAGVLD (PCIERQTAGVLD_out),
    .PCIETFCNPDAV (PCIETFCNPDAV_out),
    .PCIETFCNPHAV (PCIETFCNPHAV_out),
    .PIPERX0EQCONTROL (PIPERX0EQCONTROL_out),
    .PIPERX0EQLPLFFS (PIPERX0EQLPLFFS_out),
    .PIPERX0EQLPTXPRESET (PIPERX0EQLPTXPRESET_out),
    .PIPERX0EQPRESET (PIPERX0EQPRESET_out),
    .PIPERX0POLARITY (PIPERX0POLARITY_out),
    .PIPERX1EQCONTROL (PIPERX1EQCONTROL_out),
    .PIPERX1EQLPLFFS (PIPERX1EQLPLFFS_out),
    .PIPERX1EQLPTXPRESET (PIPERX1EQLPTXPRESET_out),
    .PIPERX1EQPRESET (PIPERX1EQPRESET_out),
    .PIPERX1POLARITY (PIPERX1POLARITY_out),
    .PIPERX2EQCONTROL (PIPERX2EQCONTROL_out),
    .PIPERX2EQLPLFFS (PIPERX2EQLPLFFS_out),
    .PIPERX2EQLPTXPRESET (PIPERX2EQLPTXPRESET_out),
    .PIPERX2EQPRESET (PIPERX2EQPRESET_out),
    .PIPERX2POLARITY (PIPERX2POLARITY_out),
    .PIPERX3EQCONTROL (PIPERX3EQCONTROL_out),
    .PIPERX3EQLPLFFS (PIPERX3EQLPLFFS_out),
    .PIPERX3EQLPTXPRESET (PIPERX3EQLPTXPRESET_out),
    .PIPERX3EQPRESET (PIPERX3EQPRESET_out),
    .PIPERX3POLARITY (PIPERX3POLARITY_out),
    .PIPERX4EQCONTROL (PIPERX4EQCONTROL_out),
    .PIPERX4EQLPLFFS (PIPERX4EQLPLFFS_out),
    .PIPERX4EQLPTXPRESET (PIPERX4EQLPTXPRESET_out),
    .PIPERX4EQPRESET (PIPERX4EQPRESET_out),
    .PIPERX4POLARITY (PIPERX4POLARITY_out),
    .PIPERX5EQCONTROL (PIPERX5EQCONTROL_out),
    .PIPERX5EQLPLFFS (PIPERX5EQLPLFFS_out),
    .PIPERX5EQLPTXPRESET (PIPERX5EQLPTXPRESET_out),
    .PIPERX5EQPRESET (PIPERX5EQPRESET_out),
    .PIPERX5POLARITY (PIPERX5POLARITY_out),
    .PIPERX6EQCONTROL (PIPERX6EQCONTROL_out),
    .PIPERX6EQLPLFFS (PIPERX6EQLPLFFS_out),
    .PIPERX6EQLPTXPRESET (PIPERX6EQLPTXPRESET_out),
    .PIPERX6EQPRESET (PIPERX6EQPRESET_out),
    .PIPERX6POLARITY (PIPERX6POLARITY_out),
    .PIPERX7EQCONTROL (PIPERX7EQCONTROL_out),
    .PIPERX7EQLPLFFS (PIPERX7EQLPLFFS_out),
    .PIPERX7EQLPTXPRESET (PIPERX7EQLPTXPRESET_out),
    .PIPERX7EQPRESET (PIPERX7EQPRESET_out),
    .PIPERX7POLARITY (PIPERX7POLARITY_out),
    .PIPETX0CHARISK (PIPETX0CHARISK_out),
    .PIPETX0COMPLIANCE (PIPETX0COMPLIANCE_out),
    .PIPETX0DATA (PIPETX0DATA_out),
    .PIPETX0DATAVALID (PIPETX0DATAVALID_out),
    .PIPETX0DEEMPH (PIPETX0DEEMPH_out),
    .PIPETX0ELECIDLE (PIPETX0ELECIDLE_out),
    .PIPETX0EQCONTROL (PIPETX0EQCONTROL_out),
    .PIPETX0EQDEEMPH (PIPETX0EQDEEMPH_out),
    .PIPETX0EQPRESET (PIPETX0EQPRESET_out),
    .PIPETX0MARGIN (PIPETX0MARGIN_out),
    .PIPETX0POWERDOWN (PIPETX0POWERDOWN_out),
    .PIPETX0RATE (PIPETX0RATE_out),
    .PIPETX0RCVRDET (PIPETX0RCVRDET_out),
    .PIPETX0RESET (PIPETX0RESET_out),
    .PIPETX0STARTBLOCK (PIPETX0STARTBLOCK_out),
    .PIPETX0SWING (PIPETX0SWING_out),
    .PIPETX0SYNCHEADER (PIPETX0SYNCHEADER_out),
    .PIPETX1CHARISK (PIPETX1CHARISK_out),
    .PIPETX1COMPLIANCE (PIPETX1COMPLIANCE_out),
    .PIPETX1DATA (PIPETX1DATA_out),
    .PIPETX1DATAVALID (PIPETX1DATAVALID_out),
    .PIPETX1DEEMPH (PIPETX1DEEMPH_out),
    .PIPETX1ELECIDLE (PIPETX1ELECIDLE_out),
    .PIPETX1EQCONTROL (PIPETX1EQCONTROL_out),
    .PIPETX1EQDEEMPH (PIPETX1EQDEEMPH_out),
    .PIPETX1EQPRESET (PIPETX1EQPRESET_out),
    .PIPETX1MARGIN (PIPETX1MARGIN_out),
    .PIPETX1POWERDOWN (PIPETX1POWERDOWN_out),
    .PIPETX1RATE (PIPETX1RATE_out),
    .PIPETX1RCVRDET (PIPETX1RCVRDET_out),
    .PIPETX1RESET (PIPETX1RESET_out),
    .PIPETX1STARTBLOCK (PIPETX1STARTBLOCK_out),
    .PIPETX1SWING (PIPETX1SWING_out),
    .PIPETX1SYNCHEADER (PIPETX1SYNCHEADER_out),
    .PIPETX2CHARISK (PIPETX2CHARISK_out),
    .PIPETX2COMPLIANCE (PIPETX2COMPLIANCE_out),
    .PIPETX2DATA (PIPETX2DATA_out),
    .PIPETX2DATAVALID (PIPETX2DATAVALID_out),
    .PIPETX2DEEMPH (PIPETX2DEEMPH_out),
    .PIPETX2ELECIDLE (PIPETX2ELECIDLE_out),
    .PIPETX2EQCONTROL (PIPETX2EQCONTROL_out),
    .PIPETX2EQDEEMPH (PIPETX2EQDEEMPH_out),
    .PIPETX2EQPRESET (PIPETX2EQPRESET_out),
    .PIPETX2MARGIN (PIPETX2MARGIN_out),
    .PIPETX2POWERDOWN (PIPETX2POWERDOWN_out),
    .PIPETX2RATE (PIPETX2RATE_out),
    .PIPETX2RCVRDET (PIPETX2RCVRDET_out),
    .PIPETX2RESET (PIPETX2RESET_out),
    .PIPETX2STARTBLOCK (PIPETX2STARTBLOCK_out),
    .PIPETX2SWING (PIPETX2SWING_out),
    .PIPETX2SYNCHEADER (PIPETX2SYNCHEADER_out),
    .PIPETX3CHARISK (PIPETX3CHARISK_out),
    .PIPETX3COMPLIANCE (PIPETX3COMPLIANCE_out),
    .PIPETX3DATA (PIPETX3DATA_out),
    .PIPETX3DATAVALID (PIPETX3DATAVALID_out),
    .PIPETX3DEEMPH (PIPETX3DEEMPH_out),
    .PIPETX3ELECIDLE (PIPETX3ELECIDLE_out),
    .PIPETX3EQCONTROL (PIPETX3EQCONTROL_out),
    .PIPETX3EQDEEMPH (PIPETX3EQDEEMPH_out),
    .PIPETX3EQPRESET (PIPETX3EQPRESET_out),
    .PIPETX3MARGIN (PIPETX3MARGIN_out),
    .PIPETX3POWERDOWN (PIPETX3POWERDOWN_out),
    .PIPETX3RATE (PIPETX3RATE_out),
    .PIPETX3RCVRDET (PIPETX3RCVRDET_out),
    .PIPETX3RESET (PIPETX3RESET_out),
    .PIPETX3STARTBLOCK (PIPETX3STARTBLOCK_out),
    .PIPETX3SWING (PIPETX3SWING_out),
    .PIPETX3SYNCHEADER (PIPETX3SYNCHEADER_out),
    .PIPETX4CHARISK (PIPETX4CHARISK_out),
    .PIPETX4COMPLIANCE (PIPETX4COMPLIANCE_out),
    .PIPETX4DATA (PIPETX4DATA_out),
    .PIPETX4DATAVALID (PIPETX4DATAVALID_out),
    .PIPETX4DEEMPH (PIPETX4DEEMPH_out),
    .PIPETX4ELECIDLE (PIPETX4ELECIDLE_out),
    .PIPETX4EQCONTROL (PIPETX4EQCONTROL_out),
    .PIPETX4EQDEEMPH (PIPETX4EQDEEMPH_out),
    .PIPETX4EQPRESET (PIPETX4EQPRESET_out),
    .PIPETX4MARGIN (PIPETX4MARGIN_out),
    .PIPETX4POWERDOWN (PIPETX4POWERDOWN_out),
    .PIPETX4RATE (PIPETX4RATE_out),
    .PIPETX4RCVRDET (PIPETX4RCVRDET_out),
    .PIPETX4RESET (PIPETX4RESET_out),
    .PIPETX4STARTBLOCK (PIPETX4STARTBLOCK_out),
    .PIPETX4SWING (PIPETX4SWING_out),
    .PIPETX4SYNCHEADER (PIPETX4SYNCHEADER_out),
    .PIPETX5CHARISK (PIPETX5CHARISK_out),
    .PIPETX5COMPLIANCE (PIPETX5COMPLIANCE_out),
    .PIPETX5DATA (PIPETX5DATA_out),
    .PIPETX5DATAVALID (PIPETX5DATAVALID_out),
    .PIPETX5DEEMPH (PIPETX5DEEMPH_out),
    .PIPETX5ELECIDLE (PIPETX5ELECIDLE_out),
    .PIPETX5EQCONTROL (PIPETX5EQCONTROL_out),
    .PIPETX5EQDEEMPH (PIPETX5EQDEEMPH_out),
    .PIPETX5EQPRESET (PIPETX5EQPRESET_out),
    .PIPETX5MARGIN (PIPETX5MARGIN_out),
    .PIPETX5POWERDOWN (PIPETX5POWERDOWN_out),
    .PIPETX5RATE (PIPETX5RATE_out),
    .PIPETX5RCVRDET (PIPETX5RCVRDET_out),
    .PIPETX5RESET (PIPETX5RESET_out),
    .PIPETX5STARTBLOCK (PIPETX5STARTBLOCK_out),
    .PIPETX5SWING (PIPETX5SWING_out),
    .PIPETX5SYNCHEADER (PIPETX5SYNCHEADER_out),
    .PIPETX6CHARISK (PIPETX6CHARISK_out),
    .PIPETX6COMPLIANCE (PIPETX6COMPLIANCE_out),
    .PIPETX6DATA (PIPETX6DATA_out),
    .PIPETX6DATAVALID (PIPETX6DATAVALID_out),
    .PIPETX6DEEMPH (PIPETX6DEEMPH_out),
    .PIPETX6ELECIDLE (PIPETX6ELECIDLE_out),
    .PIPETX6EQCONTROL (PIPETX6EQCONTROL_out),
    .PIPETX6EQDEEMPH (PIPETX6EQDEEMPH_out),
    .PIPETX6EQPRESET (PIPETX6EQPRESET_out),
    .PIPETX6MARGIN (PIPETX6MARGIN_out),
    .PIPETX6POWERDOWN (PIPETX6POWERDOWN_out),
    .PIPETX6RATE (PIPETX6RATE_out),
    .PIPETX6RCVRDET (PIPETX6RCVRDET_out),
    .PIPETX6RESET (PIPETX6RESET_out),
    .PIPETX6STARTBLOCK (PIPETX6STARTBLOCK_out),
    .PIPETX6SWING (PIPETX6SWING_out),
    .PIPETX6SYNCHEADER (PIPETX6SYNCHEADER_out),
    .PIPETX7CHARISK (PIPETX7CHARISK_out),
    .PIPETX7COMPLIANCE (PIPETX7COMPLIANCE_out),
    .PIPETX7DATA (PIPETX7DATA_out),
    .PIPETX7DATAVALID (PIPETX7DATAVALID_out),
    .PIPETX7DEEMPH (PIPETX7DEEMPH_out),
    .PIPETX7ELECIDLE (PIPETX7ELECIDLE_out),
    .PIPETX7EQCONTROL (PIPETX7EQCONTROL_out),
    .PIPETX7EQDEEMPH (PIPETX7EQDEEMPH_out),
    .PIPETX7EQPRESET (PIPETX7EQPRESET_out),
    .PIPETX7MARGIN (PIPETX7MARGIN_out),
    .PIPETX7POWERDOWN (PIPETX7POWERDOWN_out),
    .PIPETX7RATE (PIPETX7RATE_out),
    .PIPETX7RCVRDET (PIPETX7RCVRDET_out),
    .PIPETX7RESET (PIPETX7RESET_out),
    .PIPETX7STARTBLOCK (PIPETX7STARTBLOCK_out),
    .PIPETX7SWING (PIPETX7SWING_out),
    .PIPETX7SYNCHEADER (PIPETX7SYNCHEADER_out),
    .PLEQINPROGRESS (PLEQINPROGRESS_out),
    .PLEQPHASE (PLEQPHASE_out),
    .PMVOUT (PMVOUT_out),
    .SAXISCCTREADY (SAXISCCTREADY_out),
    .SAXISRQTREADY (SAXISRQTREADY_out),
    .SCANOUT (SCANOUT_out),
    .SPAREOUT (SPAREOUT_out),
    .XILUNCONNBOUT (XILUNCONNBOUT_out),
    .XILUNCONNOUT (XILUNCONNOUT_out),
    .CFGCONFIGSPACEENABLE (CFGCONFIGSPACEENABLE_in),
    .CFGDEVID (CFGDEVID_in),
    .CFGDSBUSNUMBER (CFGDSBUSNUMBER_in),
    .CFGDSDEVICENUMBER (CFGDSDEVICENUMBER_in),
    .CFGDSFUNCTIONNUMBER (CFGDSFUNCTIONNUMBER_in),
    .CFGDSN (CFGDSN_in),
    .CFGDSPORTNUMBER (CFGDSPORTNUMBER_in),
    .CFGERRCORIN (CFGERRCORIN_in),
    .CFGERRUNCORIN (CFGERRUNCORIN_in),
    .CFGEXTREADDATA (CFGEXTREADDATA_in),
    .CFGEXTREADDATAVALID (CFGEXTREADDATAVALID_in),
    .CFGFCSEL (CFGFCSEL_in),
    .CFGFLRDONE (CFGFLRDONE_in),
    .CFGHOTRESETIN (CFGHOTRESETIN_in),
    .CFGINTERRUPTINT (CFGINTERRUPTINT_in),
    .CFGINTERRUPTMSIATTR (CFGINTERRUPTMSIATTR_in),
    .CFGINTERRUPTMSIFUNCTIONNUMBER (CFGINTERRUPTMSIFUNCTIONNUMBER_in),
    .CFGINTERRUPTMSIINT (CFGINTERRUPTMSIINT_in),
    .CFGINTERRUPTMSIPENDINGSTATUS (CFGINTERRUPTMSIPENDINGSTATUS_in),
    .CFGINTERRUPTMSIPENDINGSTATUSDATAENABLE (CFGINTERRUPTMSIPENDINGSTATUSDATAENABLE_in),
    .CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM (CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM_in),
    .CFGINTERRUPTMSISELECT (CFGINTERRUPTMSISELECT_in),
    .CFGINTERRUPTMSITPHPRESENT (CFGINTERRUPTMSITPHPRESENT_in),
    .CFGINTERRUPTMSITPHSTTAG (CFGINTERRUPTMSITPHSTTAG_in),
    .CFGINTERRUPTMSITPHTYPE (CFGINTERRUPTMSITPHTYPE_in),
    .CFGINTERRUPTMSIXADDRESS (CFGINTERRUPTMSIXADDRESS_in),
    .CFGINTERRUPTMSIXDATA (CFGINTERRUPTMSIXDATA_in),
    .CFGINTERRUPTMSIXINT (CFGINTERRUPTMSIXINT_in),
    .CFGINTERRUPTPENDING (CFGINTERRUPTPENDING_in),
    .CFGLINKTRAININGENABLE (CFGLINKTRAININGENABLE_in),
    .CFGMGMTADDR (CFGMGMTADDR_in),
    .CFGMGMTBYTEENABLE (CFGMGMTBYTEENABLE_in),
    .CFGMGMTREAD (CFGMGMTREAD_in),
    .CFGMGMTTYPE1CFGREGACCESS (CFGMGMTTYPE1CFGREGACCESS_in),
    .CFGMGMTWRITE (CFGMGMTWRITE_in),
    .CFGMGMTWRITEDATA (CFGMGMTWRITEDATA_in),
    .CFGMSGTRANSMIT (CFGMSGTRANSMIT_in),
    .CFGMSGTRANSMITDATA (CFGMSGTRANSMITDATA_in),
    .CFGMSGTRANSMITTYPE (CFGMSGTRANSMITTYPE_in),
    .CFGPERFUNCSTATUSCONTROL (CFGPERFUNCSTATUSCONTROL_in),
    .CFGPERFUNCTIONNUMBER (CFGPERFUNCTIONNUMBER_in),
    .CFGPERFUNCTIONOUTPUTREQUEST (CFGPERFUNCTIONOUTPUTREQUEST_in),
    .CFGPOWERSTATECHANGEACK (CFGPOWERSTATECHANGEACK_in),
    .CFGREQPMTRANSITIONL23READY (CFGREQPMTRANSITIONL23READY_in),
    .CFGREVID (CFGREVID_in),
    .CFGSUBSYSID (CFGSUBSYSID_in),
    .CFGSUBSYSVENDID (CFGSUBSYSVENDID_in),
    .CFGTPHSTTREADDATA (CFGTPHSTTREADDATA_in),
    .CFGTPHSTTREADDATAVALID (CFGTPHSTTREADDATAVALID_in),
    .CFGVENDID (CFGVENDID_in),
    .CFGVFFLRDONE (CFGVFFLRDONE_in),
    .CONFMCAPREQUESTBYCONF (CONFMCAPREQUESTBYCONF_in),
    .CONFREQDATA (CONFREQDATA_in),
    .CONFREQREGNUM (CONFREQREGNUM_in),
    .CONFREQTYPE (CONFREQTYPE_in),
    .CONFREQVALID (CONFREQVALID_in),
    .CORECLK (CORECLK_in),
    .CORECLKMICOMPLETIONRAML (CORECLKMICOMPLETIONRAML_in),
    .CORECLKMICOMPLETIONRAMU (CORECLKMICOMPLETIONRAMU_in),
    .CORECLKMIREPLAYRAM (CORECLKMIREPLAYRAM_in),
    .CORECLKMIREQUESTRAM (CORECLKMIREQUESTRAM_in),
    .DBGCFGLOCALMGMTREGOVERRIDE (DBGCFGLOCALMGMTREGOVERRIDE_in),
    .DBGDATASEL (DBGDATASEL_in),
    .DRPADDR (DRPADDR_in),
    .DRPCLK (DRPCLK_in),
    .DRPDI (DRPDI_in),
    .DRPEN (DRPEN_in),
    .DRPWE (DRPWE_in),
    .LL2LMSAXISTXTUSER (LL2LMSAXISTXTUSER_in),
    .LL2LMSAXISTXTVALID (LL2LMSAXISTXTVALID_in),
    .LL2LMTXTLPID0 (LL2LMTXTLPID0_in),
    .LL2LMTXTLPID1 (LL2LMTXTLPID1_in),
    .MAXISCQTREADY (MAXISCQTREADY_in),
    .MAXISRCTREADY (MAXISRCTREADY_in),
    .MCAPCLK (MCAPCLK_in),
    .MCAPPERST0B (MCAPPERST0B_in),
    .MCAPPERST1B (MCAPPERST1B_in),
    .MGMTRESETN (MGMTRESETN_in),
    .MGMTSTICKYRESETN (MGMTSTICKYRESETN_in),
    .MICOMPLETIONRAMREADDATA (MICOMPLETIONRAMREADDATA_in),
    .MIREPLAYRAMREADDATA (MIREPLAYRAMREADDATA_in),
    .MIREQUESTRAMREADDATA (MIREQUESTRAMREADDATA_in),
    .PCIECQNPREQ (PCIECQNPREQ_in),
    .PIPECLK (PIPECLK_in),
    .PIPEEQFS (PIPEEQFS_in),
    .PIPEEQLF (PIPEEQLF_in),
    .PIPERESETN (PIPERESETN_in),
    .PIPERX0CHARISK (PIPERX0CHARISK_in),
    .PIPERX0DATA (PIPERX0DATA_in),
    .PIPERX0DATAVALID (PIPERX0DATAVALID_in),
    .PIPERX0ELECIDLE (PIPERX0ELECIDLE_in),
    .PIPERX0EQDONE (PIPERX0EQDONE_in),
    .PIPERX0EQLPADAPTDONE (PIPERX0EQLPADAPTDONE_in),
    .PIPERX0EQLPLFFSSEL (PIPERX0EQLPLFFSSEL_in),
    .PIPERX0EQLPNEWTXCOEFFORPRESET (PIPERX0EQLPNEWTXCOEFFORPRESET_in),
    .PIPERX0PHYSTATUS (PIPERX0PHYSTATUS_in),
    .PIPERX0STARTBLOCK (PIPERX0STARTBLOCK_in),
    .PIPERX0STATUS (PIPERX0STATUS_in),
    .PIPERX0SYNCHEADER (PIPERX0SYNCHEADER_in),
    .PIPERX0VALID (PIPERX0VALID_in),
    .PIPERX1CHARISK (PIPERX1CHARISK_in),
    .PIPERX1DATA (PIPERX1DATA_in),
    .PIPERX1DATAVALID (PIPERX1DATAVALID_in),
    .PIPERX1ELECIDLE (PIPERX1ELECIDLE_in),
    .PIPERX1EQDONE (PIPERX1EQDONE_in),
    .PIPERX1EQLPADAPTDONE (PIPERX1EQLPADAPTDONE_in),
    .PIPERX1EQLPLFFSSEL (PIPERX1EQLPLFFSSEL_in),
    .PIPERX1EQLPNEWTXCOEFFORPRESET (PIPERX1EQLPNEWTXCOEFFORPRESET_in),
    .PIPERX1PHYSTATUS (PIPERX1PHYSTATUS_in),
    .PIPERX1STARTBLOCK (PIPERX1STARTBLOCK_in),
    .PIPERX1STATUS (PIPERX1STATUS_in),
    .PIPERX1SYNCHEADER (PIPERX1SYNCHEADER_in),
    .PIPERX1VALID (PIPERX1VALID_in),
    .PIPERX2CHARISK (PIPERX2CHARISK_in),
    .PIPERX2DATA (PIPERX2DATA_in),
    .PIPERX2DATAVALID (PIPERX2DATAVALID_in),
    .PIPERX2ELECIDLE (PIPERX2ELECIDLE_in),
    .PIPERX2EQDONE (PIPERX2EQDONE_in),
    .PIPERX2EQLPADAPTDONE (PIPERX2EQLPADAPTDONE_in),
    .PIPERX2EQLPLFFSSEL (PIPERX2EQLPLFFSSEL_in),
    .PIPERX2EQLPNEWTXCOEFFORPRESET (PIPERX2EQLPNEWTXCOEFFORPRESET_in),
    .PIPERX2PHYSTATUS (PIPERX2PHYSTATUS_in),
    .PIPERX2STARTBLOCK (PIPERX2STARTBLOCK_in),
    .PIPERX2STATUS (PIPERX2STATUS_in),
    .PIPERX2SYNCHEADER (PIPERX2SYNCHEADER_in),
    .PIPERX2VALID (PIPERX2VALID_in),
    .PIPERX3CHARISK (PIPERX3CHARISK_in),
    .PIPERX3DATA (PIPERX3DATA_in),
    .PIPERX3DATAVALID (PIPERX3DATAVALID_in),
    .PIPERX3ELECIDLE (PIPERX3ELECIDLE_in),
    .PIPERX3EQDONE (PIPERX3EQDONE_in),
    .PIPERX3EQLPADAPTDONE (PIPERX3EQLPADAPTDONE_in),
    .PIPERX3EQLPLFFSSEL (PIPERX3EQLPLFFSSEL_in),
    .PIPERX3EQLPNEWTXCOEFFORPRESET (PIPERX3EQLPNEWTXCOEFFORPRESET_in),
    .PIPERX3PHYSTATUS (PIPERX3PHYSTATUS_in),
    .PIPERX3STARTBLOCK (PIPERX3STARTBLOCK_in),
    .PIPERX3STATUS (PIPERX3STATUS_in),
    .PIPERX3SYNCHEADER (PIPERX3SYNCHEADER_in),
    .PIPERX3VALID (PIPERX3VALID_in),
    .PIPERX4CHARISK (PIPERX4CHARISK_in),
    .PIPERX4DATA (PIPERX4DATA_in),
    .PIPERX4DATAVALID (PIPERX4DATAVALID_in),
    .PIPERX4ELECIDLE (PIPERX4ELECIDLE_in),
    .PIPERX4EQDONE (PIPERX4EQDONE_in),
    .PIPERX4EQLPADAPTDONE (PIPERX4EQLPADAPTDONE_in),
    .PIPERX4EQLPLFFSSEL (PIPERX4EQLPLFFSSEL_in),
    .PIPERX4EQLPNEWTXCOEFFORPRESET (PIPERX4EQLPNEWTXCOEFFORPRESET_in),
    .PIPERX4PHYSTATUS (PIPERX4PHYSTATUS_in),
    .PIPERX4STARTBLOCK (PIPERX4STARTBLOCK_in),
    .PIPERX4STATUS (PIPERX4STATUS_in),
    .PIPERX4SYNCHEADER (PIPERX4SYNCHEADER_in),
    .PIPERX4VALID (PIPERX4VALID_in),
    .PIPERX5CHARISK (PIPERX5CHARISK_in),
    .PIPERX5DATA (PIPERX5DATA_in),
    .PIPERX5DATAVALID (PIPERX5DATAVALID_in),
    .PIPERX5ELECIDLE (PIPERX5ELECIDLE_in),
    .PIPERX5EQDONE (PIPERX5EQDONE_in),
    .PIPERX5EQLPADAPTDONE (PIPERX5EQLPADAPTDONE_in),
    .PIPERX5EQLPLFFSSEL (PIPERX5EQLPLFFSSEL_in),
    .PIPERX5EQLPNEWTXCOEFFORPRESET (PIPERX5EQLPNEWTXCOEFFORPRESET_in),
    .PIPERX5PHYSTATUS (PIPERX5PHYSTATUS_in),
    .PIPERX5STARTBLOCK (PIPERX5STARTBLOCK_in),
    .PIPERX5STATUS (PIPERX5STATUS_in),
    .PIPERX5SYNCHEADER (PIPERX5SYNCHEADER_in),
    .PIPERX5VALID (PIPERX5VALID_in),
    .PIPERX6CHARISK (PIPERX6CHARISK_in),
    .PIPERX6DATA (PIPERX6DATA_in),
    .PIPERX6DATAVALID (PIPERX6DATAVALID_in),
    .PIPERX6ELECIDLE (PIPERX6ELECIDLE_in),
    .PIPERX6EQDONE (PIPERX6EQDONE_in),
    .PIPERX6EQLPADAPTDONE (PIPERX6EQLPADAPTDONE_in),
    .PIPERX6EQLPLFFSSEL (PIPERX6EQLPLFFSSEL_in),
    .PIPERX6EQLPNEWTXCOEFFORPRESET (PIPERX6EQLPNEWTXCOEFFORPRESET_in),
    .PIPERX6PHYSTATUS (PIPERX6PHYSTATUS_in),
    .PIPERX6STARTBLOCK (PIPERX6STARTBLOCK_in),
    .PIPERX6STATUS (PIPERX6STATUS_in),
    .PIPERX6SYNCHEADER (PIPERX6SYNCHEADER_in),
    .PIPERX6VALID (PIPERX6VALID_in),
    .PIPERX7CHARISK (PIPERX7CHARISK_in),
    .PIPERX7DATA (PIPERX7DATA_in),
    .PIPERX7DATAVALID (PIPERX7DATAVALID_in),
    .PIPERX7ELECIDLE (PIPERX7ELECIDLE_in),
    .PIPERX7EQDONE (PIPERX7EQDONE_in),
    .PIPERX7EQLPADAPTDONE (PIPERX7EQLPADAPTDONE_in),
    .PIPERX7EQLPLFFSSEL (PIPERX7EQLPLFFSSEL_in),
    .PIPERX7EQLPNEWTXCOEFFORPRESET (PIPERX7EQLPNEWTXCOEFFORPRESET_in),
    .PIPERX7PHYSTATUS (PIPERX7PHYSTATUS_in),
    .PIPERX7STARTBLOCK (PIPERX7STARTBLOCK_in),
    .PIPERX7STATUS (PIPERX7STATUS_in),
    .PIPERX7SYNCHEADER (PIPERX7SYNCHEADER_in),
    .PIPERX7VALID (PIPERX7VALID_in),
    .PIPETX0EQCOEFF (PIPETX0EQCOEFF_in),
    .PIPETX0EQDONE (PIPETX0EQDONE_in),
    .PIPETX1EQCOEFF (PIPETX1EQCOEFF_in),
    .PIPETX1EQDONE (PIPETX1EQDONE_in),
    .PIPETX2EQCOEFF (PIPETX2EQCOEFF_in),
    .PIPETX2EQDONE (PIPETX2EQDONE_in),
    .PIPETX3EQCOEFF (PIPETX3EQCOEFF_in),
    .PIPETX3EQDONE (PIPETX3EQDONE_in),
    .PIPETX4EQCOEFF (PIPETX4EQCOEFF_in),
    .PIPETX4EQDONE (PIPETX4EQDONE_in),
    .PIPETX5EQCOEFF (PIPETX5EQCOEFF_in),
    .PIPETX5EQDONE (PIPETX5EQDONE_in),
    .PIPETX6EQCOEFF (PIPETX6EQCOEFF_in),
    .PIPETX6EQDONE (PIPETX6EQDONE_in),
    .PIPETX7EQCOEFF (PIPETX7EQCOEFF_in),
    .PIPETX7EQDONE (PIPETX7EQDONE_in),
    .PLEQRESETEIEOSCOUNT (PLEQRESETEIEOSCOUNT_in),
    .PLGEN2UPSTREAMPREFERDEEMPH (PLGEN2UPSTREAMPREFERDEEMPH_in),
    .PMVDIVIDE (PMVDIVIDE_in),
    .PMVENABLEN (PMVENABLEN_in),
    .PMVSELECT (PMVSELECT_in),
    .RESETN (RESETN_in),
    .SAXISCCTDATA (SAXISCCTDATA_in),
    .SAXISCCTKEEP (SAXISCCTKEEP_in),
    .SAXISCCTLAST (SAXISCCTLAST_in),
    .SAXISCCTUSER (SAXISCCTUSER_in),
    .SAXISCCTVALID (SAXISCCTVALID_in),
    .SAXISRQTDATA (SAXISRQTDATA_in),
    .SAXISRQTKEEP (SAXISRQTKEEP_in),
    .SAXISRQTLAST (SAXISRQTLAST_in),
    .SAXISRQTUSER (SAXISRQTUSER_in),
    .SAXISRQTVALID (SAXISRQTVALID_in),
    .SCANENABLEN (SCANENABLEN_in),
    .SCANIN (SCANIN_in),
    .SCANMODEN (SCANMODEN_in),
    .SPAREIN (SPAREIN_in),
    .USERCLK (USERCLK_in),
    .XILUNCONNBYP (XILUNCONNBYP_in),
    .XILUNCONNCLK (XILUNCONNCLK_in),
    .XILUNCONNIN (XILUNCONNIN_in),
    .GSR (glblGSR)
  );

    specify
    (CORECLK => DBGDATAOUT[0]) = (0:0:0, 0:0:0);
    (CORECLK => DBGDATAOUT[10]) = (0:0:0, 0:0:0);
    (CORECLK => DBGDATAOUT[11]) = (0:0:0, 0:0:0);
    (CORECLK => DBGDATAOUT[12]) = (0:0:0, 0:0:0);
    (CORECLK => DBGDATAOUT[13]) = (0:0:0, 0:0:0);
    (CORECLK => DBGDATAOUT[14]) = (0:0:0, 0:0:0);
    (CORECLK => DBGDATAOUT[15]) = (0:0:0, 0:0:0);
    (CORECLK => DBGDATAOUT[1]) = (0:0:0, 0:0:0);
    (CORECLK => DBGDATAOUT[2]) = (0:0:0, 0:0:0);
    (CORECLK => DBGDATAOUT[3]) = (0:0:0, 0:0:0);
    (CORECLK => DBGDATAOUT[4]) = (0:0:0, 0:0:0);
    (CORECLK => DBGDATAOUT[5]) = (0:0:0, 0:0:0);
    (CORECLK => DBGDATAOUT[6]) = (0:0:0, 0:0:0);
    (CORECLK => DBGDATAOUT[7]) = (0:0:0, 0:0:0);
    (CORECLK => DBGDATAOUT[8]) = (0:0:0, 0:0:0);
    (CORECLK => DBGDATAOUT[9]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMREADADDRESSAL[0]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMREADADDRESSAL[1]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMREADADDRESSAL[2]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMREADADDRESSAL[3]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMREADADDRESSAL[4]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMREADADDRESSAL[5]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMREADADDRESSAL[6]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMREADADDRESSAL[7]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMREADADDRESSAL[8]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMREADADDRESSAL[9]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMREADADDRESSBL[0]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMREADADDRESSBL[1]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMREADADDRESSBL[2]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMREADADDRESSBL[3]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMREADADDRESSBL[4]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMREADADDRESSBL[5]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMREADADDRESSBL[6]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMREADADDRESSBL[7]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMREADADDRESSBL[8]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMREADADDRESSBL[9]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMREADENABLEL[0]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMREADENABLEL[1]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMREADENABLEL[2]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMREADENABLEL[3]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEADDRESSAL[0]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEADDRESSAL[1]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEADDRESSAL[2]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEADDRESSAL[3]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEADDRESSAL[4]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEADDRESSAL[5]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEADDRESSAL[6]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEADDRESSAL[7]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEADDRESSAL[8]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEADDRESSAL[9]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEADDRESSBL[0]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEADDRESSBL[1]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEADDRESSBL[2]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEADDRESSBL[3]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEADDRESSBL[4]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEADDRESSBL[5]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEADDRESSBL[6]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEADDRESSBL[7]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEADDRESSBL[8]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEADDRESSBL[9]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[0]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[10]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[11]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[12]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[13]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[14]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[15]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[16]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[17]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[18]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[19]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[1]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[20]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[21]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[22]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[23]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[24]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[25]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[26]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[27]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[28]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[29]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[2]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[30]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[31]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[32]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[33]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[34]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[35]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[36]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[37]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[38]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[39]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[3]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[40]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[41]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[42]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[43]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[44]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[45]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[46]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[47]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[48]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[49]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[4]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[50]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[51]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[52]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[53]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[54]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[55]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[56]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[57]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[58]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[59]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[5]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[60]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[61]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[62]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[63]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[64]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[65]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[66]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[67]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[68]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[69]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[6]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[70]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[71]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[7]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[8]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEDATAL[9]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEENABLEL[0]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEENABLEL[1]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEENABLEL[2]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAML => MICOMPLETIONRAMWRITEENABLEL[3]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMREADADDRESSAU[0]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMREADADDRESSAU[1]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMREADADDRESSAU[2]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMREADADDRESSAU[3]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMREADADDRESSAU[4]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMREADADDRESSAU[5]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMREADADDRESSAU[6]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMREADADDRESSAU[7]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMREADADDRESSAU[8]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMREADADDRESSAU[9]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMREADADDRESSBU[0]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMREADADDRESSBU[1]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMREADADDRESSBU[2]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMREADADDRESSBU[3]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMREADADDRESSBU[4]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMREADADDRESSBU[5]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMREADADDRESSBU[6]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMREADADDRESSBU[7]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMREADADDRESSBU[8]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMREADADDRESSBU[9]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMREADENABLEU[0]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMREADENABLEU[1]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMREADENABLEU[2]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMREADENABLEU[3]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEADDRESSAU[0]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEADDRESSAU[1]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEADDRESSAU[2]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEADDRESSAU[3]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEADDRESSAU[4]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEADDRESSAU[5]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEADDRESSAU[6]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEADDRESSAU[7]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEADDRESSAU[8]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEADDRESSAU[9]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEADDRESSBU[0]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEADDRESSBU[1]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEADDRESSBU[2]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEADDRESSBU[3]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEADDRESSBU[4]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEADDRESSBU[5]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEADDRESSBU[6]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEADDRESSBU[7]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEADDRESSBU[8]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEADDRESSBU[9]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[0]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[10]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[11]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[12]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[13]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[14]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[15]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[16]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[17]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[18]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[19]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[1]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[20]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[21]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[22]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[23]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[24]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[25]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[26]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[27]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[28]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[29]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[2]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[30]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[31]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[32]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[33]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[34]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[35]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[36]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[37]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[38]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[39]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[3]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[40]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[41]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[42]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[43]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[44]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[45]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[46]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[47]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[48]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[49]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[4]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[50]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[51]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[52]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[53]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[54]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[55]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[56]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[57]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[58]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[59]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[5]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[60]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[61]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[62]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[63]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[64]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[65]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[66]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[67]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[68]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[69]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[6]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[70]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[71]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[7]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[8]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEDATAU[9]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEENABLEU[0]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEENABLEU[1]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEENABLEU[2]) = (0:0:0, 0:0:0);
    (CORECLKMICOMPLETIONRAMU => MICOMPLETIONRAMWRITEENABLEU[3]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMADDRESS[0]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMADDRESS[1]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMADDRESS[2]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMADDRESS[3]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMADDRESS[4]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMADDRESS[5]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMADDRESS[6]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMADDRESS[7]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMADDRESS[8]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMREADENABLE[0]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMREADENABLE[1]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[0]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[100]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[101]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[102]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[103]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[104]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[105]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[106]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[107]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[108]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[109]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[10]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[110]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[111]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[112]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[113]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[114]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[115]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[116]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[117]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[118]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[119]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[11]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[120]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[121]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[122]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[123]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[124]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[125]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[126]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[127]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[128]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[129]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[12]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[130]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[131]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[132]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[133]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[134]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[135]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[136]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[137]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[138]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[139]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[13]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[140]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[141]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[142]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[143]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[14]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[15]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[16]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[17]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[18]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[19]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[1]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[20]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[21]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[22]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[23]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[24]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[25]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[26]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[27]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[28]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[29]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[2]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[30]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[31]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[32]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[33]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[34]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[35]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[36]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[37]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[38]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[39]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[3]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[40]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[41]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[42]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[43]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[44]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[45]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[46]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[47]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[48]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[49]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[4]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[50]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[51]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[52]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[53]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[54]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[55]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[56]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[57]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[58]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[59]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[5]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[60]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[61]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[62]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[63]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[64]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[65]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[66]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[67]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[68]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[69]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[6]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[70]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[71]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[72]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[73]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[74]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[75]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[76]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[77]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[78]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[79]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[7]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[80]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[81]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[82]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[83]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[84]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[85]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[86]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[87]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[88]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[89]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[8]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[90]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[91]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[92]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[93]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[94]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[95]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[96]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[97]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[98]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[99]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEDATA[9]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEENABLE[0]) = (0:0:0, 0:0:0);
    (CORECLKMIREPLAYRAM => MIREPLAYRAMWRITEENABLE[1]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMREADADDRESSA[0]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMREADADDRESSA[1]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMREADADDRESSA[2]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMREADADDRESSA[3]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMREADADDRESSA[4]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMREADADDRESSA[5]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMREADADDRESSA[6]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMREADADDRESSA[7]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMREADADDRESSA[8]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMREADADDRESSB[0]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMREADADDRESSB[1]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMREADADDRESSB[2]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMREADADDRESSB[3]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMREADADDRESSB[4]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMREADADDRESSB[5]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMREADADDRESSB[6]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMREADADDRESSB[7]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMREADADDRESSB[8]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMREADENABLE[0]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMREADENABLE[1]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMREADENABLE[2]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMREADENABLE[3]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEADDRESSA[0]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEADDRESSA[1]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEADDRESSA[2]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEADDRESSA[3]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEADDRESSA[4]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEADDRESSA[5]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEADDRESSA[6]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEADDRESSA[7]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEADDRESSA[8]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEADDRESSB[0]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEADDRESSB[1]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEADDRESSB[2]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEADDRESSB[3]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEADDRESSB[4]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEADDRESSB[5]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEADDRESSB[6]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEADDRESSB[7]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEADDRESSB[8]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[0]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[100]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[101]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[102]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[103]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[104]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[105]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[106]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[107]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[108]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[109]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[10]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[110]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[111]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[112]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[113]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[114]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[115]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[116]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[117]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[118]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[119]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[11]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[120]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[121]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[122]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[123]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[124]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[125]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[126]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[127]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[128]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[129]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[12]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[130]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[131]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[132]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[133]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[134]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[135]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[136]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[137]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[138]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[139]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[13]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[140]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[141]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[142]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[143]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[14]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[15]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[16]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[17]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[18]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[19]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[1]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[20]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[21]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[22]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[23]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[24]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[25]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[26]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[27]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[28]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[29]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[2]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[30]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[31]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[32]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[33]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[34]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[35]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[36]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[37]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[38]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[39]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[3]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[40]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[41]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[42]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[43]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[44]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[45]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[46]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[47]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[48]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[49]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[4]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[50]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[51]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[52]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[53]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[54]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[55]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[56]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[57]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[58]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[59]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[5]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[60]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[61]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[62]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[63]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[64]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[65]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[66]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[67]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[68]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[69]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[6]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[70]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[71]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[72]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[73]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[74]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[75]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[76]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[77]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[78]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[79]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[7]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[80]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[81]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[82]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[83]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[84]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[85]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[86]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[87]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[88]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[89]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[8]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[90]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[91]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[92]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[93]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[94]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[95]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[96]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[97]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[98]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[99]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEDATA[9]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEENABLE[0]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEENABLE[1]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEENABLE[2]) = (0:0:0, 0:0:0);
    (CORECLKMIREQUESTRAM => MIREQUESTRAMWRITEENABLE[3]) = (0:0:0, 0:0:0);
    (DRPCLK => DRPDO[0]) = (0:0:0, 0:0:0);
    (DRPCLK => DRPDO[10]) = (0:0:0, 0:0:0);
    (DRPCLK => DRPDO[11]) = (0:0:0, 0:0:0);
    (DRPCLK => DRPDO[12]) = (0:0:0, 0:0:0);
    (DRPCLK => DRPDO[13]) = (0:0:0, 0:0:0);
    (DRPCLK => DRPDO[14]) = (0:0:0, 0:0:0);
    (DRPCLK => DRPDO[15]) = (0:0:0, 0:0:0);
    (DRPCLK => DRPDO[1]) = (0:0:0, 0:0:0);
    (DRPCLK => DRPDO[2]) = (0:0:0, 0:0:0);
    (DRPCLK => DRPDO[3]) = (0:0:0, 0:0:0);
    (DRPCLK => DRPDO[4]) = (0:0:0, 0:0:0);
    (DRPCLK => DRPDO[5]) = (0:0:0, 0:0:0);
    (DRPCLK => DRPDO[6]) = (0:0:0, 0:0:0);
    (DRPCLK => DRPDO[7]) = (0:0:0, 0:0:0);
    (DRPCLK => DRPDO[8]) = (0:0:0, 0:0:0);
    (DRPCLK => DRPDO[9]) = (0:0:0, 0:0:0);
    (DRPCLK => DRPRDY) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPCSB) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[0]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[10]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[11]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[12]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[13]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[14]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[15]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[16]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[17]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[18]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[19]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[1]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[20]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[21]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[22]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[23]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[24]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[25]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[26]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[27]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[28]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[29]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[2]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[30]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[31]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[3]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[4]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[5]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[6]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[7]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[8]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPDATA[9]) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPEOS) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPERROR) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPMODE) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPRDATAVALID) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPRDWRB) = (0:0:0, 0:0:0);
    (MCAPCLK => DBGMCAPRESET) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX0EQCONTROL[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX0EQCONTROL[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX0EQLPLFFS[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX0EQLPLFFS[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX0EQLPLFFS[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX0EQLPLFFS[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX0EQLPLFFS[4]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX0EQLPLFFS[5]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX0EQLPTXPRESET[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX0EQLPTXPRESET[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX0EQLPTXPRESET[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX0EQLPTXPRESET[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX0EQPRESET[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX0EQPRESET[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX0EQPRESET[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX0POLARITY) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX1EQCONTROL[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX1EQCONTROL[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX1EQLPLFFS[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX1EQLPLFFS[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX1EQLPLFFS[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX1EQLPLFFS[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX1EQLPLFFS[4]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX1EQLPLFFS[5]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX1EQLPTXPRESET[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX1EQLPTXPRESET[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX1EQLPTXPRESET[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX1EQLPTXPRESET[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX1EQPRESET[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX1EQPRESET[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX1EQPRESET[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX1POLARITY) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX2EQCONTROL[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX2EQCONTROL[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX2EQLPLFFS[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX2EQLPLFFS[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX2EQLPLFFS[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX2EQLPLFFS[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX2EQLPLFFS[4]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX2EQLPLFFS[5]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX2EQLPTXPRESET[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX2EQLPTXPRESET[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX2EQLPTXPRESET[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX2EQLPTXPRESET[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX2EQPRESET[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX2EQPRESET[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX2EQPRESET[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX2POLARITY) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX3EQCONTROL[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX3EQCONTROL[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX3EQLPLFFS[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX3EQLPLFFS[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX3EQLPLFFS[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX3EQLPLFFS[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX3EQLPLFFS[4]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX3EQLPLFFS[5]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX3EQLPTXPRESET[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX3EQLPTXPRESET[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX3EQLPTXPRESET[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX3EQLPTXPRESET[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX3EQPRESET[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX3EQPRESET[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX3EQPRESET[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX3POLARITY) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX4EQCONTROL[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX4EQCONTROL[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX4EQLPLFFS[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX4EQLPLFFS[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX4EQLPLFFS[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX4EQLPLFFS[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX4EQLPLFFS[4]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX4EQLPLFFS[5]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX4EQLPTXPRESET[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX4EQLPTXPRESET[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX4EQLPTXPRESET[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX4EQLPTXPRESET[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX4EQPRESET[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX4EQPRESET[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX4EQPRESET[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX4POLARITY) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX5EQCONTROL[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX5EQCONTROL[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX5EQLPLFFS[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX5EQLPLFFS[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX5EQLPLFFS[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX5EQLPLFFS[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX5EQLPLFFS[4]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX5EQLPLFFS[5]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX5EQLPTXPRESET[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX5EQLPTXPRESET[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX5EQLPTXPRESET[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX5EQLPTXPRESET[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX5EQPRESET[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX5EQPRESET[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX5EQPRESET[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX5POLARITY) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX6EQCONTROL[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX6EQCONTROL[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX6EQLPLFFS[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX6EQLPLFFS[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX6EQLPLFFS[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX6EQLPLFFS[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX6EQLPLFFS[4]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX6EQLPLFFS[5]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX6EQLPTXPRESET[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX6EQLPTXPRESET[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX6EQLPTXPRESET[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX6EQLPTXPRESET[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX6EQPRESET[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX6EQPRESET[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX6EQPRESET[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX6POLARITY) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX7EQCONTROL[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX7EQCONTROL[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX7EQLPLFFS[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX7EQLPLFFS[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX7EQLPLFFS[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX7EQLPLFFS[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX7EQLPLFFS[4]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX7EQLPLFFS[5]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX7EQLPTXPRESET[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX7EQLPTXPRESET[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX7EQLPTXPRESET[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX7EQLPTXPRESET[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX7EQPRESET[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX7EQPRESET[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX7EQPRESET[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPERX7POLARITY) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0CHARISK[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0CHARISK[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0COMPLIANCE) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATAVALID) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[10]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[11]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[12]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[13]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[14]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[15]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[16]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[17]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[18]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[19]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[20]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[21]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[22]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[23]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[24]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[25]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[26]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[27]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[28]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[29]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[30]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[31]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[4]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[5]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[6]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[7]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[8]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DATA[9]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0DEEMPH) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0ELECIDLE) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0EQCONTROL[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0EQCONTROL[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0EQDEEMPH[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0EQDEEMPH[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0EQDEEMPH[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0EQDEEMPH[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0EQDEEMPH[4]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0EQDEEMPH[5]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0EQPRESET[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0EQPRESET[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0EQPRESET[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0EQPRESET[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0MARGIN[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0MARGIN[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0MARGIN[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0POWERDOWN[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0POWERDOWN[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0RATE[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0RATE[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0RCVRDET) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0RESET) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0STARTBLOCK) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0SWING) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0SYNCHEADER[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX0SYNCHEADER[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1CHARISK[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1CHARISK[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1COMPLIANCE) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATAVALID) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[10]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[11]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[12]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[13]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[14]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[15]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[16]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[17]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[18]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[19]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[20]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[21]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[22]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[23]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[24]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[25]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[26]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[27]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[28]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[29]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[30]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[31]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[4]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[5]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[6]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[7]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[8]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DATA[9]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1DEEMPH) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1ELECIDLE) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1EQCONTROL[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1EQCONTROL[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1EQDEEMPH[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1EQDEEMPH[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1EQDEEMPH[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1EQDEEMPH[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1EQDEEMPH[4]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1EQDEEMPH[5]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1EQPRESET[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1EQPRESET[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1EQPRESET[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1EQPRESET[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1MARGIN[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1MARGIN[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1MARGIN[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1POWERDOWN[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1POWERDOWN[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1RATE[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1RATE[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1RCVRDET) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1RESET) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1STARTBLOCK) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1SWING) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1SYNCHEADER[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX1SYNCHEADER[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2CHARISK[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2CHARISK[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2COMPLIANCE) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATAVALID) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[10]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[11]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[12]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[13]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[14]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[15]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[16]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[17]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[18]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[19]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[20]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[21]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[22]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[23]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[24]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[25]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[26]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[27]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[28]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[29]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[30]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[31]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[4]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[5]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[6]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[7]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[8]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DATA[9]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2DEEMPH) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2ELECIDLE) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2EQCONTROL[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2EQCONTROL[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2EQDEEMPH[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2EQDEEMPH[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2EQDEEMPH[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2EQDEEMPH[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2EQDEEMPH[4]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2EQDEEMPH[5]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2EQPRESET[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2EQPRESET[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2EQPRESET[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2EQPRESET[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2MARGIN[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2MARGIN[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2MARGIN[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2POWERDOWN[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2POWERDOWN[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2RATE[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2RATE[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2RCVRDET) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2RESET) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2STARTBLOCK) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2SWING) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2SYNCHEADER[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX2SYNCHEADER[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3CHARISK[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3CHARISK[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3COMPLIANCE) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATAVALID) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[10]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[11]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[12]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[13]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[14]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[15]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[16]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[17]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[18]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[19]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[20]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[21]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[22]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[23]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[24]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[25]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[26]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[27]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[28]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[29]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[30]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[31]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[4]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[5]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[6]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[7]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[8]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DATA[9]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3DEEMPH) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3ELECIDLE) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3EQCONTROL[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3EQCONTROL[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3EQDEEMPH[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3EQDEEMPH[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3EQDEEMPH[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3EQDEEMPH[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3EQDEEMPH[4]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3EQDEEMPH[5]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3EQPRESET[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3EQPRESET[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3EQPRESET[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3EQPRESET[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3MARGIN[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3MARGIN[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3MARGIN[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3POWERDOWN[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3POWERDOWN[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3RATE[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3RATE[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3RCVRDET) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3RESET) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3STARTBLOCK) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3SWING) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3SYNCHEADER[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX3SYNCHEADER[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4CHARISK[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4CHARISK[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4COMPLIANCE) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATAVALID) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[10]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[11]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[12]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[13]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[14]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[15]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[16]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[17]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[18]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[19]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[20]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[21]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[22]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[23]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[24]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[25]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[26]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[27]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[28]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[29]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[30]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[31]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[4]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[5]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[6]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[7]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[8]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DATA[9]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4DEEMPH) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4ELECIDLE) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4EQCONTROL[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4EQCONTROL[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4EQDEEMPH[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4EQDEEMPH[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4EQDEEMPH[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4EQDEEMPH[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4EQDEEMPH[4]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4EQDEEMPH[5]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4EQPRESET[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4EQPRESET[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4EQPRESET[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4EQPRESET[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4MARGIN[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4MARGIN[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4MARGIN[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4POWERDOWN[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4POWERDOWN[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4RATE[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4RATE[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4RCVRDET) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4RESET) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4STARTBLOCK) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4SWING) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4SYNCHEADER[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX4SYNCHEADER[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5CHARISK[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5CHARISK[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5COMPLIANCE) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATAVALID) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[10]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[11]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[12]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[13]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[14]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[15]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[16]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[17]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[18]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[19]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[20]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[21]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[22]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[23]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[24]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[25]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[26]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[27]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[28]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[29]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[30]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[31]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[4]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[5]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[6]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[7]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[8]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DATA[9]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5DEEMPH) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5ELECIDLE) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5EQCONTROL[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5EQCONTROL[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5EQDEEMPH[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5EQDEEMPH[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5EQDEEMPH[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5EQDEEMPH[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5EQDEEMPH[4]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5EQDEEMPH[5]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5EQPRESET[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5EQPRESET[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5EQPRESET[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5EQPRESET[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5MARGIN[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5MARGIN[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5MARGIN[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5POWERDOWN[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5POWERDOWN[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5RATE[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5RATE[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5RCVRDET) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5RESET) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5STARTBLOCK) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5SWING) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5SYNCHEADER[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX5SYNCHEADER[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6CHARISK[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6CHARISK[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6COMPLIANCE) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATAVALID) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[10]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[11]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[12]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[13]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[14]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[15]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[16]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[17]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[18]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[19]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[20]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[21]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[22]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[23]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[24]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[25]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[26]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[27]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[28]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[29]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[30]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[31]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[4]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[5]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[6]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[7]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[8]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DATA[9]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6DEEMPH) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6ELECIDLE) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6EQCONTROL[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6EQCONTROL[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6EQDEEMPH[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6EQDEEMPH[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6EQDEEMPH[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6EQDEEMPH[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6EQDEEMPH[4]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6EQDEEMPH[5]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6EQPRESET[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6EQPRESET[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6EQPRESET[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6EQPRESET[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6MARGIN[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6MARGIN[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6MARGIN[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6POWERDOWN[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6POWERDOWN[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6RATE[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6RATE[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6RCVRDET) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6RESET) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6STARTBLOCK) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6SWING) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6SYNCHEADER[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX6SYNCHEADER[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7CHARISK[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7CHARISK[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7COMPLIANCE) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATAVALID) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[10]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[11]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[12]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[13]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[14]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[15]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[16]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[17]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[18]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[19]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[20]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[21]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[22]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[23]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[24]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[25]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[26]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[27]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[28]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[29]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[30]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[31]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[4]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[5]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[6]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[7]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[8]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DATA[9]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7DEEMPH) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7ELECIDLE) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7EQCONTROL[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7EQCONTROL[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7EQDEEMPH[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7EQDEEMPH[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7EQDEEMPH[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7EQDEEMPH[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7EQDEEMPH[4]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7EQDEEMPH[5]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7EQPRESET[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7EQPRESET[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7EQPRESET[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7EQPRESET[3]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7MARGIN[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7MARGIN[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7MARGIN[2]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7POWERDOWN[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7POWERDOWN[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7RATE[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7RATE[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7RCVRDET) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7RESET) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7STARTBLOCK) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7SWING) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7SYNCHEADER[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PIPETX7SYNCHEADER[1]) = (0:0:0, 0:0:0);
    (PIPECLK => PLEQINPROGRESS) = (0:0:0, 0:0:0);
    (PIPECLK => PLEQPHASE[0]) = (0:0:0, 0:0:0);
    (PIPECLK => PLEQPHASE[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGCURRENTSPEED[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGCURRENTSPEED[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGCURRENTSPEED[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGDPASUBSTATECHANGE[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGDPASUBSTATECHANGE[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGERRCOROUT) = (0:0:0, 0:0:0);
    (USERCLK => CFGERRFATALOUT) = (0:0:0, 0:0:0);
    (USERCLK => CFGERRNONFATALOUT) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTFUNCTIONNUMBER[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTFUNCTIONNUMBER[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTFUNCTIONNUMBER[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTFUNCTIONNUMBER[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTFUNCTIONNUMBER[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTFUNCTIONNUMBER[5]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTFUNCTIONNUMBER[6]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTFUNCTIONNUMBER[7]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTREADRECEIVED) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTREGISTERNUMBER[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTREGISTERNUMBER[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTREGISTERNUMBER[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTREGISTERNUMBER[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTREGISTERNUMBER[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTREGISTERNUMBER[5]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTREGISTERNUMBER[6]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTREGISTERNUMBER[7]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTREGISTERNUMBER[8]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTREGISTERNUMBER[9]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEBYTEENABLE[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEBYTEENABLE[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEBYTEENABLE[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEBYTEENABLE[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[10]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[11]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[12]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[13]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[14]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[15]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[16]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[17]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[18]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[19]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[20]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[21]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[22]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[23]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[24]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[25]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[26]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[27]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[28]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[29]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[30]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[31]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[5]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[6]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[7]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[8]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITEDATA[9]) = (0:0:0, 0:0:0);
    (USERCLK => CFGEXTWRITERECEIVED) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCCPLD[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCCPLD[10]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCCPLD[11]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCCPLD[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCCPLD[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCCPLD[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCCPLD[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCCPLD[5]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCCPLD[6]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCCPLD[7]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCCPLD[8]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCCPLD[9]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCCPLH[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCCPLH[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCCPLH[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCCPLH[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCCPLH[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCCPLH[5]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCCPLH[6]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCCPLH[7]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCNPD[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCNPD[10]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCNPD[11]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCNPD[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCNPD[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCNPD[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCNPD[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCNPD[5]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCNPD[6]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCNPD[7]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCNPD[8]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCNPD[9]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCNPH[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCNPH[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCNPH[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCNPH[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCNPH[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCNPH[5]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCNPH[6]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCNPH[7]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCPD[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCPD[10]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCPD[11]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCPD[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCPD[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCPD[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCPD[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCPD[5]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCPD[6]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCPD[7]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCPD[8]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCPD[9]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCPH[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCPH[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCPH[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCPH[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCPH[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCPH[5]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCPH[6]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFCPH[7]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFLRINPROCESS[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFLRINPROCESS[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFUNCTIONPOWERSTATE[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFUNCTIONPOWERSTATE[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFUNCTIONPOWERSTATE[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFUNCTIONPOWERSTATE[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFUNCTIONPOWERSTATE[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFUNCTIONPOWERSTATE[5]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFUNCTIONSTATUS[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFUNCTIONSTATUS[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFUNCTIONSTATUS[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFUNCTIONSTATUS[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFUNCTIONSTATUS[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFUNCTIONSTATUS[5]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFUNCTIONSTATUS[6]) = (0:0:0, 0:0:0);
    (USERCLK => CFGFUNCTIONSTATUS[7]) = (0:0:0, 0:0:0);
    (USERCLK => CFGHOTRESETOUT) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[10]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[11]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[12]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[13]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[14]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[15]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[16]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[17]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[18]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[19]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[20]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[21]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[22]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[23]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[24]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[25]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[26]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[27]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[28]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[29]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[30]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[31]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[5]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[6]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[7]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[8]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIDATA[9]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIENABLE[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIENABLE[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIFAIL) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIMASKUPDATE) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIMMENABLE[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIMMENABLE[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIMMENABLE[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIMMENABLE[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIMMENABLE[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIMMENABLE[5]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSISENT) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIVFENABLE[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIVFENABLE[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIVFENABLE[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIVFENABLE[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIVFENABLE[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIVFENABLE[5]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIXENABLE[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIXENABLE[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIXFAIL) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIXMASK[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIXMASK[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIXSENT) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIXVFENABLE[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIXVFENABLE[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIXVFENABLE[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIXVFENABLE[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIXVFENABLE[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIXVFENABLE[5]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIXVFMASK[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIXVFMASK[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIXVFMASK[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIXVFMASK[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIXVFMASK[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTMSIXVFMASK[5]) = (0:0:0, 0:0:0);
    (USERCLK => CFGINTERRUPTSENT) = (0:0:0, 0:0:0);
    (USERCLK => CFGLINKPOWERSTATE[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGLINKPOWERSTATE[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGLOCALERROR) = (0:0:0, 0:0:0);
    (USERCLK => CFGLTRENABLE) = (0:0:0, 0:0:0);
    (USERCLK => CFGLTSSMSTATE[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGLTSSMSTATE[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGLTSSMSTATE[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGLTSSMSTATE[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGLTSSMSTATE[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGLTSSMSTATE[5]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMAXPAYLOAD[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMAXPAYLOAD[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMAXPAYLOAD[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMAXREADREQ[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMAXREADREQ[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMAXREADREQ[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[10]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[11]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[12]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[13]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[14]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[15]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[16]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[17]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[18]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[19]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[20]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[21]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[22]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[23]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[24]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[25]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[26]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[27]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[28]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[29]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[30]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[31]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[5]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[6]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[7]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[8]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADDATA[9]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMGMTREADWRITEDONE) = (0:0:0, 0:0:0);
    (USERCLK => CFGMSGRECEIVED) = (0:0:0, 0:0:0);
    (USERCLK => CFGMSGRECEIVEDDATA[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMSGRECEIVEDDATA[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMSGRECEIVEDDATA[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMSGRECEIVEDDATA[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMSGRECEIVEDDATA[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMSGRECEIVEDDATA[5]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMSGRECEIVEDDATA[6]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMSGRECEIVEDDATA[7]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMSGRECEIVEDTYPE[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMSGRECEIVEDTYPE[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMSGRECEIVEDTYPE[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMSGRECEIVEDTYPE[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMSGRECEIVEDTYPE[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGMSGTRANSMITDONE) = (0:0:0, 0:0:0);
    (USERCLK => CFGNEGOTIATEDWIDTH[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGNEGOTIATEDWIDTH[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGNEGOTIATEDWIDTH[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGNEGOTIATEDWIDTH[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGOBFFENABLE[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGOBFFENABLE[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGPERFUNCSTATUSDATA[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGPERFUNCSTATUSDATA[10]) = (0:0:0, 0:0:0);
    (USERCLK => CFGPERFUNCSTATUSDATA[11]) = (0:0:0, 0:0:0);
    (USERCLK => CFGPERFUNCSTATUSDATA[12]) = (0:0:0, 0:0:0);
    (USERCLK => CFGPERFUNCSTATUSDATA[13]) = (0:0:0, 0:0:0);
    (USERCLK => CFGPERFUNCSTATUSDATA[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGPERFUNCSTATUSDATA[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGPERFUNCSTATUSDATA[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGPERFUNCSTATUSDATA[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGPERFUNCSTATUSDATA[5]) = (0:0:0, 0:0:0);
    (USERCLK => CFGPERFUNCSTATUSDATA[6]) = (0:0:0, 0:0:0);
    (USERCLK => CFGPERFUNCSTATUSDATA[7]) = (0:0:0, 0:0:0);
    (USERCLK => CFGPERFUNCSTATUSDATA[8]) = (0:0:0, 0:0:0);
    (USERCLK => CFGPERFUNCSTATUSDATA[9]) = (0:0:0, 0:0:0);
    (USERCLK => CFGPERFUNCTIONUPDATEDONE) = (0:0:0, 0:0:0);
    (USERCLK => CFGPHYLINKDOWN) = (0:0:0, 0:0:0);
    (USERCLK => CFGPHYLINKSTATUS[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGPHYLINKSTATUS[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGPLSTATUSCHANGE) = (0:0:0, 0:0:0);
    (USERCLK => CFGPOWERSTATECHANGEINTERRUPT) = (0:0:0, 0:0:0);
    (USERCLK => CFGRCBSTATUS[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGRCBSTATUS[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHFUNCTIONNUM[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHFUNCTIONNUM[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHFUNCTIONNUM[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHFUNCTIONNUM[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHREQUESTERENABLE[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHREQUESTERENABLE[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTMODE[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTMODE[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTMODE[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTMODE[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTMODE[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTMODE[5]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTADDRESS[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTADDRESS[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTADDRESS[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTADDRESS[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTADDRESS[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTREADENABLE) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEBYTEVALID[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEBYTEVALID[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEBYTEVALID[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEBYTEVALID[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[10]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[11]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[12]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[13]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[14]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[15]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[16]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[17]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[18]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[19]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[20]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[21]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[22]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[23]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[24]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[25]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[26]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[27]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[28]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[29]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[30]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[31]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[5]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[6]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[7]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[8]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEDATA[9]) = (0:0:0, 0:0:0);
    (USERCLK => CFGTPHSTTWRITEENABLE) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFFLRINPROCESS[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFFLRINPROCESS[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFFLRINPROCESS[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFFLRINPROCESS[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFFLRINPROCESS[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFFLRINPROCESS[5]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFPOWERSTATE[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFPOWERSTATE[10]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFPOWERSTATE[11]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFPOWERSTATE[12]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFPOWERSTATE[13]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFPOWERSTATE[14]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFPOWERSTATE[15]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFPOWERSTATE[16]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFPOWERSTATE[17]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFPOWERSTATE[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFPOWERSTATE[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFPOWERSTATE[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFPOWERSTATE[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFPOWERSTATE[5]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFPOWERSTATE[6]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFPOWERSTATE[7]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFPOWERSTATE[8]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFPOWERSTATE[9]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFSTATUS[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFSTATUS[10]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFSTATUS[11]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFSTATUS[12]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFSTATUS[14]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFSTATUS[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFSTATUS[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFSTATUS[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFSTATUS[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFSTATUS[5]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFSTATUS[6]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFSTATUS[7]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFSTATUS[8]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFSTATUS[9]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFTPHREQUESTERENABLE[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFTPHREQUESTERENABLE[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFTPHREQUESTERENABLE[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFTPHREQUESTERENABLE[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFTPHREQUESTERENABLE[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFTPHREQUESTERENABLE[5]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFTPHSTMODE[0]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFTPHSTMODE[10]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFTPHSTMODE[11]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFTPHSTMODE[12]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFTPHSTMODE[13]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFTPHSTMODE[14]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFTPHSTMODE[15]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFTPHSTMODE[16]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFTPHSTMODE[17]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFTPHSTMODE[1]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFTPHSTMODE[2]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFTPHSTMODE[3]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFTPHSTMODE[4]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFTPHSTMODE[5]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFTPHSTMODE[6]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFTPHSTMODE[7]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFTPHSTMODE[8]) = (0:0:0, 0:0:0);
    (USERCLK => CFGVFTPHSTMODE[9]) = (0:0:0, 0:0:0);
    (USERCLK => CONFMCAPDESIGNSWITCH) = (0:0:0, 0:0:0);
    (USERCLK => CONFMCAPEOS) = (0:0:0, 0:0:0);
    (USERCLK => CONFMCAPINUSEBYPCIE) = (0:0:0, 0:0:0);
    (USERCLK => CONFREQREADY) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[0]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[10]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[11]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[12]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[13]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[14]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[15]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[16]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[17]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[18]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[19]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[1]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[20]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[21]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[22]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[23]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[24]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[25]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[26]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[27]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[28]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[29]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[2]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[30]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[31]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[3]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[4]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[5]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[6]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[7]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[8]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPRDATA[9]) = (0:0:0, 0:0:0);
    (USERCLK => CONFRESPVALID) = (0:0:0, 0:0:0);
    (USERCLK => DBGPLDATABLOCKRECEIVEDAFTEREDS) = (0:0:0, 0:0:0);
    (USERCLK => DBGPLGEN3FRAMINGERRORDETECTED) = (0:0:0, 0:0:0);
    (USERCLK => DBGPLGEN3SYNCHEADERERRORDETECTED) = (0:0:0, 0:0:0);
    (USERCLK => DBGPLINFERREDRXELECTRICALIDLE[0]) = (0:0:0, 0:0:0);
    (USERCLK => DBGPLINFERREDRXELECTRICALIDLE[1]) = (0:0:0, 0:0:0);
    (USERCLK => DBGPLINFERREDRXELECTRICALIDLE[2]) = (0:0:0, 0:0:0);
    (USERCLK => DBGPLINFERREDRXELECTRICALIDLE[3]) = (0:0:0, 0:0:0);
    (USERCLK => DBGPLINFERREDRXELECTRICALIDLE[4]) = (0:0:0, 0:0:0);
    (USERCLK => DBGPLINFERREDRXELECTRICALIDLE[5]) = (0:0:0, 0:0:0);
    (USERCLK => DBGPLINFERREDRXELECTRICALIDLE[6]) = (0:0:0, 0:0:0);
    (USERCLK => DBGPLINFERREDRXELECTRICALIDLE[7]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMASTERTLPSENT0) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMASTERTLPSENT1) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMASTERTLPSENTTLPID0[0]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMASTERTLPSENTTLPID0[1]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMASTERTLPSENTTLPID0[2]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMASTERTLPSENTTLPID0[3]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMASTERTLPSENTTLPID1[0]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMASTERTLPSENTTLPID1[1]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMASTERTLPSENTTLPID1[2]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMASTERTLPSENTTLPID1[3]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[0]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[100]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[101]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[102]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[103]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[104]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[105]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[106]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[107]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[108]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[109]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[10]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[110]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[111]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[112]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[113]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[114]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[115]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[116]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[117]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[118]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[119]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[11]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[120]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[121]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[122]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[123]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[124]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[125]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[126]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[127]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[128]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[129]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[12]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[130]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[131]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[132]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[133]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[134]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[135]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[136]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[137]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[138]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[139]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[13]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[140]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[141]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[142]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[143]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[144]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[145]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[146]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[147]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[148]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[149]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[14]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[150]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[151]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[152]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[153]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[154]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[155]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[156]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[157]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[158]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[159]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[15]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[160]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[161]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[162]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[163]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[164]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[165]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[166]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[167]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[168]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[169]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[16]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[170]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[171]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[172]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[173]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[174]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[175]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[176]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[177]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[178]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[179]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[17]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[180]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[181]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[182]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[183]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[184]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[185]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[186]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[187]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[188]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[189]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[18]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[190]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[191]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[192]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[193]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[194]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[195]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[196]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[197]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[198]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[199]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[19]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[1]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[200]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[201]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[202]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[203]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[204]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[205]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[206]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[207]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[208]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[209]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[20]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[210]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[211]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[212]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[213]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[214]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[215]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[216]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[217]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[218]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[219]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[21]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[220]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[221]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[222]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[223]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[224]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[225]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[226]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[227]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[228]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[229]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[22]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[230]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[231]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[232]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[233]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[234]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[235]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[236]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[237]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[238]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[239]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[23]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[240]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[241]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[242]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[243]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[244]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[245]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[246]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[247]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[248]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[249]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[24]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[250]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[251]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[252]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[253]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[254]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[255]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[25]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[26]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[27]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[28]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[29]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[2]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[30]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[31]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[32]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[33]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[34]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[35]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[36]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[37]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[38]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[39]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[3]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[40]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[41]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[42]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[43]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[44]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[45]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[46]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[47]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[48]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[49]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[4]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[50]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[51]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[52]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[53]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[54]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[55]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[56]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[57]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[58]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[59]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[5]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[60]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[61]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[62]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[63]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[64]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[65]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[66]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[67]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[68]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[69]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[6]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[70]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[71]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[72]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[73]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[74]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[75]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[76]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[77]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[78]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[79]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[7]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[80]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[81]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[82]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[83]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[84]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[85]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[86]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[87]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[88]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[89]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[8]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[90]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[91]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[92]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[93]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[94]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[95]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[96]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[97]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[98]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[99]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTDATA[9]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTUSER[0]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTUSER[10]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTUSER[11]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTUSER[12]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTUSER[13]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTUSER[14]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTUSER[15]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTUSER[16]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTUSER[17]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTUSER[2]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTUSER[3]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTUSER[4]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTUSER[5]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTUSER[6]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTUSER[7]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTUSER[8]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTVALID[0]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTVALID[1]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTVALID[2]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTVALID[3]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTVALID[4]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTVALID[5]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTVALID[6]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMMAXISRXTVALID[7]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMSAXISTXTREADY[0]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMSAXISTXTREADY[1]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMSAXISTXTREADY[2]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMSAXISTXTREADY[3]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMSAXISTXTREADY[4]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMSAXISTXTREADY[5]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMSAXISTXTREADY[6]) = (0:0:0, 0:0:0);
    (USERCLK => LL2LMSAXISTXTREADY[7]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[0]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[100]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[101]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[102]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[103]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[104]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[105]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[106]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[107]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[108]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[109]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[10]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[110]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[111]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[112]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[113]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[114]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[115]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[116]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[117]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[118]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[119]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[11]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[120]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[121]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[122]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[123]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[124]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[125]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[126]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[127]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[128]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[129]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[12]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[130]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[131]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[132]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[133]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[134]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[135]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[136]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[137]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[138]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[139]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[13]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[140]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[141]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[142]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[143]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[144]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[145]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[146]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[147]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[148]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[149]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[14]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[150]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[151]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[152]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[153]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[154]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[155]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[156]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[157]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[158]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[159]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[15]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[160]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[161]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[162]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[163]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[164]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[165]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[166]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[167]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[168]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[169]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[16]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[170]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[171]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[172]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[173]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[174]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[175]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[176]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[177]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[178]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[179]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[17]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[180]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[181]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[182]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[183]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[184]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[185]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[186]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[187]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[188]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[189]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[18]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[190]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[191]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[192]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[193]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[194]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[195]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[196]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[197]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[198]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[199]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[19]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[1]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[200]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[201]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[202]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[203]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[204]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[205]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[206]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[207]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[208]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[209]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[20]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[210]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[211]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[212]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[213]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[214]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[215]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[216]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[217]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[218]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[219]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[21]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[220]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[221]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[222]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[223]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[224]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[225]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[226]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[227]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[228]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[229]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[22]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[230]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[231]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[232]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[233]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[234]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[235]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[236]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[237]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[238]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[239]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[23]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[240]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[241]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[242]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[243]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[244]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[245]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[246]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[247]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[248]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[249]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[24]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[250]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[251]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[252]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[253]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[254]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[255]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[25]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[26]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[27]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[28]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[29]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[2]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[30]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[31]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[32]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[33]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[34]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[35]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[36]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[37]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[38]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[39]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[3]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[40]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[41]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[42]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[43]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[44]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[45]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[46]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[47]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[48]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[49]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[4]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[50]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[51]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[52]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[53]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[54]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[55]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[56]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[57]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[58]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[59]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[5]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[60]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[61]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[62]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[63]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[64]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[65]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[66]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[67]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[68]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[69]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[6]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[70]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[71]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[72]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[73]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[74]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[75]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[76]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[77]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[78]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[79]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[7]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[80]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[81]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[82]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[83]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[84]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[85]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[86]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[87]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[88]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[89]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[8]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[90]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[91]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[92]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[93]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[94]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[95]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[96]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[97]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[98]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[99]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTDATA[9]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTKEEP[0]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTKEEP[1]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTKEEP[2]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTKEEP[3]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTKEEP[4]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTKEEP[5]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTKEEP[6]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTKEEP[7]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTLAST) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[0]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[10]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[11]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[12]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[13]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[14]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[15]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[16]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[17]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[18]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[19]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[1]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[20]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[21]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[22]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[23]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[24]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[25]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[26]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[27]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[28]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[29]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[2]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[30]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[31]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[32]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[33]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[34]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[35]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[36]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[37]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[38]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[39]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[3]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[40]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[41]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[42]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[43]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[44]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[45]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[46]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[47]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[48]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[49]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[4]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[50]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[51]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[52]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[53]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[54]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[55]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[56]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[57]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[58]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[59]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[5]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[60]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[61]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[62]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[63]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[64]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[65]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[66]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[67]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[68]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[69]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[6]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[70]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[71]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[72]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[73]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[74]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[75]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[76]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[77]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[78]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[79]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[7]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[80]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[81]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[82]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[83]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[84]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[8]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTUSER[9]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISCQTVALID) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[0]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[100]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[101]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[102]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[103]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[104]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[105]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[106]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[107]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[108]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[109]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[10]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[110]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[111]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[112]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[113]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[114]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[115]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[116]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[117]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[118]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[119]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[11]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[120]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[121]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[122]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[123]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[124]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[125]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[126]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[127]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[128]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[129]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[12]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[130]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[131]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[132]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[133]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[134]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[135]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[136]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[137]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[138]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[139]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[13]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[140]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[141]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[142]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[143]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[144]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[145]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[146]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[147]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[148]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[149]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[14]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[150]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[151]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[152]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[153]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[154]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[155]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[156]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[157]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[158]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[159]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[15]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[160]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[161]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[162]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[163]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[164]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[165]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[166]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[167]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[168]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[169]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[16]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[170]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[171]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[172]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[173]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[174]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[175]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[176]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[177]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[178]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[179]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[17]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[180]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[181]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[182]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[183]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[184]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[185]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[186]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[187]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[188]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[189]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[18]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[190]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[191]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[192]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[193]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[194]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[195]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[196]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[197]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[198]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[199]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[19]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[1]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[200]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[201]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[202]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[203]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[204]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[205]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[206]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[207]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[208]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[209]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[20]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[210]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[211]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[212]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[213]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[214]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[215]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[216]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[217]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[218]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[219]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[21]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[220]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[221]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[222]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[223]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[224]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[225]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[226]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[227]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[228]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[229]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[22]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[230]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[231]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[232]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[233]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[234]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[235]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[236]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[237]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[238]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[239]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[23]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[240]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[241]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[242]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[243]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[244]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[245]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[246]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[247]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[248]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[249]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[24]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[250]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[251]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[252]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[253]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[254]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[255]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[25]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[26]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[27]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[28]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[29]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[2]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[30]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[31]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[32]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[33]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[34]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[35]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[36]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[37]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[38]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[39]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[3]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[40]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[41]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[42]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[43]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[44]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[45]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[46]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[47]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[48]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[49]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[4]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[50]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[51]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[52]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[53]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[54]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[55]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[56]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[57]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[58]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[59]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[5]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[60]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[61]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[62]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[63]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[64]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[65]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[66]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[67]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[68]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[69]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[6]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[70]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[71]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[72]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[73]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[74]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[75]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[76]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[77]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[78]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[79]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[7]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[80]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[81]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[82]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[83]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[84]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[85]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[86]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[87]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[88]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[89]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[8]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[90]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[91]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[92]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[93]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[94]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[95]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[96]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[97]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[98]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[99]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTDATA[9]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTKEEP[0]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTKEEP[1]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTKEEP[2]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTKEEP[3]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTKEEP[4]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTKEEP[5]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTKEEP[6]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTKEEP[7]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTLAST) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[0]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[10]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[11]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[12]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[13]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[14]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[15]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[16]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[17]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[18]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[19]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[1]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[20]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[21]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[22]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[23]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[24]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[25]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[26]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[27]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[28]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[29]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[2]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[30]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[31]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[32]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[33]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[34]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[35]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[36]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[37]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[38]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[39]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[3]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[40]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[41]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[42]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[43]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[44]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[45]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[46]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[47]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[48]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[49]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[4]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[50]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[51]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[52]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[53]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[54]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[55]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[56]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[57]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[58]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[59]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[5]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[60]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[61]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[62]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[63]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[64]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[65]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[66]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[67]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[68]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[69]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[6]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[70]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[71]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[72]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[73]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[74]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[7]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[8]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTUSER[9]) = (0:0:0, 0:0:0);
    (USERCLK => MAXISRCTVALID) = (0:0:0, 0:0:0);
    (USERCLK => PCIECQNPREQCOUNT[0]) = (0:0:0, 0:0:0);
    (USERCLK => PCIECQNPREQCOUNT[1]) = (0:0:0, 0:0:0);
    (USERCLK => PCIECQNPREQCOUNT[2]) = (0:0:0, 0:0:0);
    (USERCLK => PCIECQNPREQCOUNT[3]) = (0:0:0, 0:0:0);
    (USERCLK => PCIECQNPREQCOUNT[4]) = (0:0:0, 0:0:0);
    (USERCLK => PCIECQNPREQCOUNT[5]) = (0:0:0, 0:0:0);
    (USERCLK => PCIERQSEQNUMVLD) = (0:0:0, 0:0:0);
    (USERCLK => PCIERQSEQNUM[0]) = (0:0:0, 0:0:0);
    (USERCLK => PCIERQSEQNUM[1]) = (0:0:0, 0:0:0);
    (USERCLK => PCIERQSEQNUM[2]) = (0:0:0, 0:0:0);
    (USERCLK => PCIERQSEQNUM[3]) = (0:0:0, 0:0:0);
    (USERCLK => PCIERQTAGAV[0]) = (0:0:0, 0:0:0);
    (USERCLK => PCIERQTAGAV[1]) = (0:0:0, 0:0:0);
    (USERCLK => PCIERQTAGVLD) = (0:0:0, 0:0:0);
    (USERCLK => PCIERQTAG[0]) = (0:0:0, 0:0:0);
    (USERCLK => PCIERQTAG[1]) = (0:0:0, 0:0:0);
    (USERCLK => PCIERQTAG[2]) = (0:0:0, 0:0:0);
    (USERCLK => PCIERQTAG[3]) = (0:0:0, 0:0:0);
    (USERCLK => PCIERQTAG[4]) = (0:0:0, 0:0:0);
    (USERCLK => PCIERQTAG[5]) = (0:0:0, 0:0:0);
    (USERCLK => PCIETFCNPDAV[0]) = (0:0:0, 0:0:0);
    (USERCLK => PCIETFCNPDAV[1]) = (0:0:0, 0:0:0);
    (USERCLK => PCIETFCNPHAV[0]) = (0:0:0, 0:0:0);
    (USERCLK => PCIETFCNPHAV[1]) = (0:0:0, 0:0:0);
    (USERCLK => SAXISCCTREADY[0]) = (0:0:0, 0:0:0);
    (USERCLK => SAXISCCTREADY[1]) = (0:0:0, 0:0:0);
    (USERCLK => SAXISCCTREADY[2]) = (0:0:0, 0:0:0);
    (USERCLK => SAXISCCTREADY[3]) = (0:0:0, 0:0:0);
    (USERCLK => SAXISRQTREADY[0]) = (0:0:0, 0:0:0);
    (USERCLK => SAXISRQTREADY[1]) = (0:0:0, 0:0:0);
    (USERCLK => SAXISRQTREADY[2]) = (0:0:0, 0:0:0);
    (USERCLK => SAXISRQTREADY[3]) = (0:0:0, 0:0:0);
`ifdef XIL_TIMING // Simprim
    $period (negedge CORECLK, 0:0:0, notifier);
    $period (negedge CORECLKMICOMPLETIONRAML, 0:0:0, notifier);
    $period (negedge CORECLKMICOMPLETIONRAMU, 0:0:0, notifier);
    $period (negedge CORECLKMIREPLAYRAM, 0:0:0, notifier);
    $period (negedge CORECLKMIREQUESTRAM, 0:0:0, notifier);
    $period (negedge DRPCLK, 0:0:0, notifier);
    $period (negedge MCAPCLK, 0:0:0, notifier);
    $period (negedge PIPECLK, 0:0:0, notifier);
    $period (negedge USERCLK, 0:0:0, notifier);
    $period (posedge CORECLK, 0:0:0, notifier);
    $period (posedge CORECLKMICOMPLETIONRAML, 0:0:0, notifier);
    $period (posedge CORECLKMICOMPLETIONRAMU, 0:0:0, notifier);
    $period (posedge CORECLKMIREPLAYRAM, 0:0:0, notifier);
    $period (posedge CORECLKMIREQUESTRAM, 0:0:0, notifier);
    $period (posedge DRPCLK, 0:0:0, notifier);
    $period (posedge MCAPCLK, 0:0:0, notifier);
    $period (posedge PIPECLK, 0:0:0, notifier);
    $period (posedge USERCLK, 0:0:0, notifier);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[0], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[0]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[100], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[100]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[101], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[101]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[102], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[102]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[103], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[103]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[104], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[104]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[105], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[105]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[106], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[106]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[107], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[107]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[108], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[108]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[109], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[109]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[10], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[10]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[110], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[110]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[111], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[111]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[112], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[112]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[113], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[113]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[114], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[114]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[115], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[115]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[116], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[116]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[117], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[117]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[118], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[118]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[119], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[119]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[11], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[11]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[120], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[120]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[121], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[121]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[122], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[122]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[123], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[123]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[124], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[124]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[125], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[125]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[126], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[126]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[127], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[127]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[128], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[128]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[129], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[129]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[12], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[12]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[130], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[130]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[131], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[131]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[132], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[132]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[133], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[133]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[134], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[134]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[135], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[135]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[136], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[136]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[137], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[137]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[138], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[138]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[139], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[139]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[13], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[13]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[140], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[140]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[141], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[141]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[142], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[142]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[143], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[143]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[14], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[14]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[15], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[15]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[16], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[16]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[17], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[17]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[18], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[18]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[19], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[19]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[1], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[1]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[20], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[20]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[21], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[21]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[22], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[22]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[23], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[23]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[24], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[24]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[25], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[25]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[26], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[26]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[27], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[27]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[28], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[28]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[29], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[29]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[2], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[2]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[30], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[30]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[31], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[31]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[32], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[32]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[33], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[33]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[34], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[34]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[35], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[35]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[36], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[36]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[37], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[37]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[38], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[38]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[39], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[39]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[3], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[3]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[40], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[40]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[41], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[41]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[42], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[42]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[43], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[43]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[44], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[44]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[45], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[45]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[46], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[46]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[47], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[47]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[48], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[48]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[49], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[49]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[4], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[4]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[50], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[50]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[51], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[51]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[52], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[52]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[53], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[53]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[54], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[54]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[55], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[55]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[56], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[56]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[57], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[57]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[58], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[58]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[59], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[59]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[5], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[5]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[60], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[60]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[61], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[61]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[62], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[62]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[63], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[63]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[64], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[64]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[65], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[65]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[66], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[66]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[67], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[67]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[68], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[68]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[69], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[69]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[6], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[6]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[70], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[70]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[71], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[71]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[72], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[72]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[73], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[73]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[74], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[74]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[75], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[75]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[76], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[76]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[77], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[77]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[78], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[78]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[79], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[79]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[7], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[7]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[80], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[80]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[81], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[81]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[82], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[82]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[83], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[83]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[84], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[84]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[85], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[85]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[86], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[86]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[87], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[87]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[88], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[88]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[89], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[89]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[8], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[8]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[90], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[90]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[91], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[91]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[92], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[92]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[93], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[93]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[94], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[94]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[95], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[95]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[96], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[96]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[97], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[97]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[98], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[98]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[99], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[99]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[9], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[9]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[0], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[0]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[100], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[100]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[101], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[101]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[102], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[102]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[103], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[103]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[104], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[104]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[105], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[105]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[106], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[106]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[107], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[107]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[108], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[108]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[109], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[109]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[10], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[10]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[110], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[110]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[111], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[111]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[112], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[112]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[113], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[113]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[114], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[114]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[115], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[115]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[116], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[116]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[117], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[117]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[118], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[118]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[119], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[119]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[11], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[11]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[120], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[120]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[121], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[121]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[122], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[122]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[123], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[123]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[124], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[124]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[125], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[125]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[126], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[126]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[127], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[127]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[128], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[128]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[129], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[129]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[12], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[12]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[130], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[130]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[131], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[131]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[132], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[132]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[133], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[133]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[134], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[134]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[135], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[135]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[136], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[136]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[137], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[137]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[138], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[138]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[139], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[139]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[13], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[13]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[140], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[140]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[141], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[141]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[142], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[142]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[143], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[143]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[14], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[14]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[15], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[15]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[16], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[16]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[17], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[17]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[18], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[18]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[19], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[19]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[1], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[1]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[20], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[20]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[21], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[21]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[22], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[22]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[23], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[23]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[24], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[24]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[25], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[25]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[26], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[26]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[27], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[27]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[28], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[28]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[29], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[29]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[2], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[2]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[30], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[30]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[31], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[31]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[32], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[32]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[33], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[33]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[34], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[34]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[35], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[35]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[36], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[36]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[37], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[37]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[38], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[38]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[39], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[39]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[3], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[3]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[40], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[40]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[41], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[41]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[42], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[42]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[43], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[43]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[44], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[44]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[45], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[45]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[46], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[46]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[47], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[47]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[48], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[48]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[49], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[49]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[4], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[4]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[50], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[50]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[51], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[51]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[52], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[52]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[53], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[53]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[54], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[54]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[55], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[55]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[56], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[56]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[57], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[57]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[58], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[58]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[59], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[59]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[5], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[5]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[60], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[60]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[61], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[61]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[62], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[62]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[63], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[63]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[64], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[64]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[65], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[65]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[66], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[66]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[67], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[67]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[68], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[68]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[69], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[69]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[6], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[6]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[70], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[70]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[71], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[71]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[72], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[72]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[73], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[73]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[74], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[74]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[75], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[75]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[76], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[76]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[77], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[77]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[78], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[78]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[79], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[79]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[7], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[7]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[80], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[80]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[81], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[81]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[82], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[82]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[83], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[83]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[84], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[84]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[85], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[85]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[86], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[86]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[87], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[87]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[88], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[88]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[89], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[89]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[8], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[8]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[90], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[90]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[91], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[91]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[92], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[92]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[93], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[93]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[94], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[94]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[95], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[95]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[96], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[96]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[97], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[97]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[98], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[98]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[99], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[99]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[9], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[9]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[0], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[0]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[100], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[100]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[101], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[101]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[102], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[102]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[103], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[103]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[104], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[104]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[105], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[105]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[106], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[106]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[107], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[107]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[108], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[108]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[109], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[109]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[10], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[10]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[110], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[110]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[111], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[111]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[112], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[112]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[113], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[113]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[114], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[114]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[115], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[115]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[116], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[116]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[117], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[117]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[118], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[118]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[119], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[119]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[11], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[11]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[120], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[120]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[121], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[121]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[122], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[122]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[123], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[123]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[124], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[124]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[125], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[125]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[126], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[126]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[127], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[127]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[128], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[128]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[129], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[129]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[12], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[12]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[130], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[130]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[131], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[131]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[132], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[132]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[133], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[133]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[134], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[134]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[135], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[135]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[136], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[136]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[137], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[137]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[138], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[138]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[139], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[139]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[13], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[13]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[140], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[140]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[141], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[141]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[142], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[142]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[143], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[143]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[14], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[14]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[15], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[15]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[16], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[16]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[17], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[17]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[18], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[18]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[19], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[19]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[1], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[1]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[20], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[20]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[21], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[21]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[22], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[22]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[23], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[23]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[24], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[24]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[25], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[25]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[26], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[26]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[27], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[27]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[28], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[28]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[29], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[29]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[2], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[2]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[30], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[30]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[31], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[31]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[32], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[32]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[33], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[33]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[34], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[34]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[35], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[35]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[36], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[36]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[37], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[37]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[38], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[38]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[39], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[39]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[3], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[3]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[40], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[40]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[41], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[41]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[42], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[42]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[43], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[43]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[44], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[44]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[45], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[45]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[46], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[46]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[47], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[47]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[48], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[48]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[49], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[49]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[4], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[4]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[50], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[50]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[51], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[51]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[52], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[52]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[53], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[53]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[54], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[54]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[55], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[55]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[56], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[56]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[57], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[57]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[58], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[58]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[59], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[59]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[5], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[5]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[60], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[60]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[61], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[61]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[62], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[62]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[63], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[63]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[64], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[64]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[65], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[65]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[66], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[66]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[67], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[67]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[68], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[68]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[69], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[69]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[6], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[6]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[70], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[70]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[71], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[71]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[72], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[72]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[73], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[73]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[74], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[74]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[75], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[75]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[76], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[76]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[77], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[77]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[78], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[78]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[79], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[79]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[7], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[7]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[80], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[80]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[81], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[81]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[82], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[82]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[83], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[83]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[84], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[84]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[85], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[85]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[86], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[86]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[87], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[87]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[88], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[88]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[89], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[89]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[8], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[8]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[90], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[90]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[91], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[91]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[92], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[92]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[93], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[93]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[94], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[94]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[95], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[95]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[96], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[96]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[97], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[97]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[98], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[98]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[99], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[99]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[9], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[9]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[0], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[0]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[100], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[100]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[101], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[101]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[102], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[102]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[103], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[103]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[104], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[104]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[105], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[105]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[106], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[106]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[107], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[107]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[108], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[108]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[109], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[109]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[10], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[10]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[110], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[110]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[111], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[111]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[112], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[112]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[113], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[113]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[114], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[114]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[115], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[115]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[116], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[116]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[117], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[117]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[118], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[118]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[119], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[119]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[11], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[11]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[120], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[120]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[121], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[121]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[122], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[122]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[123], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[123]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[124], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[124]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[125], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[125]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[126], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[126]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[127], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[127]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[128], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[128]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[129], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[129]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[12], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[12]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[130], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[130]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[131], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[131]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[132], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[132]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[133], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[133]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[134], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[134]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[135], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[135]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[136], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[136]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[137], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[137]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[138], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[138]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[139], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[139]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[13], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[13]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[140], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[140]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[141], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[141]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[142], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[142]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[143], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[143]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[14], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[14]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[15], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[15]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[16], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[16]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[17], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[17]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[18], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[18]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[19], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[19]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[1], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[1]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[20], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[20]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[21], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[21]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[22], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[22]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[23], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[23]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[24], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[24]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[25], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[25]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[26], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[26]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[27], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[27]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[28], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[28]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[29], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[29]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[2], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[2]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[30], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[30]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[31], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[31]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[32], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[32]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[33], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[33]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[34], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[34]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[35], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[35]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[36], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[36]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[37], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[37]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[38], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[38]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[39], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[39]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[3], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[3]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[40], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[40]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[41], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[41]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[42], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[42]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[43], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[43]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[44], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[44]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[45], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[45]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[46], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[46]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[47], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[47]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[48], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[48]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[49], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[49]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[4], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[4]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[50], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[50]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[51], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[51]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[52], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[52]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[53], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[53]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[54], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[54]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[55], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[55]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[56], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[56]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[57], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[57]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[58], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[58]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[59], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[59]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[5], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[5]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[60], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[60]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[61], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[61]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[62], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[62]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[63], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[63]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[64], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[64]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[65], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[65]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[66], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[66]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[67], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[67]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[68], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[68]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[69], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[69]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[6], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[6]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[70], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[70]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[71], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[71]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[72], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[72]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[73], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[73]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[74], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[74]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[75], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[75]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[76], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[76]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[77], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[77]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[78], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[78]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[79], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[79]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[7], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[7]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[80], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[80]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[81], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[81]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[82], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[82]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[83], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[83]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[84], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[84]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[85], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[85]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[86], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[86]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[87], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[87]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[88], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[88]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[89], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[89]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[8], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[8]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[90], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[90]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[91], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[91]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[92], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[92]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[93], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[93]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[94], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[94]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[95], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[95]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[96], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[96]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[97], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[97]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[98], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[98]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[99], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[99]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[9], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MICOMPLETIONRAMREADDATA_delay[9]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[0], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[0]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[100], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[100]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[101], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[101]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[102], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[102]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[103], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[103]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[104], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[104]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[105], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[105]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[106], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[106]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[107], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[107]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[108], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[108]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[109], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[109]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[10], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[10]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[110], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[110]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[111], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[111]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[112], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[112]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[113], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[113]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[114], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[114]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[115], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[115]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[116], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[116]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[117], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[117]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[118], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[118]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[119], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[119]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[11], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[11]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[120], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[120]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[121], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[121]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[122], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[122]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[123], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[123]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[124], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[124]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[125], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[125]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[126], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[126]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[127], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[127]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[128], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[128]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[129], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[129]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[12], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[12]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[130], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[130]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[131], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[131]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[132], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[132]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[133], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[133]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[134], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[134]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[135], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[135]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[136], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[136]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[137], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[137]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[138], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[138]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[139], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[139]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[13], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[13]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[140], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[140]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[141], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[141]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[142], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[142]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[143], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[143]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[14], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[14]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[15], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[15]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[16], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[16]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[17], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[17]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[18], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[18]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[19], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[19]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[1], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[1]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[20], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[20]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[21], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[21]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[22], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[22]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[23], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[23]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[24], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[24]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[25], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[25]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[26], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[26]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[27], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[27]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[28], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[28]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[29], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[29]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[2], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[2]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[30], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[30]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[31], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[31]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[32], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[32]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[33], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[33]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[34], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[34]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[35], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[35]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[36], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[36]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[37], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[37]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[38], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[38]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[39], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[39]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[3], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[3]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[40], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[40]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[41], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[41]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[42], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[42]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[43], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[43]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[44], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[44]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[45], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[45]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[46], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[46]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[47], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[47]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[48], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[48]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[49], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[49]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[4], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[4]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[50], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[50]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[51], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[51]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[52], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[52]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[53], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[53]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[54], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[54]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[55], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[55]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[56], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[56]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[57], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[57]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[58], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[58]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[59], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[59]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[5], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[5]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[60], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[60]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[61], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[61]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[62], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[62]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[63], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[63]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[64], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[64]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[65], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[65]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[66], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[66]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[67], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[67]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[68], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[68]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[69], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[69]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[6], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[6]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[70], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[70]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[71], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[71]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[72], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[72]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[73], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[73]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[74], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[74]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[75], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[75]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[76], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[76]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[77], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[77]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[78], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[78]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[79], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[79]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[7], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[7]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[80], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[80]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[81], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[81]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[82], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[82]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[83], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[83]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[84], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[84]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[85], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[85]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[86], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[86]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[87], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[87]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[88], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[88]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[89], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[89]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[8], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[8]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[90], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[90]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[91], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[91]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[92], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[92]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[93], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[93]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[94], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[94]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[95], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[95]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[96], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[96]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[97], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[97]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[98], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[98]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[99], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[99]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[9], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREPLAYRAMREADDATA_delay[9]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[0], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[0]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[100], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[100]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[101], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[101]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[102], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[102]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[103], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[103]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[104], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[104]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[105], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[105]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[106], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[106]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[107], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[107]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[108], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[108]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[109], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[109]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[10], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[10]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[110], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[110]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[111], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[111]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[112], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[112]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[113], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[113]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[114], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[114]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[115], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[115]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[116], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[116]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[117], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[117]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[118], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[118]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[119], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[119]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[11], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[11]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[120], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[120]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[121], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[121]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[122], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[122]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[123], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[123]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[124], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[124]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[125], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[125]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[126], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[126]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[127], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[127]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[128], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[128]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[129], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[129]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[12], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[12]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[130], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[130]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[131], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[131]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[132], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[132]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[133], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[133]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[134], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[134]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[135], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[135]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[136], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[136]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[137], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[137]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[138], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[138]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[139], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[139]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[13], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[13]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[140], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[140]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[141], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[141]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[142], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[142]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[143], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[143]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[14], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[14]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[15], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[15]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[16], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[16]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[17], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[17]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[18], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[18]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[19], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[19]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[1], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[1]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[20], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[20]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[21], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[21]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[22], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[22]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[23], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[23]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[24], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[24]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[25], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[25]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[26], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[26]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[27], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[27]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[28], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[28]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[29], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[29]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[2], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[2]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[30], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[30]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[31], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[31]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[32], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[32]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[33], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[33]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[34], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[34]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[35], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[35]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[36], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[36]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[37], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[37]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[38], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[38]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[39], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[39]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[3], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[3]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[40], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[40]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[41], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[41]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[42], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[42]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[43], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[43]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[44], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[44]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[45], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[45]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[46], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[46]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[47], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[47]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[48], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[48]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[49], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[49]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[4], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[4]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[50], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[50]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[51], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[51]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[52], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[52]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[53], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[53]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[54], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[54]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[55], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[55]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[56], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[56]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[57], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[57]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[58], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[58]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[59], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[59]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[5], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[5]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[60], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[60]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[61], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[61]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[62], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[62]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[63], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[63]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[64], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[64]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[65], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[65]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[66], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[66]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[67], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[67]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[68], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[68]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[69], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[69]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[6], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[6]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[70], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[70]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[71], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[71]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[72], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[72]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[73], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[73]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[74], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[74]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[75], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[75]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[76], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[76]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[77], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[77]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[78], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[78]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[79], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[79]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[7], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[7]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[80], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[80]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[81], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[81]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[82], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[82]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[83], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[83]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[84], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[84]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[85], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[85]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[86], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[86]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[87], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[87]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[88], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[88]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[89], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[89]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[8], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[8]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[90], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[90]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[91], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[91]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[92], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[92]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[93], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[93]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[94], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[94]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[95], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[95]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[96], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[96]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[97], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[97]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[98], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[98]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[99], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[99]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[9], 0:0:0, 0:0:0, notifier,,, CORECLK_delay, MIREQUESTRAMREADDATA_delay[9]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[0], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPADDR_delay[0]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[1], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPADDR_delay[1]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[2], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPADDR_delay[2]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[3], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPADDR_delay[3]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[4], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPADDR_delay[4]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[5], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPADDR_delay[5]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[6], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPADDR_delay[6]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[7], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPADDR_delay[7]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[8], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPADDR_delay[8]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[9], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPADDR_delay[9]);
    $setuphold (posedge DRPCLK, negedge DRPDI[0], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[0]);
    $setuphold (posedge DRPCLK, negedge DRPDI[10], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[10]);
    $setuphold (posedge DRPCLK, negedge DRPDI[11], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[11]);
    $setuphold (posedge DRPCLK, negedge DRPDI[12], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[12]);
    $setuphold (posedge DRPCLK, negedge DRPDI[13], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[13]);
    $setuphold (posedge DRPCLK, negedge DRPDI[14], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[14]);
    $setuphold (posedge DRPCLK, negedge DRPDI[15], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[15]);
    $setuphold (posedge DRPCLK, negedge DRPDI[1], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[1]);
    $setuphold (posedge DRPCLK, negedge DRPDI[2], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[2]);
    $setuphold (posedge DRPCLK, negedge DRPDI[3], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[3]);
    $setuphold (posedge DRPCLK, negedge DRPDI[4], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[4]);
    $setuphold (posedge DRPCLK, negedge DRPDI[5], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[5]);
    $setuphold (posedge DRPCLK, negedge DRPDI[6], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[6]);
    $setuphold (posedge DRPCLK, negedge DRPDI[7], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[7]);
    $setuphold (posedge DRPCLK, negedge DRPDI[8], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[8]);
    $setuphold (posedge DRPCLK, negedge DRPDI[9], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[9]);
    $setuphold (posedge DRPCLK, negedge DRPEN, 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPEN_delay);
    $setuphold (posedge DRPCLK, negedge DRPWE, 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPWE_delay);
    $setuphold (posedge DRPCLK, posedge DRPADDR[0], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPADDR_delay[0]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[1], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPADDR_delay[1]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[2], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPADDR_delay[2]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[3], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPADDR_delay[3]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[4], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPADDR_delay[4]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[5], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPADDR_delay[5]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[6], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPADDR_delay[6]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[7], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPADDR_delay[7]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[8], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPADDR_delay[8]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[9], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPADDR_delay[9]);
    $setuphold (posedge DRPCLK, posedge DRPDI[0], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[0]);
    $setuphold (posedge DRPCLK, posedge DRPDI[10], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[10]);
    $setuphold (posedge DRPCLK, posedge DRPDI[11], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[11]);
    $setuphold (posedge DRPCLK, posedge DRPDI[12], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[12]);
    $setuphold (posedge DRPCLK, posedge DRPDI[13], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[13]);
    $setuphold (posedge DRPCLK, posedge DRPDI[14], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[14]);
    $setuphold (posedge DRPCLK, posedge DRPDI[15], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[15]);
    $setuphold (posedge DRPCLK, posedge DRPDI[1], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[1]);
    $setuphold (posedge DRPCLK, posedge DRPDI[2], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[2]);
    $setuphold (posedge DRPCLK, posedge DRPDI[3], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[3]);
    $setuphold (posedge DRPCLK, posedge DRPDI[4], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[4]);
    $setuphold (posedge DRPCLK, posedge DRPDI[5], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[5]);
    $setuphold (posedge DRPCLK, posedge DRPDI[6], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[6]);
    $setuphold (posedge DRPCLK, posedge DRPDI[7], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[7]);
    $setuphold (posedge DRPCLK, posedge DRPDI[8], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[8]);
    $setuphold (posedge DRPCLK, posedge DRPDI[9], 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPDI_delay[9]);
    $setuphold (posedge DRPCLK, posedge DRPEN, 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPEN_delay);
    $setuphold (posedge DRPCLK, posedge DRPWE, 0:0:0, 0:0:0, notifier,,, DRPCLK_delay, DRPWE_delay);
    $setuphold (posedge PIPECLK, negedge PIPEEQFS[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPEEQFS_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPEEQFS[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPEEQFS_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPEEQFS[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPEEQFS_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPEEQFS[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPEEQFS_delay[3]);
    $setuphold (posedge PIPECLK, negedge PIPEEQFS[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPEEQFS_delay[4]);
    $setuphold (posedge PIPECLK, negedge PIPEEQFS[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPEEQFS_delay[5]);
    $setuphold (posedge PIPECLK, negedge PIPEEQLF[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPEEQLF_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPEEQLF[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPEEQLF_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPEEQLF[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPEEQLF_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPEEQLF[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPEEQLF_delay[3]);
    $setuphold (posedge PIPECLK, negedge PIPEEQLF[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPEEQLF_delay[4]);
    $setuphold (posedge PIPECLK, negedge PIPEEQLF[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPEEQLF_delay[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX0CHARISK[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0CHARISK_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX0CHARISK[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0CHARISK_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATAVALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATAVALID_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[18], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[18]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[19], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[19]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[20], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[20]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[21], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[21]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[22], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[22]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[23], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[23]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[24], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[24]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[25], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[25]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[26], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[26]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[27], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[27]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[28], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[28]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[29], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[29]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[30], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[30]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[31], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[31]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX0ELECIDLE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0ELECIDLE_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQDONE_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPADAPTDONE_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPLFFSSEL_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX0PHYSTATUS, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0PHYSTATUS_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX0STARTBLOCK, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0STARTBLOCK_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX0STATUS[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0STATUS_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX0STATUS[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0STATUS_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX0STATUS[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0STATUS_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX0SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0SYNCHEADER_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX0SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0SYNCHEADER_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX0VALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0VALID_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX1CHARISK[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1CHARISK_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX1CHARISK[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1CHARISK_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATAVALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATAVALID_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[18], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[18]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[19], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[19]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[20], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[20]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[21], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[21]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[22], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[22]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[23], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[23]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[24], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[24]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[25], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[25]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[26], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[26]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[27], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[27]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[28], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[28]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[29], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[29]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[30], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[30]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[31], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[31]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX1ELECIDLE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1ELECIDLE_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQDONE_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPADAPTDONE_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPLFFSSEL_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX1PHYSTATUS, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1PHYSTATUS_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX1STARTBLOCK, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1STARTBLOCK_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX1STATUS[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1STATUS_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX1STATUS[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1STATUS_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX1STATUS[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1STATUS_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX1SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1SYNCHEADER_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX1SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1SYNCHEADER_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX1VALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1VALID_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX2CHARISK[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2CHARISK_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX2CHARISK[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2CHARISK_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATAVALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATAVALID_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[18], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[18]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[19], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[19]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[20], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[20]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[21], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[21]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[22], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[22]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[23], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[23]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[24], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[24]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[25], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[25]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[26], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[26]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[27], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[27]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[28], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[28]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[29], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[29]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[30], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[30]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[31], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[31]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX2ELECIDLE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2ELECIDLE_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQDONE_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPADAPTDONE_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPLFFSSEL_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX2PHYSTATUS, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2PHYSTATUS_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX2STARTBLOCK, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2STARTBLOCK_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX2STATUS[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2STATUS_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX2STATUS[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2STATUS_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX2STATUS[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2STATUS_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX2SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2SYNCHEADER_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX2SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2SYNCHEADER_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX2VALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2VALID_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX3CHARISK[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3CHARISK_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX3CHARISK[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3CHARISK_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATAVALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATAVALID_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[18], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[18]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[19], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[19]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[20], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[20]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[21], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[21]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[22], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[22]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[23], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[23]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[24], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[24]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[25], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[25]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[26], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[26]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[27], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[27]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[28], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[28]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[29], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[29]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[30], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[30]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[31], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[31]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX3ELECIDLE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3ELECIDLE_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQDONE_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPADAPTDONE_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPLFFSSEL_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX3PHYSTATUS, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3PHYSTATUS_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX3STARTBLOCK, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3STARTBLOCK_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX3STATUS[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3STATUS_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX3STATUS[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3STATUS_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX3STATUS[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3STATUS_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX3SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3SYNCHEADER_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX3SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3SYNCHEADER_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX3VALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3VALID_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX4CHARISK[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4CHARISK_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX4CHARISK[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4CHARISK_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATAVALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATAVALID_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[18], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[18]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[19], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[19]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[20], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[20]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[21], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[21]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[22], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[22]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[23], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[23]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[24], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[24]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[25], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[25]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[26], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[26]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[27], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[27]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[28], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[28]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[29], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[29]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[30], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[30]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[31], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[31]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX4ELECIDLE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4ELECIDLE_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQDONE_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPADAPTDONE_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPLFFSSEL_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX4PHYSTATUS, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4PHYSTATUS_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX4STARTBLOCK, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4STARTBLOCK_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX4STATUS[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4STATUS_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX4STATUS[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4STATUS_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX4STATUS[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4STATUS_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX4SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4SYNCHEADER_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX4SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4SYNCHEADER_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX4VALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4VALID_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX5CHARISK[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5CHARISK_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX5CHARISK[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5CHARISK_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATAVALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATAVALID_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[18], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[18]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[19], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[19]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[20], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[20]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[21], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[21]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[22], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[22]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[23], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[23]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[24], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[24]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[25], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[25]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[26], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[26]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[27], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[27]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[28], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[28]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[29], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[29]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[30], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[30]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[31], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[31]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX5ELECIDLE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5ELECIDLE_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQDONE_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPADAPTDONE_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPLFFSSEL_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX5PHYSTATUS, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5PHYSTATUS_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX5STARTBLOCK, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5STARTBLOCK_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX5STATUS[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5STATUS_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX5STATUS[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5STATUS_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX5STATUS[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5STATUS_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX5SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5SYNCHEADER_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX5SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5SYNCHEADER_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX5VALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5VALID_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX6CHARISK[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6CHARISK_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX6CHARISK[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6CHARISK_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATAVALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATAVALID_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[18], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[18]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[19], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[19]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[20], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[20]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[21], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[21]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[22], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[22]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[23], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[23]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[24], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[24]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[25], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[25]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[26], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[26]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[27], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[27]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[28], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[28]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[29], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[29]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[30], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[30]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[31], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[31]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX6ELECIDLE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6ELECIDLE_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQDONE_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPADAPTDONE_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPLFFSSEL_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX6PHYSTATUS, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6PHYSTATUS_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX6STARTBLOCK, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6STARTBLOCK_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX6STATUS[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6STATUS_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX6STATUS[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6STATUS_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX6STATUS[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6STATUS_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX6SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6SYNCHEADER_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX6SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6SYNCHEADER_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX6VALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6VALID_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX7CHARISK[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7CHARISK_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX7CHARISK[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7CHARISK_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATAVALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATAVALID_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[18], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[18]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[19], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[19]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[20], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[20]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[21], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[21]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[22], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[22]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[23], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[23]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[24], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[24]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[25], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[25]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[26], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[26]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[27], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[27]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[28], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[28]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[29], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[29]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[30], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[30]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[31], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[31]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX7ELECIDLE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7ELECIDLE_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQDONE_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPADAPTDONE_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPLFFSSEL_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX7PHYSTATUS, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7PHYSTATUS_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX7STARTBLOCK, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7STARTBLOCK_delay);
    $setuphold (posedge PIPECLK, negedge PIPERX7STATUS[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7STATUS_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX7STATUS[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7STATUS_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX7STATUS[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7STATUS_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX7SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7SYNCHEADER_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX7SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7SYNCHEADER_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX7VALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7VALID_delay);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[10]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[11]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[12]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[13]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[14]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[15]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[16]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[17]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[3]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[4]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[5]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[6]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[7]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[8]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[9]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQDONE_delay);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[10]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[11]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[12]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[13]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[14]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[15]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[16]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[17]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[3]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[4]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[5]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[6]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[7]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[8]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[9]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQDONE_delay);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[10]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[11]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[12]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[13]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[14]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[15]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[16]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[17]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[3]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[4]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[5]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[6]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[7]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[8]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[9]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQDONE_delay);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[10]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[11]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[12]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[13]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[14]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[15]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[16]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[17]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[3]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[4]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[5]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[6]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[7]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[8]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[9]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQDONE_delay);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[10]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[11]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[12]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[13]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[14]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[15]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[16]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[17]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[3]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[4]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[5]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[6]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[7]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[8]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[9]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQDONE_delay);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[10]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[11]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[12]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[13]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[14]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[15]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[16]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[17]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[3]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[4]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[5]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[6]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[7]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[8]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[9]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQDONE_delay);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[10]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[11]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[12]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[13]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[14]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[15]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[16]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[17]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[3]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[4]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[5]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[6]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[7]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[8]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[9]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQDONE_delay);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[0]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[10]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[11]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[12]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[13]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[14]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[15]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[16]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[17]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[1]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[2]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[3]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[4]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[5]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[6]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[7]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[8]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[9]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQDONE_delay);
    $setuphold (posedge PIPECLK, negedge PLEQRESETEIEOSCOUNT, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PLEQRESETEIEOSCOUNT_delay);
    $setuphold (posedge PIPECLK, negedge PLGEN2UPSTREAMPREFERDEEMPH, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PLGEN2UPSTREAMPREFERDEEMPH_delay);
    $setuphold (posedge PIPECLK, posedge PIPEEQFS[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPEEQFS_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPEEQFS[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPEEQFS_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPEEQFS[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPEEQFS_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPEEQFS[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPEEQFS_delay[3]);
    $setuphold (posedge PIPECLK, posedge PIPEEQFS[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPEEQFS_delay[4]);
    $setuphold (posedge PIPECLK, posedge PIPEEQFS[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPEEQFS_delay[5]);
    $setuphold (posedge PIPECLK, posedge PIPEEQLF[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPEEQLF_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPEEQLF[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPEEQLF_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPEEQLF[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPEEQLF_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPEEQLF[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPEEQLF_delay[3]);
    $setuphold (posedge PIPECLK, posedge PIPEEQLF[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPEEQLF_delay[4]);
    $setuphold (posedge PIPECLK, posedge PIPEEQLF[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPEEQLF_delay[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX0CHARISK[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0CHARISK_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX0CHARISK[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0CHARISK_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATAVALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATAVALID_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[18], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[18]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[19], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[19]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[20], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[20]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[21], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[21]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[22], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[22]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[23], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[23]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[24], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[24]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[25], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[25]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[26], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[26]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[27], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[27]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[28], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[28]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[29], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[29]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[30], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[30]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[31], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[31]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0DATA_delay[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX0ELECIDLE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0ELECIDLE_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQDONE_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPADAPTDONE_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPLFFSSEL_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0EQLPNEWTXCOEFFORPRESET_delay[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX0PHYSTATUS, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0PHYSTATUS_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX0STARTBLOCK, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0STARTBLOCK_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX0STATUS[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0STATUS_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX0STATUS[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0STATUS_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX0STATUS[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0STATUS_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX0SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0SYNCHEADER_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX0SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0SYNCHEADER_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX0VALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX0VALID_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX1CHARISK[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1CHARISK_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX1CHARISK[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1CHARISK_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATAVALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATAVALID_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[18], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[18]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[19], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[19]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[20], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[20]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[21], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[21]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[22], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[22]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[23], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[23]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[24], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[24]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[25], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[25]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[26], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[26]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[27], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[27]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[28], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[28]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[29], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[29]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[30], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[30]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[31], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[31]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1DATA_delay[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX1ELECIDLE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1ELECIDLE_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQDONE_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPADAPTDONE_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPLFFSSEL_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1EQLPNEWTXCOEFFORPRESET_delay[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX1PHYSTATUS, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1PHYSTATUS_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX1STARTBLOCK, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1STARTBLOCK_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX1STATUS[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1STATUS_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX1STATUS[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1STATUS_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX1STATUS[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1STATUS_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX1SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1SYNCHEADER_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX1SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1SYNCHEADER_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX1VALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX1VALID_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX2CHARISK[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2CHARISK_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX2CHARISK[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2CHARISK_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATAVALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATAVALID_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[18], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[18]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[19], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[19]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[20], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[20]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[21], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[21]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[22], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[22]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[23], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[23]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[24], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[24]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[25], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[25]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[26], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[26]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[27], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[27]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[28], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[28]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[29], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[29]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[30], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[30]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[31], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[31]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2DATA_delay[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX2ELECIDLE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2ELECIDLE_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQDONE_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPADAPTDONE_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPLFFSSEL_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2EQLPNEWTXCOEFFORPRESET_delay[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX2PHYSTATUS, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2PHYSTATUS_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX2STARTBLOCK, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2STARTBLOCK_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX2STATUS[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2STATUS_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX2STATUS[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2STATUS_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX2STATUS[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2STATUS_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX2SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2SYNCHEADER_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX2SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2SYNCHEADER_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX2VALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX2VALID_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX3CHARISK[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3CHARISK_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX3CHARISK[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3CHARISK_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATAVALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATAVALID_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[18], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[18]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[19], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[19]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[20], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[20]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[21], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[21]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[22], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[22]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[23], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[23]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[24], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[24]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[25], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[25]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[26], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[26]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[27], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[27]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[28], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[28]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[29], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[29]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[30], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[30]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[31], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[31]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3DATA_delay[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX3ELECIDLE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3ELECIDLE_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQDONE_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPADAPTDONE_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPLFFSSEL_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3EQLPNEWTXCOEFFORPRESET_delay[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX3PHYSTATUS, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3PHYSTATUS_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX3STARTBLOCK, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3STARTBLOCK_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX3STATUS[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3STATUS_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX3STATUS[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3STATUS_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX3STATUS[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3STATUS_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX3SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3SYNCHEADER_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX3SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3SYNCHEADER_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX3VALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX3VALID_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX4CHARISK[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4CHARISK_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX4CHARISK[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4CHARISK_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATAVALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATAVALID_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[18], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[18]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[19], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[19]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[20], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[20]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[21], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[21]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[22], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[22]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[23], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[23]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[24], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[24]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[25], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[25]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[26], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[26]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[27], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[27]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[28], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[28]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[29], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[29]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[30], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[30]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[31], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[31]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4DATA_delay[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX4ELECIDLE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4ELECIDLE_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQDONE_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPADAPTDONE_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPLFFSSEL_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4EQLPNEWTXCOEFFORPRESET_delay[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX4PHYSTATUS, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4PHYSTATUS_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX4STARTBLOCK, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4STARTBLOCK_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX4STATUS[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4STATUS_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX4STATUS[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4STATUS_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX4STATUS[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4STATUS_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX4SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4SYNCHEADER_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX4SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4SYNCHEADER_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX4VALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX4VALID_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX5CHARISK[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5CHARISK_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX5CHARISK[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5CHARISK_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATAVALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATAVALID_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[18], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[18]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[19], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[19]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[20], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[20]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[21], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[21]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[22], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[22]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[23], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[23]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[24], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[24]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[25], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[25]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[26], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[26]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[27], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[27]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[28], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[28]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[29], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[29]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[30], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[30]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[31], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[31]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5DATA_delay[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX5ELECIDLE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5ELECIDLE_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQDONE_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPADAPTDONE_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPLFFSSEL_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5EQLPNEWTXCOEFFORPRESET_delay[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX5PHYSTATUS, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5PHYSTATUS_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX5STARTBLOCK, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5STARTBLOCK_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX5STATUS[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5STATUS_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX5STATUS[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5STATUS_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX5STATUS[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5STATUS_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX5SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5SYNCHEADER_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX5SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5SYNCHEADER_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX5VALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX5VALID_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX6CHARISK[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6CHARISK_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX6CHARISK[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6CHARISK_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATAVALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATAVALID_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[18], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[18]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[19], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[19]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[20], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[20]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[21], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[21]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[22], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[22]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[23], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[23]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[24], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[24]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[25], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[25]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[26], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[26]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[27], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[27]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[28], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[28]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[29], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[29]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[30], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[30]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[31], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[31]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6DATA_delay[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX6ELECIDLE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6ELECIDLE_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQDONE_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPADAPTDONE_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPLFFSSEL_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6EQLPNEWTXCOEFFORPRESET_delay[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX6PHYSTATUS, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6PHYSTATUS_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX6STARTBLOCK, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6STARTBLOCK_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX6STATUS[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6STATUS_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX6STATUS[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6STATUS_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX6STATUS[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6STATUS_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX6SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6SYNCHEADER_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX6SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6SYNCHEADER_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX6VALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX6VALID_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX7CHARISK[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7CHARISK_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX7CHARISK[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7CHARISK_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATAVALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATAVALID_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[18], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[18]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[19], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[19]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[20], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[20]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[21], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[21]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[22], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[22]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[23], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[23]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[24], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[24]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[25], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[25]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[26], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[26]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[27], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[27]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[28], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[28]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[29], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[29]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[30], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[30]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[31], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[31]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7DATA_delay[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX7ELECIDLE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7ELECIDLE_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQDONE_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPADAPTDONE_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPLFFSSEL_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7EQLPNEWTXCOEFFORPRESET_delay[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX7PHYSTATUS, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7PHYSTATUS_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX7STARTBLOCK, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7STARTBLOCK_delay);
    $setuphold (posedge PIPECLK, posedge PIPERX7STATUS[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7STATUS_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX7STATUS[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7STATUS_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX7STATUS[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7STATUS_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX7SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7SYNCHEADER_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX7SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7SYNCHEADER_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX7VALID, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPERX7VALID_delay);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[10]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[11]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[12]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[13]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[14]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[15]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[16]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[17]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[3]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[4]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[5]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[6]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[7]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[8]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQCOEFF_delay[9]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX0EQDONE_delay);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[10]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[11]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[12]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[13]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[14]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[15]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[16]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[17]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[3]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[4]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[5]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[6]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[7]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[8]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQCOEFF_delay[9]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX1EQDONE_delay);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[10]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[11]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[12]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[13]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[14]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[15]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[16]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[17]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[3]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[4]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[5]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[6]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[7]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[8]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQCOEFF_delay[9]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX2EQDONE_delay);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[10]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[11]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[12]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[13]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[14]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[15]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[16]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[17]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[3]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[4]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[5]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[6]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[7]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[8]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQCOEFF_delay[9]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX3EQDONE_delay);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[10]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[11]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[12]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[13]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[14]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[15]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[16]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[17]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[3]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[4]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[5]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[6]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[7]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[8]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQCOEFF_delay[9]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX4EQDONE_delay);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[10]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[11]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[12]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[13]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[14]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[15]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[16]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[17]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[3]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[4]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[5]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[6]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[7]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[8]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQCOEFF_delay[9]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX5EQDONE_delay);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[10]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[11]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[12]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[13]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[14]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[15]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[16]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[17]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[3]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[4]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[5]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[6]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[7]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[8]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQCOEFF_delay[9]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX6EQDONE_delay);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[0]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[10]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[11]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[12]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[13]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[14]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[15]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[16]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[17]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[1]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[2]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[3]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[4]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[5]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[6]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[7]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[8]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQCOEFF_delay[9]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQDONE, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PIPETX7EQDONE_delay);
    $setuphold (posedge PIPECLK, posedge PLEQRESETEIEOSCOUNT, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PLEQRESETEIEOSCOUNT_delay);
    $setuphold (posedge PIPECLK, posedge PLGEN2UPSTREAMPREFERDEEMPH, 0:0:0, 0:0:0, notifier,,, PIPECLK_delay, PLGEN2UPSTREAMPREFERDEEMPH_delay);
    $setuphold (posedge USERCLK, negedge CFGCONFIGSPACEENABLE, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGCONFIGSPACEENABLE_delay);
    $setuphold (posedge USERCLK, negedge CFGDEVID[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[10]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[11]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[12]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[13]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[14]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[15]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[3]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[4]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[5]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[6]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[7]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[8]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[9]);
    $setuphold (posedge USERCLK, negedge CFGDSBUSNUMBER[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSBUSNUMBER_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGDSBUSNUMBER[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSBUSNUMBER_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGDSBUSNUMBER[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSBUSNUMBER_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGDSBUSNUMBER[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSBUSNUMBER_delay[3]);
    $setuphold (posedge USERCLK, negedge CFGDSBUSNUMBER[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSBUSNUMBER_delay[4]);
    $setuphold (posedge USERCLK, negedge CFGDSBUSNUMBER[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSBUSNUMBER_delay[5]);
    $setuphold (posedge USERCLK, negedge CFGDSBUSNUMBER[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSBUSNUMBER_delay[6]);
    $setuphold (posedge USERCLK, negedge CFGDSBUSNUMBER[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSBUSNUMBER_delay[7]);
    $setuphold (posedge USERCLK, negedge CFGDSDEVICENUMBER[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSDEVICENUMBER_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGDSDEVICENUMBER[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSDEVICENUMBER_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGDSDEVICENUMBER[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSDEVICENUMBER_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGDSDEVICENUMBER[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSDEVICENUMBER_delay[3]);
    $setuphold (posedge USERCLK, negedge CFGDSDEVICENUMBER[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSDEVICENUMBER_delay[4]);
    $setuphold (posedge USERCLK, negedge CFGDSFUNCTIONNUMBER[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSFUNCTIONNUMBER_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGDSFUNCTIONNUMBER[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSFUNCTIONNUMBER_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGDSFUNCTIONNUMBER[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSFUNCTIONNUMBER_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGDSN[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGDSN[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[10]);
    $setuphold (posedge USERCLK, negedge CFGDSN[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[11]);
    $setuphold (posedge USERCLK, negedge CFGDSN[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[12]);
    $setuphold (posedge USERCLK, negedge CFGDSN[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[13]);
    $setuphold (posedge USERCLK, negedge CFGDSN[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[14]);
    $setuphold (posedge USERCLK, negedge CFGDSN[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[15]);
    $setuphold (posedge USERCLK, negedge CFGDSN[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[16]);
    $setuphold (posedge USERCLK, negedge CFGDSN[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[17]);
    $setuphold (posedge USERCLK, negedge CFGDSN[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[18]);
    $setuphold (posedge USERCLK, negedge CFGDSN[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[19]);
    $setuphold (posedge USERCLK, negedge CFGDSN[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGDSN[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[20]);
    $setuphold (posedge USERCLK, negedge CFGDSN[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[21]);
    $setuphold (posedge USERCLK, negedge CFGDSN[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[22]);
    $setuphold (posedge USERCLK, negedge CFGDSN[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[23]);
    $setuphold (posedge USERCLK, negedge CFGDSN[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[24]);
    $setuphold (posedge USERCLK, negedge CFGDSN[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[25]);
    $setuphold (posedge USERCLK, negedge CFGDSN[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[26]);
    $setuphold (posedge USERCLK, negedge CFGDSN[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[27]);
    $setuphold (posedge USERCLK, negedge CFGDSN[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[28]);
    $setuphold (posedge USERCLK, negedge CFGDSN[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[29]);
    $setuphold (posedge USERCLK, negedge CFGDSN[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGDSN[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[30]);
    $setuphold (posedge USERCLK, negedge CFGDSN[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[31]);
    $setuphold (posedge USERCLK, negedge CFGDSN[32], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[32]);
    $setuphold (posedge USERCLK, negedge CFGDSN[33], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[33]);
    $setuphold (posedge USERCLK, negedge CFGDSN[34], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[34]);
    $setuphold (posedge USERCLK, negedge CFGDSN[35], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[35]);
    $setuphold (posedge USERCLK, negedge CFGDSN[36], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[36]);
    $setuphold (posedge USERCLK, negedge CFGDSN[37], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[37]);
    $setuphold (posedge USERCLK, negedge CFGDSN[38], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[38]);
    $setuphold (posedge USERCLK, negedge CFGDSN[39], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[39]);
    $setuphold (posedge USERCLK, negedge CFGDSN[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[3]);
    $setuphold (posedge USERCLK, negedge CFGDSN[40], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[40]);
    $setuphold (posedge USERCLK, negedge CFGDSN[41], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[41]);
    $setuphold (posedge USERCLK, negedge CFGDSN[42], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[42]);
    $setuphold (posedge USERCLK, negedge CFGDSN[43], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[43]);
    $setuphold (posedge USERCLK, negedge CFGDSN[44], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[44]);
    $setuphold (posedge USERCLK, negedge CFGDSN[45], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[45]);
    $setuphold (posedge USERCLK, negedge CFGDSN[46], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[46]);
    $setuphold (posedge USERCLK, negedge CFGDSN[47], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[47]);
    $setuphold (posedge USERCLK, negedge CFGDSN[48], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[48]);
    $setuphold (posedge USERCLK, negedge CFGDSN[49], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[49]);
    $setuphold (posedge USERCLK, negedge CFGDSN[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[4]);
    $setuphold (posedge USERCLK, negedge CFGDSN[50], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[50]);
    $setuphold (posedge USERCLK, negedge CFGDSN[51], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[51]);
    $setuphold (posedge USERCLK, negedge CFGDSN[52], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[52]);
    $setuphold (posedge USERCLK, negedge CFGDSN[53], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[53]);
    $setuphold (posedge USERCLK, negedge CFGDSN[54], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[54]);
    $setuphold (posedge USERCLK, negedge CFGDSN[55], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[55]);
    $setuphold (posedge USERCLK, negedge CFGDSN[56], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[56]);
    $setuphold (posedge USERCLK, negedge CFGDSN[57], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[57]);
    $setuphold (posedge USERCLK, negedge CFGDSN[58], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[58]);
    $setuphold (posedge USERCLK, negedge CFGDSN[59], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[59]);
    $setuphold (posedge USERCLK, negedge CFGDSN[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[5]);
    $setuphold (posedge USERCLK, negedge CFGDSN[60], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[60]);
    $setuphold (posedge USERCLK, negedge CFGDSN[61], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[61]);
    $setuphold (posedge USERCLK, negedge CFGDSN[62], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[62]);
    $setuphold (posedge USERCLK, negedge CFGDSN[63], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[63]);
    $setuphold (posedge USERCLK, negedge CFGDSN[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[6]);
    $setuphold (posedge USERCLK, negedge CFGDSN[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[7]);
    $setuphold (posedge USERCLK, negedge CFGDSN[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[8]);
    $setuphold (posedge USERCLK, negedge CFGDSN[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[9]);
    $setuphold (posedge USERCLK, negedge CFGDSPORTNUMBER[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSPORTNUMBER_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGDSPORTNUMBER[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSPORTNUMBER_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGDSPORTNUMBER[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSPORTNUMBER_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGDSPORTNUMBER[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSPORTNUMBER_delay[3]);
    $setuphold (posedge USERCLK, negedge CFGDSPORTNUMBER[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSPORTNUMBER_delay[4]);
    $setuphold (posedge USERCLK, negedge CFGDSPORTNUMBER[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSPORTNUMBER_delay[5]);
    $setuphold (posedge USERCLK, negedge CFGDSPORTNUMBER[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSPORTNUMBER_delay[6]);
    $setuphold (posedge USERCLK, negedge CFGDSPORTNUMBER[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSPORTNUMBER_delay[7]);
    $setuphold (posedge USERCLK, negedge CFGERRCORIN, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGERRCORIN_delay);
    $setuphold (posedge USERCLK, negedge CFGERRUNCORIN, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGERRUNCORIN_delay);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATAVALID, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATAVALID_delay);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[10]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[11]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[12]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[13]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[14]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[15]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[16]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[17]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[18]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[19]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[20]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[21]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[22]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[23]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[24]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[25]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[26]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[27]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[28]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[29]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[30]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[31]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[3]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[4]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[5]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[6]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[7]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[8]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[9]);
    $setuphold (posedge USERCLK, negedge CFGFCSEL[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGFCSEL_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGFCSEL[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGFCSEL_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGFCSEL[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGFCSEL_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGFLRDONE[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGFLRDONE_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGFLRDONE[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGFLRDONE_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGHOTRESETIN, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGHOTRESETIN_delay);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTINT[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTINT_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTINT[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTINT_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTINT[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTINT_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTINT[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTINT_delay[3]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIATTR[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIATTR_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIATTR[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIATTR_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIATTR[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIATTR_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIFUNCTIONNUMBER[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIFUNCTIONNUMBER_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIFUNCTIONNUMBER[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIFUNCTIONNUMBER_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIFUNCTIONNUMBER[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIFUNCTIONNUMBER_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIFUNCTIONNUMBER[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIFUNCTIONNUMBER_delay[3]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[10]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[11]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[12]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[13]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[14]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[15]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[16]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[17]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[18]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[19]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[20]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[21]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[22]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[23]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[24]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[25]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[26]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[27]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[28]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[29]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[30]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[31]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[3]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[4]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[5]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[6]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[7]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[8]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[9]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUSDATAENABLE, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUSDATAENABLE_delay);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM_delay[3]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[10]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[11]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[12]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[13]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[14]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[15]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[16]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[17]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[18]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[19]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[20]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[21]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[22]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[23]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[24]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[25]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[26]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[27]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[28]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[29]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[30]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[31]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[3]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[4]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[5]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[6]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[7]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[8]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[9]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSISELECT[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSISELECT_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSISELECT[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSISELECT_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSISELECT[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSISELECT_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSISELECT[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSISELECT_delay[3]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHPRESENT, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSITPHPRESENT_delay);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHSTTAG[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSITPHSTTAG_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHSTTAG[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSITPHSTTAG_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHSTTAG[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSITPHSTTAG_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHSTTAG[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSITPHSTTAG_delay[3]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHSTTAG[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSITPHSTTAG_delay[4]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHSTTAG[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSITPHSTTAG_delay[5]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHSTTAG[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSITPHSTTAG_delay[6]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHSTTAG[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSITPHSTTAG_delay[7]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHSTTAG[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSITPHSTTAG_delay[8]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHTYPE[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSITPHTYPE_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHTYPE[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSITPHTYPE_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[10]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[11]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[12]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[13]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[14]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[15]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[16]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[17]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[18]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[19]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[20]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[21]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[22]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[23]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[24]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[25]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[26]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[27]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[28]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[29]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[30]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[31]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[32], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[32]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[33], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[33]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[34], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[34]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[35], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[35]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[36], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[36]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[37], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[37]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[38], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[38]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[39], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[39]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[3]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[40], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[40]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[41], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[41]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[42], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[42]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[43], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[43]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[44], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[44]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[45], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[45]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[46], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[46]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[47], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[47]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[48], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[48]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[49], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[49]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[4]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[50], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[50]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[51], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[51]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[52], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[52]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[53], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[53]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[54], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[54]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[55], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[55]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[56], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[56]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[57], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[57]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[58], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[58]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[59], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[59]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[5]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[60], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[60]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[61], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[61]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[62], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[62]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[63], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[63]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[6]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[7]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[8]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[9]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[10]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[11]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[12]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[13]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[14]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[15]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[16]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[17]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[18]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[19]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[20]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[21]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[22]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[23]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[24]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[25]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[26]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[27]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[28]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[29]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[30]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[31]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[3]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[4]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[5]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[6]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[7]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[8]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[9]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXINT, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXINT_delay);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTPENDING[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTPENDING_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTPENDING[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTPENDING_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGLINKTRAININGENABLE, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGLINKTRAININGENABLE_delay);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[10]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[11]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[12]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[13]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[14]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[15]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[16]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[17]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[18]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[3]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[4]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[5]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[6]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[7]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[8]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[9]);
    $setuphold (posedge USERCLK, negedge CFGMGMTBYTEENABLE[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTBYTEENABLE_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGMGMTBYTEENABLE[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTBYTEENABLE_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGMGMTBYTEENABLE[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTBYTEENABLE_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGMGMTBYTEENABLE[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTBYTEENABLE_delay[3]);
    $setuphold (posedge USERCLK, negedge CFGMGMTREAD, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTREAD_delay);
    $setuphold (posedge USERCLK, negedge CFGMGMTTYPE1CFGREGACCESS, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTTYPE1CFGREGACCESS_delay);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITE, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITE_delay);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[10]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[11]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[12]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[13]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[14]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[15]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[16]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[17]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[18]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[19]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[20]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[21]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[22]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[23]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[24]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[25]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[26]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[27]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[28]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[29]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[30]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[31]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[3]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[4]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[5]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[6]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[7]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[8]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[9]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMIT, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMIT_delay);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[10]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[11]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[12]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[13]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[14]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[15]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[16]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[17]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[18]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[19]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[20]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[21]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[22]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[23]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[24]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[25]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[26]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[27]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[28]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[29]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[30]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[31]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[3]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[4]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[5]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[6]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[7]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[8]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[9]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITTYPE[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITTYPE_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITTYPE[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITTYPE_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITTYPE[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITTYPE_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGPERFUNCSTATUSCONTROL[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGPERFUNCSTATUSCONTROL_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGPERFUNCSTATUSCONTROL[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGPERFUNCSTATUSCONTROL_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGPERFUNCSTATUSCONTROL[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGPERFUNCSTATUSCONTROL_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGPERFUNCTIONNUMBER[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGPERFUNCTIONNUMBER_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGPERFUNCTIONNUMBER[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGPERFUNCTIONNUMBER_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGPERFUNCTIONNUMBER[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGPERFUNCTIONNUMBER_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGPERFUNCTIONNUMBER[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGPERFUNCTIONNUMBER_delay[3]);
    $setuphold (posedge USERCLK, negedge CFGPERFUNCTIONOUTPUTREQUEST, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGPERFUNCTIONOUTPUTREQUEST_delay);
    $setuphold (posedge USERCLK, negedge CFGPOWERSTATECHANGEACK, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGPOWERSTATECHANGEACK_delay);
    $setuphold (posedge USERCLK, negedge CFGREQPMTRANSITIONL23READY, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGREQPMTRANSITIONL23READY_delay);
    $setuphold (posedge USERCLK, negedge CFGREVID[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGREVID_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGREVID[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGREVID_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGREVID[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGREVID_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGREVID[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGREVID_delay[3]);
    $setuphold (posedge USERCLK, negedge CFGREVID[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGREVID_delay[4]);
    $setuphold (posedge USERCLK, negedge CFGREVID[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGREVID_delay[5]);
    $setuphold (posedge USERCLK, negedge CFGREVID[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGREVID_delay[6]);
    $setuphold (posedge USERCLK, negedge CFGREVID[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGREVID_delay[7]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[10]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[11]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[12]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[13]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[14]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[15]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[3]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[4]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[5]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[6]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[7]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[8]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[9]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[10]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[11]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[12]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[13]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[14]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[15]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[3]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[4]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[5]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[6]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[7]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[8]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[9]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATAVALID, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATAVALID_delay);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[10]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[11]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[12]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[13]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[14]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[15]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[16]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[17]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[18]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[19]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[20]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[21]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[22]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[23]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[24]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[25]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[26]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[27]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[28]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[29]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[30]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[31]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[3]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[4]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[5]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[6]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[7]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[8]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[9]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[10]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[11]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[12]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[13]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[14]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[15]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[3]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[4]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[5]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[6]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[7]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[8]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[9]);
    $setuphold (posedge USERCLK, negedge CFGVFFLRDONE[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVFFLRDONE_delay[0]);
    $setuphold (posedge USERCLK, negedge CFGVFFLRDONE[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVFFLRDONE_delay[1]);
    $setuphold (posedge USERCLK, negedge CFGVFFLRDONE[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVFFLRDONE_delay[2]);
    $setuphold (posedge USERCLK, negedge CFGVFFLRDONE[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVFFLRDONE_delay[3]);
    $setuphold (posedge USERCLK, negedge CFGVFFLRDONE[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVFFLRDONE_delay[4]);
    $setuphold (posedge USERCLK, negedge CFGVFFLRDONE[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVFFLRDONE_delay[5]);
    $setuphold (posedge USERCLK, negedge CONFMCAPREQUESTBYCONF, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFMCAPREQUESTBYCONF_delay);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[0]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[10]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[11]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[12]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[13]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[14]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[15]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[16]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[17]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[18]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[19]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[1]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[20]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[21]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[22]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[23]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[24]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[25]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[26]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[27]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[28]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[29]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[2]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[30]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[31]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[3]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[4]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[5]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[6]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[7]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[8]);
    $setuphold (posedge USERCLK, negedge CONFREQDATA[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[9]);
    $setuphold (posedge USERCLK, negedge CONFREQREGNUM[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQREGNUM_delay[0]);
    $setuphold (posedge USERCLK, negedge CONFREQREGNUM[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQREGNUM_delay[1]);
    $setuphold (posedge USERCLK, negedge CONFREQREGNUM[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQREGNUM_delay[2]);
    $setuphold (posedge USERCLK, negedge CONFREQREGNUM[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQREGNUM_delay[3]);
    $setuphold (posedge USERCLK, negedge CONFREQTYPE[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQTYPE_delay[0]);
    $setuphold (posedge USERCLK, negedge CONFREQTYPE[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQTYPE_delay[1]);
    $setuphold (posedge USERCLK, negedge CONFREQVALID, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQVALID_delay);
    $setuphold (posedge USERCLK, negedge DBGCFGLOCALMGMTREGOVERRIDE, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, DBGCFGLOCALMGMTREGOVERRIDE_delay);
    $setuphold (posedge USERCLK, negedge DBGDATASEL[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, DBGDATASEL_delay[0]);
    $setuphold (posedge USERCLK, negedge DBGDATASEL[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, DBGDATASEL_delay[1]);
    $setuphold (posedge USERCLK, negedge DBGDATASEL[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, DBGDATASEL_delay[2]);
    $setuphold (posedge USERCLK, negedge DBGDATASEL[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, DBGDATASEL_delay[3]);
    $setuphold (posedge USERCLK, negedge LL2LMSAXISTXTUSER[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[0]);
    $setuphold (posedge USERCLK, negedge LL2LMSAXISTXTUSER[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[10]);
    $setuphold (posedge USERCLK, negedge LL2LMSAXISTXTUSER[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[11]);
    $setuphold (posedge USERCLK, negedge LL2LMSAXISTXTUSER[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[12]);
    $setuphold (posedge USERCLK, negedge LL2LMSAXISTXTUSER[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[13]);
    $setuphold (posedge USERCLK, negedge LL2LMSAXISTXTUSER[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[1]);
    $setuphold (posedge USERCLK, negedge LL2LMSAXISTXTUSER[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[2]);
    $setuphold (posedge USERCLK, negedge LL2LMSAXISTXTUSER[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[3]);
    $setuphold (posedge USERCLK, negedge LL2LMSAXISTXTUSER[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[4]);
    $setuphold (posedge USERCLK, negedge LL2LMSAXISTXTUSER[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[5]);
    $setuphold (posedge USERCLK, negedge LL2LMSAXISTXTUSER[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[6]);
    $setuphold (posedge USERCLK, negedge LL2LMSAXISTXTUSER[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[7]);
    $setuphold (posedge USERCLK, negedge LL2LMSAXISTXTUSER[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[8]);
    $setuphold (posedge USERCLK, negedge LL2LMSAXISTXTUSER[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[9]);
    $setuphold (posedge USERCLK, negedge LL2LMSAXISTXTVALID, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTVALID_delay);
    $setuphold (posedge USERCLK, negedge LL2LMTXTLPID0[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMTXTLPID0_delay[0]);
    $setuphold (posedge USERCLK, negedge LL2LMTXTLPID0[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMTXTLPID0_delay[1]);
    $setuphold (posedge USERCLK, negedge LL2LMTXTLPID0[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMTXTLPID0_delay[2]);
    $setuphold (posedge USERCLK, negedge LL2LMTXTLPID0[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMTXTLPID0_delay[3]);
    $setuphold (posedge USERCLK, negedge LL2LMTXTLPID1[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMTXTLPID1_delay[0]);
    $setuphold (posedge USERCLK, negedge LL2LMTXTLPID1[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMTXTLPID1_delay[1]);
    $setuphold (posedge USERCLK, negedge LL2LMTXTLPID1[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMTXTLPID1_delay[2]);
    $setuphold (posedge USERCLK, negedge LL2LMTXTLPID1[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMTXTLPID1_delay[3]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[0]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[10]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[11]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[12]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[13]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[14]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[15]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[16]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[17]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[18]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[19]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[1]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[20]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[21]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[2]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[3]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[4]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[5]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[6]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[7]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[8]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[9]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[0]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[10]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[11]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[12]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[13]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[14]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[15]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[16]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[17]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[18]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[19]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[1]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[20]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[21]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[2]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[3]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[4]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[5]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[6]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[7]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[8]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[9]);
    $setuphold (posedge USERCLK, negedge PCIECQNPREQ, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, PCIECQNPREQ_delay);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[0]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[100], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[100]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[101], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[101]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[102], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[102]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[103], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[103]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[104], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[104]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[105], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[105]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[106], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[106]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[107], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[107]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[108], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[108]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[109], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[109]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[10]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[110], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[110]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[111], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[111]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[112], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[112]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[113], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[113]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[114], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[114]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[115], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[115]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[116], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[116]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[117], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[117]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[118], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[118]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[119], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[119]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[11]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[120], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[120]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[121], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[121]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[122], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[122]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[123], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[123]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[124], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[124]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[125], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[125]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[126], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[126]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[127], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[127]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[128], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[128]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[129], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[129]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[12]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[130], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[130]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[131], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[131]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[132], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[132]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[133], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[133]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[134], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[134]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[135], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[135]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[136], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[136]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[137], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[137]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[138], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[138]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[139], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[139]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[13]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[140], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[140]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[141], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[141]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[142], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[142]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[143], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[143]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[144], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[144]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[145], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[145]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[146], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[146]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[147], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[147]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[148], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[148]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[149], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[149]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[14]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[150], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[150]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[151], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[151]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[152], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[152]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[153], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[153]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[154], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[154]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[155], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[155]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[156], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[156]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[157], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[157]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[158], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[158]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[159], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[159]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[15]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[160], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[160]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[161], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[161]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[162], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[162]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[163], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[163]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[164], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[164]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[165], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[165]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[166], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[166]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[167], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[167]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[168], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[168]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[169], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[169]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[16]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[170], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[170]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[171], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[171]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[172], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[172]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[173], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[173]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[174], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[174]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[175], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[175]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[176], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[176]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[177], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[177]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[178], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[178]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[179], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[179]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[17]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[180], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[180]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[181], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[181]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[182], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[182]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[183], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[183]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[184], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[184]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[185], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[185]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[186], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[186]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[187], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[187]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[188], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[188]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[189], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[189]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[18]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[190], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[190]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[191], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[191]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[192], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[192]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[193], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[193]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[194], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[194]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[195], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[195]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[196], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[196]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[197], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[197]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[198], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[198]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[199], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[199]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[19]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[1]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[200], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[200]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[201], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[201]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[202], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[202]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[203], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[203]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[204], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[204]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[205], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[205]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[206], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[206]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[207], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[207]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[208], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[208]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[209], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[209]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[20]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[210], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[210]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[211], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[211]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[212], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[212]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[213], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[213]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[214], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[214]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[215], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[215]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[216], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[216]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[217], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[217]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[218], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[218]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[219], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[219]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[21]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[220], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[220]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[221], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[221]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[222], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[222]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[223], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[223]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[224], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[224]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[225], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[225]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[226], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[226]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[227], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[227]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[228], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[228]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[229], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[229]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[22]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[230], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[230]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[231], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[231]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[232], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[232]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[233], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[233]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[234], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[234]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[235], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[235]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[236], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[236]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[237], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[237]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[238], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[238]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[239], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[239]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[23]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[240], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[240]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[241], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[241]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[242], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[242]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[243], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[243]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[244], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[244]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[245], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[245]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[246], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[246]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[247], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[247]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[248], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[248]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[249], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[249]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[24]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[250], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[250]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[251], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[251]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[252], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[252]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[253], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[253]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[254], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[254]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[255], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[255]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[25]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[26]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[27]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[28]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[29]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[2]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[30]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[31]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[32], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[32]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[33], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[33]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[34], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[34]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[35], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[35]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[36], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[36]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[37], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[37]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[38], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[38]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[39], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[39]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[3]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[40], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[40]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[41], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[41]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[42], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[42]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[43], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[43]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[44], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[44]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[45], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[45]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[46], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[46]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[47], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[47]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[48], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[48]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[49], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[49]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[4]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[50], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[50]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[51], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[51]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[52], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[52]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[53], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[53]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[54], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[54]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[55], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[55]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[56], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[56]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[57], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[57]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[58], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[58]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[59], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[59]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[5]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[60], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[60]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[61], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[61]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[62], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[62]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[63], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[63]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[64], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[64]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[65], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[65]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[66], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[66]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[67], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[67]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[68], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[68]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[69], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[69]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[6]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[70], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[70]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[71], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[71]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[72], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[72]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[73], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[73]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[74], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[74]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[75], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[75]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[76], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[76]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[77], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[77]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[78], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[78]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[79], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[79]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[7]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[80], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[80]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[81], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[81]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[82], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[82]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[83], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[83]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[84], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[84]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[85], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[85]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[86], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[86]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[87], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[87]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[88], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[88]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[89], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[89]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[8]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[90], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[90]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[91], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[91]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[92], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[92]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[93], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[93]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[94], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[94]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[95], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[95]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[96], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[96]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[97], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[97]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[98], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[98]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[99], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[99]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[9]);
    $setuphold (posedge USERCLK, negedge SAXISCCTKEEP[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTKEEP_delay[0]);
    $setuphold (posedge USERCLK, negedge SAXISCCTKEEP[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTKEEP_delay[1]);
    $setuphold (posedge USERCLK, negedge SAXISCCTKEEP[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTKEEP_delay[2]);
    $setuphold (posedge USERCLK, negedge SAXISCCTKEEP[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTKEEP_delay[3]);
    $setuphold (posedge USERCLK, negedge SAXISCCTKEEP[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTKEEP_delay[4]);
    $setuphold (posedge USERCLK, negedge SAXISCCTKEEP[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTKEEP_delay[5]);
    $setuphold (posedge USERCLK, negedge SAXISCCTKEEP[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTKEEP_delay[6]);
    $setuphold (posedge USERCLK, negedge SAXISCCTKEEP[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTKEEP_delay[7]);
    $setuphold (posedge USERCLK, negedge SAXISCCTLAST, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTLAST_delay);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[0]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[10]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[11]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[12]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[13]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[14]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[15]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[16]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[17]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[18]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[19]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[1]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[20]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[21]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[22]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[23]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[24]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[25]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[26]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[27]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[28]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[29]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[2]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[30]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[31]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[32], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[32]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[3]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[4]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[5]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[6]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[7]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[8]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[9]);
    $setuphold (posedge USERCLK, negedge SAXISCCTVALID, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTVALID_delay);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[0]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[100], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[100]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[101], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[101]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[102], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[102]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[103], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[103]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[104], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[104]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[105], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[105]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[106], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[106]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[107], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[107]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[108], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[108]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[109], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[109]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[10]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[110], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[110]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[111], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[111]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[112], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[112]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[113], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[113]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[114], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[114]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[115], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[115]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[116], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[116]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[117], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[117]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[118], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[118]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[119], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[119]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[11]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[120], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[120]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[121], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[121]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[122], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[122]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[123], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[123]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[124], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[124]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[125], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[125]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[126], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[126]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[127], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[127]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[128], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[128]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[129], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[129]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[12]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[130], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[130]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[131], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[131]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[132], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[132]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[133], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[133]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[134], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[134]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[135], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[135]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[136], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[136]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[137], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[137]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[138], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[138]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[139], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[139]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[13]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[140], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[140]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[141], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[141]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[142], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[142]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[143], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[143]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[144], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[144]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[145], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[145]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[146], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[146]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[147], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[147]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[148], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[148]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[149], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[149]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[14]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[150], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[150]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[151], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[151]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[152], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[152]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[153], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[153]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[154], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[154]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[155], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[155]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[156], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[156]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[157], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[157]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[158], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[158]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[159], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[159]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[15]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[160], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[160]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[161], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[161]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[162], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[162]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[163], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[163]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[164], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[164]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[165], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[165]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[166], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[166]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[167], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[167]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[168], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[168]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[169], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[169]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[16]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[170], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[170]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[171], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[171]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[172], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[172]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[173], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[173]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[174], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[174]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[175], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[175]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[176], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[176]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[177], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[177]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[178], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[178]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[179], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[179]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[17]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[180], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[180]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[181], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[181]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[182], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[182]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[183], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[183]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[184], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[184]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[185], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[185]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[186], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[186]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[187], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[187]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[188], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[188]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[189], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[189]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[18]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[190], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[190]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[191], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[191]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[192], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[192]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[193], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[193]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[194], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[194]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[195], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[195]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[196], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[196]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[197], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[197]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[198], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[198]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[199], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[199]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[19]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[1]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[200], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[200]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[201], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[201]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[202], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[202]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[203], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[203]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[204], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[204]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[205], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[205]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[206], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[206]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[207], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[207]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[208], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[208]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[209], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[209]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[20]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[210], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[210]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[211], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[211]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[212], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[212]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[213], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[213]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[214], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[214]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[215], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[215]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[216], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[216]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[217], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[217]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[218], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[218]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[219], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[219]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[21]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[220], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[220]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[221], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[221]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[222], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[222]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[223], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[223]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[224], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[224]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[225], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[225]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[226], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[226]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[227], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[227]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[228], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[228]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[229], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[229]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[22]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[230], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[230]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[231], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[231]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[232], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[232]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[233], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[233]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[234], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[234]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[235], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[235]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[236], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[236]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[237], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[237]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[238], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[238]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[239], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[239]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[23]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[240], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[240]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[241], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[241]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[242], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[242]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[243], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[243]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[244], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[244]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[245], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[245]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[246], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[246]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[247], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[247]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[248], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[248]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[249], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[249]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[24]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[250], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[250]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[251], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[251]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[252], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[252]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[253], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[253]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[254], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[254]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[255], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[255]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[25]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[26]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[27]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[28]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[29]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[2]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[30]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[31]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[32], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[32]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[33], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[33]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[34], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[34]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[35], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[35]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[36], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[36]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[37], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[37]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[38], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[38]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[39], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[39]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[3]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[40], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[40]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[41], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[41]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[42], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[42]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[43], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[43]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[44], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[44]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[45], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[45]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[46], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[46]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[47], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[47]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[48], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[48]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[49], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[49]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[4]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[50], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[50]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[51], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[51]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[52], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[52]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[53], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[53]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[54], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[54]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[55], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[55]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[56], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[56]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[57], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[57]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[58], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[58]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[59], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[59]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[5]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[60], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[60]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[61], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[61]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[62], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[62]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[63], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[63]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[64], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[64]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[65], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[65]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[66], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[66]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[67], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[67]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[68], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[68]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[69], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[69]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[6]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[70], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[70]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[71], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[71]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[72], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[72]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[73], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[73]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[74], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[74]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[75], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[75]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[76], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[76]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[77], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[77]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[78], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[78]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[79], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[79]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[7]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[80], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[80]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[81], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[81]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[82], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[82]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[83], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[83]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[84], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[84]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[85], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[85]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[86], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[86]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[87], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[87]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[88], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[88]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[89], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[89]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[8]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[90], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[90]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[91], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[91]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[92], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[92]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[93], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[93]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[94], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[94]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[95], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[95]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[96], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[96]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[97], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[97]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[98], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[98]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[99], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[99]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[9]);
    $setuphold (posedge USERCLK, negedge SAXISRQTKEEP[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTKEEP_delay[0]);
    $setuphold (posedge USERCLK, negedge SAXISRQTKEEP[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTKEEP_delay[1]);
    $setuphold (posedge USERCLK, negedge SAXISRQTKEEP[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTKEEP_delay[2]);
    $setuphold (posedge USERCLK, negedge SAXISRQTKEEP[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTKEEP_delay[3]);
    $setuphold (posedge USERCLK, negedge SAXISRQTKEEP[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTKEEP_delay[4]);
    $setuphold (posedge USERCLK, negedge SAXISRQTKEEP[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTKEEP_delay[5]);
    $setuphold (posedge USERCLK, negedge SAXISRQTKEEP[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTKEEP_delay[6]);
    $setuphold (posedge USERCLK, negedge SAXISRQTKEEP[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTKEEP_delay[7]);
    $setuphold (posedge USERCLK, negedge SAXISRQTLAST, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTLAST_delay);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[0]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[10]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[11]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[12]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[13]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[14]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[15]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[16]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[17]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[18]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[19]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[1]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[20]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[21]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[22]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[23]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[24]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[25]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[26]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[27]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[28]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[29]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[2]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[30]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[31]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[32], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[32]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[33], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[33]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[34], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[34]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[35], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[35]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[36], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[36]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[37], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[37]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[38], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[38]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[39], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[39]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[3]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[40], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[40]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[41], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[41]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[42], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[42]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[43], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[43]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[44], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[44]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[45], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[45]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[46], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[46]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[47], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[47]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[48], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[48]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[49], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[49]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[4]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[50], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[50]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[51], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[51]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[52], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[52]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[53], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[53]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[54], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[54]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[55], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[55]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[56], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[56]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[57], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[57]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[58], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[58]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[59], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[59]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[5]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[6]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[7]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[8]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[9]);
    $setuphold (posedge USERCLK, negedge SAXISRQTVALID, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTVALID_delay);
    $setuphold (posedge USERCLK, posedge CFGCONFIGSPACEENABLE, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGCONFIGSPACEENABLE_delay);
    $setuphold (posedge USERCLK, posedge CFGDEVID[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[10]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[11]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[12]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[13]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[14]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[15]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[3]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[4]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[5]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[6]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[7]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[8]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDEVID_delay[9]);
    $setuphold (posedge USERCLK, posedge CFGDSBUSNUMBER[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSBUSNUMBER_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGDSBUSNUMBER[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSBUSNUMBER_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGDSBUSNUMBER[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSBUSNUMBER_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGDSBUSNUMBER[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSBUSNUMBER_delay[3]);
    $setuphold (posedge USERCLK, posedge CFGDSBUSNUMBER[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSBUSNUMBER_delay[4]);
    $setuphold (posedge USERCLK, posedge CFGDSBUSNUMBER[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSBUSNUMBER_delay[5]);
    $setuphold (posedge USERCLK, posedge CFGDSBUSNUMBER[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSBUSNUMBER_delay[6]);
    $setuphold (posedge USERCLK, posedge CFGDSBUSNUMBER[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSBUSNUMBER_delay[7]);
    $setuphold (posedge USERCLK, posedge CFGDSDEVICENUMBER[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSDEVICENUMBER_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGDSDEVICENUMBER[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSDEVICENUMBER_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGDSDEVICENUMBER[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSDEVICENUMBER_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGDSDEVICENUMBER[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSDEVICENUMBER_delay[3]);
    $setuphold (posedge USERCLK, posedge CFGDSDEVICENUMBER[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSDEVICENUMBER_delay[4]);
    $setuphold (posedge USERCLK, posedge CFGDSFUNCTIONNUMBER[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSFUNCTIONNUMBER_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGDSFUNCTIONNUMBER[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSFUNCTIONNUMBER_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGDSFUNCTIONNUMBER[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSFUNCTIONNUMBER_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGDSN[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGDSN[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[10]);
    $setuphold (posedge USERCLK, posedge CFGDSN[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[11]);
    $setuphold (posedge USERCLK, posedge CFGDSN[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[12]);
    $setuphold (posedge USERCLK, posedge CFGDSN[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[13]);
    $setuphold (posedge USERCLK, posedge CFGDSN[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[14]);
    $setuphold (posedge USERCLK, posedge CFGDSN[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[15]);
    $setuphold (posedge USERCLK, posedge CFGDSN[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[16]);
    $setuphold (posedge USERCLK, posedge CFGDSN[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[17]);
    $setuphold (posedge USERCLK, posedge CFGDSN[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[18]);
    $setuphold (posedge USERCLK, posedge CFGDSN[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[19]);
    $setuphold (posedge USERCLK, posedge CFGDSN[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGDSN[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[20]);
    $setuphold (posedge USERCLK, posedge CFGDSN[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[21]);
    $setuphold (posedge USERCLK, posedge CFGDSN[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[22]);
    $setuphold (posedge USERCLK, posedge CFGDSN[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[23]);
    $setuphold (posedge USERCLK, posedge CFGDSN[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[24]);
    $setuphold (posedge USERCLK, posedge CFGDSN[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[25]);
    $setuphold (posedge USERCLK, posedge CFGDSN[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[26]);
    $setuphold (posedge USERCLK, posedge CFGDSN[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[27]);
    $setuphold (posedge USERCLK, posedge CFGDSN[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[28]);
    $setuphold (posedge USERCLK, posedge CFGDSN[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[29]);
    $setuphold (posedge USERCLK, posedge CFGDSN[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGDSN[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[30]);
    $setuphold (posedge USERCLK, posedge CFGDSN[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[31]);
    $setuphold (posedge USERCLK, posedge CFGDSN[32], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[32]);
    $setuphold (posedge USERCLK, posedge CFGDSN[33], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[33]);
    $setuphold (posedge USERCLK, posedge CFGDSN[34], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[34]);
    $setuphold (posedge USERCLK, posedge CFGDSN[35], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[35]);
    $setuphold (posedge USERCLK, posedge CFGDSN[36], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[36]);
    $setuphold (posedge USERCLK, posedge CFGDSN[37], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[37]);
    $setuphold (posedge USERCLK, posedge CFGDSN[38], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[38]);
    $setuphold (posedge USERCLK, posedge CFGDSN[39], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[39]);
    $setuphold (posedge USERCLK, posedge CFGDSN[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[3]);
    $setuphold (posedge USERCLK, posedge CFGDSN[40], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[40]);
    $setuphold (posedge USERCLK, posedge CFGDSN[41], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[41]);
    $setuphold (posedge USERCLK, posedge CFGDSN[42], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[42]);
    $setuphold (posedge USERCLK, posedge CFGDSN[43], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[43]);
    $setuphold (posedge USERCLK, posedge CFGDSN[44], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[44]);
    $setuphold (posedge USERCLK, posedge CFGDSN[45], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[45]);
    $setuphold (posedge USERCLK, posedge CFGDSN[46], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[46]);
    $setuphold (posedge USERCLK, posedge CFGDSN[47], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[47]);
    $setuphold (posedge USERCLK, posedge CFGDSN[48], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[48]);
    $setuphold (posedge USERCLK, posedge CFGDSN[49], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[49]);
    $setuphold (posedge USERCLK, posedge CFGDSN[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[4]);
    $setuphold (posedge USERCLK, posedge CFGDSN[50], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[50]);
    $setuphold (posedge USERCLK, posedge CFGDSN[51], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[51]);
    $setuphold (posedge USERCLK, posedge CFGDSN[52], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[52]);
    $setuphold (posedge USERCLK, posedge CFGDSN[53], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[53]);
    $setuphold (posedge USERCLK, posedge CFGDSN[54], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[54]);
    $setuphold (posedge USERCLK, posedge CFGDSN[55], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[55]);
    $setuphold (posedge USERCLK, posedge CFGDSN[56], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[56]);
    $setuphold (posedge USERCLK, posedge CFGDSN[57], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[57]);
    $setuphold (posedge USERCLK, posedge CFGDSN[58], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[58]);
    $setuphold (posedge USERCLK, posedge CFGDSN[59], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[59]);
    $setuphold (posedge USERCLK, posedge CFGDSN[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[5]);
    $setuphold (posedge USERCLK, posedge CFGDSN[60], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[60]);
    $setuphold (posedge USERCLK, posedge CFGDSN[61], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[61]);
    $setuphold (posedge USERCLK, posedge CFGDSN[62], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[62]);
    $setuphold (posedge USERCLK, posedge CFGDSN[63], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[63]);
    $setuphold (posedge USERCLK, posedge CFGDSN[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[6]);
    $setuphold (posedge USERCLK, posedge CFGDSN[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[7]);
    $setuphold (posedge USERCLK, posedge CFGDSN[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[8]);
    $setuphold (posedge USERCLK, posedge CFGDSN[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSN_delay[9]);
    $setuphold (posedge USERCLK, posedge CFGDSPORTNUMBER[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSPORTNUMBER_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGDSPORTNUMBER[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSPORTNUMBER_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGDSPORTNUMBER[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSPORTNUMBER_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGDSPORTNUMBER[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSPORTNUMBER_delay[3]);
    $setuphold (posedge USERCLK, posedge CFGDSPORTNUMBER[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSPORTNUMBER_delay[4]);
    $setuphold (posedge USERCLK, posedge CFGDSPORTNUMBER[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSPORTNUMBER_delay[5]);
    $setuphold (posedge USERCLK, posedge CFGDSPORTNUMBER[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSPORTNUMBER_delay[6]);
    $setuphold (posedge USERCLK, posedge CFGDSPORTNUMBER[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGDSPORTNUMBER_delay[7]);
    $setuphold (posedge USERCLK, posedge CFGERRCORIN, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGERRCORIN_delay);
    $setuphold (posedge USERCLK, posedge CFGERRUNCORIN, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGERRUNCORIN_delay);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATAVALID, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATAVALID_delay);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[10]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[11]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[12]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[13]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[14]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[15]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[16]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[17]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[18]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[19]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[20]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[21]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[22]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[23]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[24]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[25]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[26]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[27]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[28]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[29]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[30]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[31]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[3]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[4]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[5]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[6]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[7]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[8]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGEXTREADDATA_delay[9]);
    $setuphold (posedge USERCLK, posedge CFGFCSEL[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGFCSEL_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGFCSEL[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGFCSEL_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGFCSEL[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGFCSEL_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGFLRDONE[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGFLRDONE_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGFLRDONE[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGFLRDONE_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGHOTRESETIN, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGHOTRESETIN_delay);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTINT[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTINT_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTINT[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTINT_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTINT[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTINT_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTINT[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTINT_delay[3]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIATTR[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIATTR_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIATTR[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIATTR_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIATTR[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIATTR_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIFUNCTIONNUMBER[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIFUNCTIONNUMBER_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIFUNCTIONNUMBER[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIFUNCTIONNUMBER_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIFUNCTIONNUMBER[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIFUNCTIONNUMBER_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIFUNCTIONNUMBER[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIFUNCTIONNUMBER_delay[3]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[10]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[11]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[12]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[13]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[14]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[15]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[16]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[17]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[18]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[19]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[20]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[21]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[22]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[23]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[24]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[25]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[26]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[27]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[28]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[29]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[30]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[31]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[3]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[4]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[5]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[6]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[7]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[8]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIINT_delay[9]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUSDATAENABLE, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUSDATAENABLE_delay);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUSFUNCTIONNUM_delay[3]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[10]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[11]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[12]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[13]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[14]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[15]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[16]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[17]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[18]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[19]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[20]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[21]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[22]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[23]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[24]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[25]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[26]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[27]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[28]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[29]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[30]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[31]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[3]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[4]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[5]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[6]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[7]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[8]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIPENDINGSTATUS_delay[9]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSISELECT[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSISELECT_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSISELECT[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSISELECT_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSISELECT[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSISELECT_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSISELECT[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSISELECT_delay[3]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHPRESENT, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSITPHPRESENT_delay);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHSTTAG[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSITPHSTTAG_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHSTTAG[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSITPHSTTAG_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHSTTAG[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSITPHSTTAG_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHSTTAG[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSITPHSTTAG_delay[3]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHSTTAG[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSITPHSTTAG_delay[4]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHSTTAG[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSITPHSTTAG_delay[5]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHSTTAG[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSITPHSTTAG_delay[6]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHSTTAG[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSITPHSTTAG_delay[7]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHSTTAG[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSITPHSTTAG_delay[8]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHTYPE[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSITPHTYPE_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHTYPE[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSITPHTYPE_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[10]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[11]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[12]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[13]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[14]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[15]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[16]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[17]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[18]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[19]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[20]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[21]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[22]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[23]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[24]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[25]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[26]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[27]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[28]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[29]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[30]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[31]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[32], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[32]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[33], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[33]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[34], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[34]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[35], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[35]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[36], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[36]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[37], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[37]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[38], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[38]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[39], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[39]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[3]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[40], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[40]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[41], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[41]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[42], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[42]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[43], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[43]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[44], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[44]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[45], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[45]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[46], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[46]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[47], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[47]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[48], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[48]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[49], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[49]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[4]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[50], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[50]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[51], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[51]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[52], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[52]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[53], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[53]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[54], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[54]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[55], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[55]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[56], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[56]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[57], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[57]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[58], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[58]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[59], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[59]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[5]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[60], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[60]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[61], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[61]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[62], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[62]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[63], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[63]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[6]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[7]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[8]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXADDRESS_delay[9]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[10]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[11]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[12]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[13]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[14]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[15]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[16]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[17]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[18]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[19]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[20]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[21]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[22]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[23]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[24]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[25]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[26]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[27]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[28]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[29]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[30]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[31]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[3]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[4]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[5]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[6]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[7]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[8]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXDATA_delay[9]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXINT, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTMSIXINT_delay);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTPENDING[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTPENDING_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTPENDING[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGINTERRUPTPENDING_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGLINKTRAININGENABLE, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGLINKTRAININGENABLE_delay);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[10]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[11]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[12]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[13]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[14]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[15]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[16]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[17]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[18]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[3]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[4]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[5]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[6]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[7]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[8]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTADDR_delay[9]);
    $setuphold (posedge USERCLK, posedge CFGMGMTBYTEENABLE[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTBYTEENABLE_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGMGMTBYTEENABLE[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTBYTEENABLE_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGMGMTBYTEENABLE[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTBYTEENABLE_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGMGMTBYTEENABLE[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTBYTEENABLE_delay[3]);
    $setuphold (posedge USERCLK, posedge CFGMGMTREAD, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTREAD_delay);
    $setuphold (posedge USERCLK, posedge CFGMGMTTYPE1CFGREGACCESS, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTTYPE1CFGREGACCESS_delay);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITE, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITE_delay);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[10]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[11]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[12]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[13]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[14]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[15]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[16]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[17]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[18]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[19]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[20]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[21]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[22]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[23]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[24]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[25]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[26]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[27]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[28]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[29]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[30]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[31]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[3]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[4]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[5]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[6]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[7]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[8]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMGMTWRITEDATA_delay[9]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMIT, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMIT_delay);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[10]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[11]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[12]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[13]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[14]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[15]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[16]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[17]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[18]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[19]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[20]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[21]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[22]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[23]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[24]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[25]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[26]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[27]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[28]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[29]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[30]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[31]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[3]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[4]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[5]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[6]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[7]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[8]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITDATA_delay[9]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITTYPE[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITTYPE_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITTYPE[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITTYPE_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITTYPE[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGMSGTRANSMITTYPE_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGPERFUNCSTATUSCONTROL[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGPERFUNCSTATUSCONTROL_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGPERFUNCSTATUSCONTROL[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGPERFUNCSTATUSCONTROL_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGPERFUNCSTATUSCONTROL[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGPERFUNCSTATUSCONTROL_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGPERFUNCTIONNUMBER[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGPERFUNCTIONNUMBER_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGPERFUNCTIONNUMBER[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGPERFUNCTIONNUMBER_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGPERFUNCTIONNUMBER[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGPERFUNCTIONNUMBER_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGPERFUNCTIONNUMBER[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGPERFUNCTIONNUMBER_delay[3]);
    $setuphold (posedge USERCLK, posedge CFGPERFUNCTIONOUTPUTREQUEST, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGPERFUNCTIONOUTPUTREQUEST_delay);
    $setuphold (posedge USERCLK, posedge CFGPOWERSTATECHANGEACK, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGPOWERSTATECHANGEACK_delay);
    $setuphold (posedge USERCLK, posedge CFGREQPMTRANSITIONL23READY, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGREQPMTRANSITIONL23READY_delay);
    $setuphold (posedge USERCLK, posedge CFGREVID[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGREVID_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGREVID[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGREVID_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGREVID[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGREVID_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGREVID[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGREVID_delay[3]);
    $setuphold (posedge USERCLK, posedge CFGREVID[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGREVID_delay[4]);
    $setuphold (posedge USERCLK, posedge CFGREVID[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGREVID_delay[5]);
    $setuphold (posedge USERCLK, posedge CFGREVID[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGREVID_delay[6]);
    $setuphold (posedge USERCLK, posedge CFGREVID[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGREVID_delay[7]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[10]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[11]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[12]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[13]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[14]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[15]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[3]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[4]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[5]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[6]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[7]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[8]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSID_delay[9]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[10]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[11]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[12]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[13]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[14]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[15]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[3]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[4]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[5]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[6]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[7]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[8]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGSUBSYSVENDID_delay[9]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATAVALID, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATAVALID_delay);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[10]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[11]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[12]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[13]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[14]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[15]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[16]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[17]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[18]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[19]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[20]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[21]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[22]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[23]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[24]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[25]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[26]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[27]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[28]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[29]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[30]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[31]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[3]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[4]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[5]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[6]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[7]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[8]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGTPHSTTREADDATA_delay[9]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[10]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[11]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[12]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[13]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[14]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[15]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[3]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[4]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[5]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[6]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[7]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[8]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVENDID_delay[9]);
    $setuphold (posedge USERCLK, posedge CFGVFFLRDONE[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVFFLRDONE_delay[0]);
    $setuphold (posedge USERCLK, posedge CFGVFFLRDONE[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVFFLRDONE_delay[1]);
    $setuphold (posedge USERCLK, posedge CFGVFFLRDONE[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVFFLRDONE_delay[2]);
    $setuphold (posedge USERCLK, posedge CFGVFFLRDONE[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVFFLRDONE_delay[3]);
    $setuphold (posedge USERCLK, posedge CFGVFFLRDONE[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVFFLRDONE_delay[4]);
    $setuphold (posedge USERCLK, posedge CFGVFFLRDONE[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CFGVFFLRDONE_delay[5]);
    $setuphold (posedge USERCLK, posedge CONFMCAPREQUESTBYCONF, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFMCAPREQUESTBYCONF_delay);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[0]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[10]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[11]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[12]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[13]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[14]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[15]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[16]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[17]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[18]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[19]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[1]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[20]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[21]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[22]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[23]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[24]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[25]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[26]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[27]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[28]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[29]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[2]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[30]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[31]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[3]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[4]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[5]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[6]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[7]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[8]);
    $setuphold (posedge USERCLK, posedge CONFREQDATA[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQDATA_delay[9]);
    $setuphold (posedge USERCLK, posedge CONFREQREGNUM[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQREGNUM_delay[0]);
    $setuphold (posedge USERCLK, posedge CONFREQREGNUM[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQREGNUM_delay[1]);
    $setuphold (posedge USERCLK, posedge CONFREQREGNUM[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQREGNUM_delay[2]);
    $setuphold (posedge USERCLK, posedge CONFREQREGNUM[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQREGNUM_delay[3]);
    $setuphold (posedge USERCLK, posedge CONFREQTYPE[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQTYPE_delay[0]);
    $setuphold (posedge USERCLK, posedge CONFREQTYPE[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQTYPE_delay[1]);
    $setuphold (posedge USERCLK, posedge CONFREQVALID, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, CONFREQVALID_delay);
    $setuphold (posedge USERCLK, posedge DBGCFGLOCALMGMTREGOVERRIDE, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, DBGCFGLOCALMGMTREGOVERRIDE_delay);
    $setuphold (posedge USERCLK, posedge DBGDATASEL[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, DBGDATASEL_delay[0]);
    $setuphold (posedge USERCLK, posedge DBGDATASEL[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, DBGDATASEL_delay[1]);
    $setuphold (posedge USERCLK, posedge DBGDATASEL[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, DBGDATASEL_delay[2]);
    $setuphold (posedge USERCLK, posedge DBGDATASEL[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, DBGDATASEL_delay[3]);
    $setuphold (posedge USERCLK, posedge LL2LMSAXISTXTUSER[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[0]);
    $setuphold (posedge USERCLK, posedge LL2LMSAXISTXTUSER[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[10]);
    $setuphold (posedge USERCLK, posedge LL2LMSAXISTXTUSER[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[11]);
    $setuphold (posedge USERCLK, posedge LL2LMSAXISTXTUSER[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[12]);
    $setuphold (posedge USERCLK, posedge LL2LMSAXISTXTUSER[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[13]);
    $setuphold (posedge USERCLK, posedge LL2LMSAXISTXTUSER[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[1]);
    $setuphold (posedge USERCLK, posedge LL2LMSAXISTXTUSER[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[2]);
    $setuphold (posedge USERCLK, posedge LL2LMSAXISTXTUSER[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[3]);
    $setuphold (posedge USERCLK, posedge LL2LMSAXISTXTUSER[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[4]);
    $setuphold (posedge USERCLK, posedge LL2LMSAXISTXTUSER[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[5]);
    $setuphold (posedge USERCLK, posedge LL2LMSAXISTXTUSER[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[6]);
    $setuphold (posedge USERCLK, posedge LL2LMSAXISTXTUSER[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[7]);
    $setuphold (posedge USERCLK, posedge LL2LMSAXISTXTUSER[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[8]);
    $setuphold (posedge USERCLK, posedge LL2LMSAXISTXTUSER[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTUSER_delay[9]);
    $setuphold (posedge USERCLK, posedge LL2LMSAXISTXTVALID, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMSAXISTXTVALID_delay);
    $setuphold (posedge USERCLK, posedge LL2LMTXTLPID0[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMTXTLPID0_delay[0]);
    $setuphold (posedge USERCLK, posedge LL2LMTXTLPID0[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMTXTLPID0_delay[1]);
    $setuphold (posedge USERCLK, posedge LL2LMTXTLPID0[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMTXTLPID0_delay[2]);
    $setuphold (posedge USERCLK, posedge LL2LMTXTLPID0[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMTXTLPID0_delay[3]);
    $setuphold (posedge USERCLK, posedge LL2LMTXTLPID1[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMTXTLPID1_delay[0]);
    $setuphold (posedge USERCLK, posedge LL2LMTXTLPID1[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMTXTLPID1_delay[1]);
    $setuphold (posedge USERCLK, posedge LL2LMTXTLPID1[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMTXTLPID1_delay[2]);
    $setuphold (posedge USERCLK, posedge LL2LMTXTLPID1[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, LL2LMTXTLPID1_delay[3]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[0]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[10]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[11]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[12]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[13]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[14]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[15]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[16]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[17]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[18]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[19]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[1]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[20]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[21]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[2]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[3]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[4]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[5]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[6]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[7]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[8]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISCQTREADY_delay[9]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[0]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[10]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[11]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[12]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[13]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[14]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[15]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[16]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[17]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[18]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[19]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[1]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[20]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[21]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[2]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[3]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[4]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[5]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[6]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[7]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[8]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, MAXISRCTREADY_delay[9]);
    $setuphold (posedge USERCLK, posedge PCIECQNPREQ, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, PCIECQNPREQ_delay);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[0]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[100], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[100]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[101], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[101]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[102], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[102]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[103], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[103]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[104], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[104]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[105], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[105]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[106], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[106]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[107], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[107]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[108], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[108]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[109], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[109]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[10]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[110], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[110]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[111], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[111]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[112], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[112]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[113], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[113]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[114], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[114]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[115], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[115]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[116], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[116]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[117], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[117]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[118], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[118]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[119], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[119]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[11]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[120], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[120]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[121], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[121]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[122], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[122]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[123], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[123]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[124], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[124]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[125], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[125]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[126], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[126]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[127], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[127]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[128], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[128]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[129], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[129]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[12]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[130], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[130]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[131], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[131]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[132], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[132]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[133], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[133]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[134], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[134]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[135], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[135]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[136], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[136]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[137], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[137]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[138], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[138]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[139], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[139]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[13]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[140], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[140]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[141], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[141]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[142], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[142]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[143], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[143]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[144], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[144]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[145], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[145]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[146], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[146]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[147], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[147]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[148], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[148]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[149], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[149]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[14]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[150], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[150]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[151], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[151]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[152], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[152]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[153], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[153]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[154], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[154]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[155], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[155]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[156], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[156]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[157], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[157]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[158], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[158]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[159], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[159]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[15]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[160], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[160]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[161], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[161]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[162], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[162]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[163], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[163]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[164], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[164]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[165], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[165]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[166], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[166]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[167], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[167]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[168], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[168]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[169], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[169]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[16]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[170], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[170]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[171], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[171]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[172], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[172]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[173], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[173]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[174], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[174]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[175], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[175]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[176], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[176]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[177], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[177]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[178], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[178]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[179], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[179]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[17]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[180], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[180]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[181], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[181]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[182], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[182]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[183], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[183]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[184], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[184]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[185], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[185]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[186], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[186]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[187], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[187]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[188], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[188]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[189], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[189]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[18]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[190], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[190]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[191], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[191]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[192], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[192]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[193], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[193]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[194], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[194]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[195], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[195]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[196], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[196]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[197], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[197]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[198], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[198]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[199], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[199]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[19]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[1]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[200], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[200]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[201], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[201]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[202], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[202]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[203], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[203]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[204], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[204]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[205], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[205]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[206], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[206]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[207], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[207]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[208], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[208]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[209], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[209]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[20]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[210], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[210]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[211], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[211]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[212], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[212]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[213], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[213]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[214], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[214]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[215], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[215]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[216], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[216]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[217], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[217]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[218], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[218]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[219], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[219]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[21]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[220], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[220]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[221], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[221]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[222], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[222]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[223], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[223]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[224], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[224]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[225], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[225]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[226], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[226]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[227], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[227]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[228], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[228]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[229], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[229]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[22]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[230], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[230]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[231], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[231]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[232], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[232]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[233], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[233]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[234], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[234]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[235], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[235]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[236], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[236]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[237], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[237]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[238], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[238]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[239], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[239]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[23]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[240], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[240]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[241], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[241]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[242], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[242]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[243], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[243]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[244], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[244]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[245], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[245]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[246], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[246]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[247], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[247]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[248], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[248]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[249], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[249]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[24]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[250], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[250]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[251], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[251]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[252], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[252]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[253], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[253]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[254], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[254]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[255], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[255]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[25]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[26]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[27]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[28]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[29]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[2]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[30]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[31]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[32], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[32]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[33], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[33]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[34], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[34]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[35], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[35]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[36], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[36]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[37], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[37]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[38], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[38]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[39], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[39]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[3]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[40], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[40]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[41], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[41]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[42], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[42]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[43], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[43]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[44], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[44]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[45], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[45]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[46], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[46]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[47], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[47]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[48], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[48]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[49], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[49]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[4]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[50], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[50]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[51], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[51]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[52], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[52]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[53], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[53]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[54], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[54]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[55], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[55]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[56], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[56]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[57], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[57]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[58], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[58]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[59], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[59]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[5]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[60], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[60]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[61], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[61]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[62], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[62]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[63], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[63]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[64], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[64]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[65], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[65]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[66], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[66]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[67], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[67]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[68], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[68]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[69], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[69]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[6]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[70], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[70]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[71], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[71]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[72], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[72]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[73], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[73]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[74], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[74]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[75], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[75]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[76], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[76]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[77], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[77]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[78], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[78]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[79], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[79]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[7]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[80], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[80]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[81], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[81]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[82], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[82]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[83], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[83]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[84], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[84]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[85], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[85]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[86], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[86]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[87], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[87]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[88], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[88]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[89], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[89]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[8]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[90], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[90]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[91], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[91]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[92], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[92]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[93], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[93]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[94], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[94]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[95], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[95]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[96], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[96]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[97], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[97]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[98], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[98]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[99], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[99]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTDATA_delay[9]);
    $setuphold (posedge USERCLK, posedge SAXISCCTKEEP[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTKEEP_delay[0]);
    $setuphold (posedge USERCLK, posedge SAXISCCTKEEP[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTKEEP_delay[1]);
    $setuphold (posedge USERCLK, posedge SAXISCCTKEEP[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTKEEP_delay[2]);
    $setuphold (posedge USERCLK, posedge SAXISCCTKEEP[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTKEEP_delay[3]);
    $setuphold (posedge USERCLK, posedge SAXISCCTKEEP[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTKEEP_delay[4]);
    $setuphold (posedge USERCLK, posedge SAXISCCTKEEP[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTKEEP_delay[5]);
    $setuphold (posedge USERCLK, posedge SAXISCCTKEEP[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTKEEP_delay[6]);
    $setuphold (posedge USERCLK, posedge SAXISCCTKEEP[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTKEEP_delay[7]);
    $setuphold (posedge USERCLK, posedge SAXISCCTLAST, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTLAST_delay);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[0]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[10]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[11]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[12]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[13]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[14]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[15]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[16]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[17]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[18]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[19]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[1]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[20]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[21]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[22]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[23]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[24]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[25]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[26]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[27]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[28]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[29]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[2]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[30]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[31]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[32], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[32]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[3]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[4]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[5]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[6]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[7]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[8]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTUSER_delay[9]);
    $setuphold (posedge USERCLK, posedge SAXISCCTVALID, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISCCTVALID_delay);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[0]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[100], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[100]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[101], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[101]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[102], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[102]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[103], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[103]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[104], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[104]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[105], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[105]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[106], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[106]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[107], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[107]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[108], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[108]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[109], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[109]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[10]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[110], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[110]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[111], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[111]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[112], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[112]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[113], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[113]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[114], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[114]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[115], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[115]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[116], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[116]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[117], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[117]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[118], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[118]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[119], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[119]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[11]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[120], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[120]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[121], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[121]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[122], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[122]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[123], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[123]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[124], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[124]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[125], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[125]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[126], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[126]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[127], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[127]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[128], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[128]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[129], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[129]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[12]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[130], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[130]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[131], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[131]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[132], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[132]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[133], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[133]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[134], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[134]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[135], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[135]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[136], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[136]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[137], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[137]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[138], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[138]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[139], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[139]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[13]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[140], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[140]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[141], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[141]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[142], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[142]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[143], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[143]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[144], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[144]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[145], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[145]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[146], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[146]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[147], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[147]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[148], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[148]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[149], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[149]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[14]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[150], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[150]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[151], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[151]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[152], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[152]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[153], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[153]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[154], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[154]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[155], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[155]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[156], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[156]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[157], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[157]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[158], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[158]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[159], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[159]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[15]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[160], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[160]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[161], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[161]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[162], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[162]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[163], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[163]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[164], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[164]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[165], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[165]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[166], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[166]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[167], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[167]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[168], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[168]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[169], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[169]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[16]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[170], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[170]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[171], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[171]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[172], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[172]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[173], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[173]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[174], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[174]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[175], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[175]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[176], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[176]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[177], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[177]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[178], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[178]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[179], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[179]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[17]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[180], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[180]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[181], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[181]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[182], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[182]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[183], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[183]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[184], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[184]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[185], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[185]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[186], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[186]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[187], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[187]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[188], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[188]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[189], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[189]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[18]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[190], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[190]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[191], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[191]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[192], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[192]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[193], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[193]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[194], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[194]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[195], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[195]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[196], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[196]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[197], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[197]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[198], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[198]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[199], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[199]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[19]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[1]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[200], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[200]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[201], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[201]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[202], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[202]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[203], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[203]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[204], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[204]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[205], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[205]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[206], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[206]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[207], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[207]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[208], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[208]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[209], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[209]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[20]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[210], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[210]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[211], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[211]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[212], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[212]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[213], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[213]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[214], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[214]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[215], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[215]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[216], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[216]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[217], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[217]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[218], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[218]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[219], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[219]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[21]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[220], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[220]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[221], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[221]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[222], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[222]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[223], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[223]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[224], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[224]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[225], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[225]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[226], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[226]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[227], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[227]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[228], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[228]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[229], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[229]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[22]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[230], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[230]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[231], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[231]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[232], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[232]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[233], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[233]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[234], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[234]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[235], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[235]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[236], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[236]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[237], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[237]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[238], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[238]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[239], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[239]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[23]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[240], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[240]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[241], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[241]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[242], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[242]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[243], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[243]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[244], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[244]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[245], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[245]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[246], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[246]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[247], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[247]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[248], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[248]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[249], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[249]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[24]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[250], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[250]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[251], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[251]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[252], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[252]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[253], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[253]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[254], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[254]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[255], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[255]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[25]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[26]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[27]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[28]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[29]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[2]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[30]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[31]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[32], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[32]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[33], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[33]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[34], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[34]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[35], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[35]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[36], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[36]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[37], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[37]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[38], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[38]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[39], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[39]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[3]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[40], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[40]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[41], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[41]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[42], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[42]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[43], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[43]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[44], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[44]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[45], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[45]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[46], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[46]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[47], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[47]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[48], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[48]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[49], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[49]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[4]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[50], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[50]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[51], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[51]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[52], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[52]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[53], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[53]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[54], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[54]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[55], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[55]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[56], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[56]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[57], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[57]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[58], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[58]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[59], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[59]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[5]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[60], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[60]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[61], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[61]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[62], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[62]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[63], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[63]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[64], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[64]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[65], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[65]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[66], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[66]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[67], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[67]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[68], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[68]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[69], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[69]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[6]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[70], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[70]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[71], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[71]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[72], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[72]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[73], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[73]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[74], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[74]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[75], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[75]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[76], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[76]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[77], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[77]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[78], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[78]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[79], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[79]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[7]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[80], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[80]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[81], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[81]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[82], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[82]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[83], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[83]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[84], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[84]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[85], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[85]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[86], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[86]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[87], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[87]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[88], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[88]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[89], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[89]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[8]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[90], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[90]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[91], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[91]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[92], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[92]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[93], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[93]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[94], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[94]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[95], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[95]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[96], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[96]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[97], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[97]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[98], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[98]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[99], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[99]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTDATA_delay[9]);
    $setuphold (posedge USERCLK, posedge SAXISRQTKEEP[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTKEEP_delay[0]);
    $setuphold (posedge USERCLK, posedge SAXISRQTKEEP[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTKEEP_delay[1]);
    $setuphold (posedge USERCLK, posedge SAXISRQTKEEP[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTKEEP_delay[2]);
    $setuphold (posedge USERCLK, posedge SAXISRQTKEEP[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTKEEP_delay[3]);
    $setuphold (posedge USERCLK, posedge SAXISRQTKEEP[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTKEEP_delay[4]);
    $setuphold (posedge USERCLK, posedge SAXISRQTKEEP[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTKEEP_delay[5]);
    $setuphold (posedge USERCLK, posedge SAXISRQTKEEP[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTKEEP_delay[6]);
    $setuphold (posedge USERCLK, posedge SAXISRQTKEEP[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTKEEP_delay[7]);
    $setuphold (posedge USERCLK, posedge SAXISRQTLAST, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTLAST_delay);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[0], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[0]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[10], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[10]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[11], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[11]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[12], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[12]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[13], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[13]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[14], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[14]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[15], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[15]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[16], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[16]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[17], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[17]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[18], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[18]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[19], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[19]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[1], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[1]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[20], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[20]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[21], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[21]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[22], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[22]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[23], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[23]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[24], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[24]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[25], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[25]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[26], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[26]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[27], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[27]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[28], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[28]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[29], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[29]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[2], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[2]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[30], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[30]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[31], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[31]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[32], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[32]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[33], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[33]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[34], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[34]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[35], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[35]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[36], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[36]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[37], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[37]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[38], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[38]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[39], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[39]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[3], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[3]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[40], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[40]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[41], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[41]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[42], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[42]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[43], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[43]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[44], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[44]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[45], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[45]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[46], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[46]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[47], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[47]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[48], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[48]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[49], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[49]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[4], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[4]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[50], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[50]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[51], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[51]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[52], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[52]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[53], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[53]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[54], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[54]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[55], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[55]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[56], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[56]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[57], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[57]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[58], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[58]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[59], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[59]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[5], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[5]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[6], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[6]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[7], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[7]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[8], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[8]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[9], 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTUSER_delay[9]);
    $setuphold (posedge USERCLK, posedge SAXISRQTVALID, 0:0:0, 0:0:0, notifier,,, USERCLK_delay, SAXISRQTVALID_delay);
`endif
    specparam PATHPULSE$ = 0;
  endspecify

endmodule

`endcelldefine
