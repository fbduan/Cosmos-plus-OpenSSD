`include "B_OSERDESE3_ODDR_defines.vh"

reg [`OSERDESE3_ODDR_DATA_SZ-1:0] ATTR [0:`OSERDESE3_ODDR_ADDR_N-1];
reg [3:0] DATA_WIDTH_REG;
reg [0:0] INIT_REG;
reg [0:0] IS_CLKDIV_INVERTED_REG;
reg [0:0] IS_CLK_INVERTED_REG;
reg [0:0] IS_RST_INVERTED_REG;
reg [8*5:1] ODDR_MODE_REG;
reg [8*5:1] OSERDES_D_BYPASS_REG;
reg [8*5:1] OSERDES_T_BYPASS_REG;

initial begin
  ATTR[`OSERDESE3_ODDR__DATA_WIDTH] = DATA_WIDTH;
  ATTR[`OSERDESE3_ODDR__INIT] = INIT;
  ATTR[`OSERDESE3_ODDR__IS_CLKDIV_INVERTED] = IS_CLKDIV_INVERTED;
  ATTR[`OSERDESE3_ODDR__IS_CLK_INVERTED] = IS_CLK_INVERTED;
  ATTR[`OSERDESE3_ODDR__IS_RST_INVERTED] = IS_RST_INVERTED;
  ATTR[`OSERDESE3_ODDR__ODDR_MODE] = ODDR_MODE;
  ATTR[`OSERDESE3_ODDR__OSERDES_D_BYPASS] = OSERDES_D_BYPASS;
  ATTR[`OSERDESE3_ODDR__OSERDES_T_BYPASS] = OSERDES_T_BYPASS;
end

always @(trig_attr) begin
  DATA_WIDTH_REG = ATTR[`OSERDESE3_ODDR__DATA_WIDTH];
  INIT_REG = ATTR[`OSERDESE3_ODDR__INIT];
  IS_CLKDIV_INVERTED_REG = ATTR[`OSERDESE3_ODDR__IS_CLKDIV_INVERTED];
  IS_CLK_INVERTED_REG = ATTR[`OSERDESE3_ODDR__IS_CLK_INVERTED];
  IS_RST_INVERTED_REG = ATTR[`OSERDESE3_ODDR__IS_RST_INVERTED];
  ODDR_MODE_REG = ATTR[`OSERDESE3_ODDR__ODDR_MODE];
  OSERDES_D_BYPASS_REG = ATTR[`OSERDESE3_ODDR__OSERDES_D_BYPASS];
  OSERDES_T_BYPASS_REG = ATTR[`OSERDESE3_ODDR__OSERDES_T_BYPASS];
end

// procedures to override, read attribute values

task write_attr;
  input  [`OSERDESE3_ODDR_ADDR_SZ-1:0] addr;
  input  [`OSERDESE3_ODDR_DATA_SZ-1:0] data;
  begin
    ATTR[addr] = data;
    trig_attr = ~trig_attr; // to be removed
  end
endtask

function [`OSERDESE3_ODDR_DATA_SZ-1:0] read_attr;
  input  [`OSERDESE3_ODDR_ADDR_SZ-1:0] addr;
  begin
    read_attr = ATTR[addr];
  end
endfunction

task commit_attr;
  begin
    trig_attr = ~trig_attr;
  end
endtask
